module vedic32x32 (ground,
    overflow,
    A,
    B,
    Prod);
 input ground;
 output overflow;
 input [31:0] A;
 input [31:0] B;
 output [63:0] Prod;

 wire c1;
 wire c2;
 wire c3;
 wire \A1/c1 ;
 wire \A1/A1/c1 ;
 wire \A1/A1/A1/c1 ;
 wire \A1/A1/A1/A1/c1 ;
 wire \A1/A1/A1/A1/c2 ;
 wire \A1/A1/A1/A1/c3 ;
 wire \A1/A1/A1/A1/M1/c1 ;
 wire \A1/A1/A1/A1/M1/c2 ;
 wire \A1/A1/A1/A1/M1/s1 ;
 wire \A1/A1/A1/A1/M2/c1 ;
 wire \A1/A1/A1/A1/M2/c2 ;
 wire \A1/A1/A1/A1/M2/s1 ;
 wire \A1/A1/A1/A1/M3/c1 ;
 wire \A1/A1/A1/A1/M3/c2 ;
 wire \A1/A1/A1/A1/M3/s1 ;
 wire \A1/A1/A1/A1/M4/c1 ;
 wire \A1/A1/A1/A1/M4/c2 ;
 wire \A1/A1/A1/A1/M4/s1 ;
 wire \A1/A1/A1/A2/c1 ;
 wire \A1/A1/A1/A2/c2 ;
 wire \A1/A1/A1/A2/c3 ;
 wire \A1/A1/A1/A2/M1/c1 ;
 wire \A1/A1/A1/A2/M1/c2 ;
 wire \A1/A1/A1/A2/M1/s1 ;
 wire \A1/A1/A1/A2/M2/c1 ;
 wire \A1/A1/A1/A2/M2/c2 ;
 wire \A1/A1/A1/A2/M2/s1 ;
 wire \A1/A1/A1/A2/M3/c1 ;
 wire \A1/A1/A1/A2/M3/c2 ;
 wire \A1/A1/A1/A2/M3/s1 ;
 wire \A1/A1/A1/A2/M4/c1 ;
 wire \A1/A1/A1/A2/M4/c2 ;
 wire \A1/A1/A1/A2/M4/s1 ;
 wire \A1/A1/A2/c1 ;
 wire \A1/A1/A2/A1/c1 ;
 wire \A1/A1/A2/A1/c2 ;
 wire \A1/A1/A2/A1/c3 ;
 wire \A1/A1/A2/A1/M1/c1 ;
 wire \A1/A1/A2/A1/M1/c2 ;
 wire \A1/A1/A2/A1/M1/s1 ;
 wire \A1/A1/A2/A1/M2/c1 ;
 wire \A1/A1/A2/A1/M2/c2 ;
 wire \A1/A1/A2/A1/M2/s1 ;
 wire \A1/A1/A2/A1/M3/c1 ;
 wire \A1/A1/A2/A1/M3/c2 ;
 wire \A1/A1/A2/A1/M3/s1 ;
 wire \A1/A1/A2/A1/M4/c1 ;
 wire \A1/A1/A2/A1/M4/c2 ;
 wire \A1/A1/A2/A1/M4/s1 ;
 wire \A1/A1/A2/A2/c1 ;
 wire \A1/A1/A2/A2/c2 ;
 wire \A1/A1/A2/A2/c3 ;
 wire \A1/A1/A2/A2/M1/c1 ;
 wire \A1/A1/A2/A2/M1/c2 ;
 wire \A1/A1/A2/A2/M1/s1 ;
 wire \A1/A1/A2/A2/M2/c1 ;
 wire \A1/A1/A2/A2/M2/c2 ;
 wire \A1/A1/A2/A2/M2/s1 ;
 wire \A1/A1/A2/A2/M3/c1 ;
 wire \A1/A1/A2/A2/M3/c2 ;
 wire \A1/A1/A2/A2/M3/s1 ;
 wire \A1/A1/A2/A2/M4/c1 ;
 wire \A1/A1/A2/A2/M4/c2 ;
 wire \A1/A1/A2/A2/M4/s1 ;
 wire \A1/A2/c1 ;
 wire \A1/A2/A1/c1 ;
 wire \A1/A2/A1/A1/c1 ;
 wire \A1/A2/A1/A1/c2 ;
 wire \A1/A2/A1/A1/c3 ;
 wire \A1/A2/A1/A1/M1/c1 ;
 wire \A1/A2/A1/A1/M1/c2 ;
 wire \A1/A2/A1/A1/M1/s1 ;
 wire \A1/A2/A1/A1/M2/c1 ;
 wire \A1/A2/A1/A1/M2/c2 ;
 wire \A1/A2/A1/A1/M2/s1 ;
 wire \A1/A2/A1/A1/M3/c1 ;
 wire \A1/A2/A1/A1/M3/c2 ;
 wire \A1/A2/A1/A1/M3/s1 ;
 wire \A1/A2/A1/A1/M4/c1 ;
 wire \A1/A2/A1/A1/M4/c2 ;
 wire \A1/A2/A1/A1/M4/s1 ;
 wire \A1/A2/A1/A2/c1 ;
 wire \A1/A2/A1/A2/c2 ;
 wire \A1/A2/A1/A2/c3 ;
 wire \A1/A2/A1/A2/M1/c1 ;
 wire \A1/A2/A1/A2/M1/c2 ;
 wire \A1/A2/A1/A2/M1/s1 ;
 wire \A1/A2/A1/A2/M2/c1 ;
 wire \A1/A2/A1/A2/M2/c2 ;
 wire \A1/A2/A1/A2/M2/s1 ;
 wire \A1/A2/A1/A2/M3/c1 ;
 wire \A1/A2/A1/A2/M3/c2 ;
 wire \A1/A2/A1/A2/M3/s1 ;
 wire \A1/A2/A1/A2/M4/c1 ;
 wire \A1/A2/A1/A2/M4/c2 ;
 wire \A1/A2/A1/A2/M4/s1 ;
 wire \A1/A2/A2/c1 ;
 wire \A1/A2/A2/A1/c1 ;
 wire \A1/A2/A2/A1/c2 ;
 wire \A1/A2/A2/A1/c3 ;
 wire \A1/A2/A2/A1/M1/c1 ;
 wire \A1/A2/A2/A1/M1/c2 ;
 wire \A1/A2/A2/A1/M1/s1 ;
 wire \A1/A2/A2/A1/M2/c1 ;
 wire \A1/A2/A2/A1/M2/c2 ;
 wire \A1/A2/A2/A1/M2/s1 ;
 wire \A1/A2/A2/A1/M3/c1 ;
 wire \A1/A2/A2/A1/M3/c2 ;
 wire \A1/A2/A2/A1/M3/s1 ;
 wire \A1/A2/A2/A1/M4/c1 ;
 wire \A1/A2/A2/A1/M4/c2 ;
 wire \A1/A2/A2/A1/M4/s1 ;
 wire \A1/A2/A2/A2/c1 ;
 wire \A1/A2/A2/A2/c2 ;
 wire \A1/A2/A2/A2/c3 ;
 wire \A1/A2/A2/A2/M1/c1 ;
 wire \A1/A2/A2/A2/M1/c2 ;
 wire \A1/A2/A2/A2/M1/s1 ;
 wire \A1/A2/A2/A2/M2/c1 ;
 wire \A1/A2/A2/A2/M2/c2 ;
 wire \A1/A2/A2/A2/M2/s1 ;
 wire \A1/A2/A2/A2/M3/c1 ;
 wire \A1/A2/A2/A2/M3/c2 ;
 wire \A1/A2/A2/A2/M3/s1 ;
 wire \A1/A2/A2/A2/M4/c1 ;
 wire \A1/A2/A2/A2/M4/c2 ;
 wire \A1/A2/A2/A2/M4/s1 ;
 wire \A2/c1 ;
 wire \A2/A1/c1 ;
 wire \A2/A1/A1/c1 ;
 wire \A2/A1/A1/A1/c1 ;
 wire \A2/A1/A1/A1/c2 ;
 wire \A2/A1/A1/A1/c3 ;
 wire \A2/A1/A1/A1/M1/c1 ;
 wire \A2/A1/A1/A1/M1/c2 ;
 wire \A2/A1/A1/A1/M1/s1 ;
 wire \A2/A1/A1/A1/M2/c1 ;
 wire \A2/A1/A1/A1/M2/c2 ;
 wire \A2/A1/A1/A1/M2/s1 ;
 wire \A2/A1/A1/A1/M3/c1 ;
 wire \A2/A1/A1/A1/M3/c2 ;
 wire \A2/A1/A1/A1/M3/s1 ;
 wire \A2/A1/A1/A1/M4/c1 ;
 wire \A2/A1/A1/A1/M4/c2 ;
 wire \A2/A1/A1/A1/M4/s1 ;
 wire \A2/A1/A1/A2/c1 ;
 wire \A2/A1/A1/A2/c2 ;
 wire \A2/A1/A1/A2/c3 ;
 wire \A2/A1/A1/A2/M1/c1 ;
 wire \A2/A1/A1/A2/M1/c2 ;
 wire \A2/A1/A1/A2/M1/s1 ;
 wire \A2/A1/A1/A2/M2/c1 ;
 wire \A2/A1/A1/A2/M2/c2 ;
 wire \A2/A1/A1/A2/M2/s1 ;
 wire \A2/A1/A1/A2/M3/c1 ;
 wire \A2/A1/A1/A2/M3/c2 ;
 wire \A2/A1/A1/A2/M3/s1 ;
 wire \A2/A1/A1/A2/M4/c1 ;
 wire \A2/A1/A1/A2/M4/c2 ;
 wire \A2/A1/A1/A2/M4/s1 ;
 wire \A2/A1/A2/c1 ;
 wire \A2/A1/A2/A1/c1 ;
 wire \A2/A1/A2/A1/c2 ;
 wire \A2/A1/A2/A1/c3 ;
 wire \A2/A1/A2/A1/M1/c1 ;
 wire \A2/A1/A2/A1/M1/c2 ;
 wire \A2/A1/A2/A1/M1/s1 ;
 wire \A2/A1/A2/A1/M2/c1 ;
 wire \A2/A1/A2/A1/M2/c2 ;
 wire \A2/A1/A2/A1/M2/s1 ;
 wire \A2/A1/A2/A1/M3/c1 ;
 wire \A2/A1/A2/A1/M3/c2 ;
 wire \A2/A1/A2/A1/M3/s1 ;
 wire \A2/A1/A2/A1/M4/c1 ;
 wire \A2/A1/A2/A1/M4/c2 ;
 wire \A2/A1/A2/A1/M4/s1 ;
 wire \A2/A1/A2/A2/c1 ;
 wire \A2/A1/A2/A2/c2 ;
 wire \A2/A1/A2/A2/c3 ;
 wire \A2/A1/A2/A2/M1/c1 ;
 wire \A2/A1/A2/A2/M1/c2 ;
 wire \A2/A1/A2/A2/M1/s1 ;
 wire \A2/A1/A2/A2/M2/c1 ;
 wire \A2/A1/A2/A2/M2/c2 ;
 wire \A2/A1/A2/A2/M2/s1 ;
 wire \A2/A1/A2/A2/M3/c1 ;
 wire \A2/A1/A2/A2/M3/c2 ;
 wire \A2/A1/A2/A2/M3/s1 ;
 wire \A2/A1/A2/A2/M4/c1 ;
 wire \A2/A1/A2/A2/M4/c2 ;
 wire \A2/A1/A2/A2/M4/s1 ;
 wire \A2/A2/c1 ;
 wire \A2/A2/A1/c1 ;
 wire \A2/A2/A1/A1/c1 ;
 wire \A2/A2/A1/A1/c2 ;
 wire \A2/A2/A1/A1/c3 ;
 wire \A2/A2/A1/A1/M1/c1 ;
 wire \A2/A2/A1/A1/M1/c2 ;
 wire \A2/A2/A1/A1/M1/s1 ;
 wire \A2/A2/A1/A1/M2/c1 ;
 wire \A2/A2/A1/A1/M2/c2 ;
 wire \A2/A2/A1/A1/M2/s1 ;
 wire \A2/A2/A1/A1/M3/c1 ;
 wire \A2/A2/A1/A1/M3/c2 ;
 wire \A2/A2/A1/A1/M3/s1 ;
 wire \A2/A2/A1/A1/M4/c1 ;
 wire \A2/A2/A1/A1/M4/c2 ;
 wire \A2/A2/A1/A1/M4/s1 ;
 wire \A2/A2/A1/A2/c1 ;
 wire \A2/A2/A1/A2/c2 ;
 wire \A2/A2/A1/A2/c3 ;
 wire \A2/A2/A1/A2/M1/c1 ;
 wire \A2/A2/A1/A2/M1/c2 ;
 wire \A2/A2/A1/A2/M1/s1 ;
 wire \A2/A2/A1/A2/M2/c1 ;
 wire \A2/A2/A1/A2/M2/c2 ;
 wire \A2/A2/A1/A2/M2/s1 ;
 wire \A2/A2/A1/A2/M3/c1 ;
 wire \A2/A2/A1/A2/M3/c2 ;
 wire \A2/A2/A1/A2/M3/s1 ;
 wire \A2/A2/A1/A2/M4/c1 ;
 wire \A2/A2/A1/A2/M4/c2 ;
 wire \A2/A2/A1/A2/M4/s1 ;
 wire \A2/A2/A2/c1 ;
 wire \A2/A2/A2/A1/c1 ;
 wire \A2/A2/A2/A1/c2 ;
 wire \A2/A2/A2/A1/c3 ;
 wire \A2/A2/A2/A1/M1/c1 ;
 wire \A2/A2/A2/A1/M1/c2 ;
 wire \A2/A2/A2/A1/M1/s1 ;
 wire \A2/A2/A2/A1/M2/c1 ;
 wire \A2/A2/A2/A1/M2/c2 ;
 wire \A2/A2/A2/A1/M2/s1 ;
 wire \A2/A2/A2/A1/M3/c1 ;
 wire \A2/A2/A2/A1/M3/c2 ;
 wire \A2/A2/A2/A1/M3/s1 ;
 wire \A2/A2/A2/A1/M4/c1 ;
 wire \A2/A2/A2/A1/M4/c2 ;
 wire \A2/A2/A2/A1/M4/s1 ;
 wire \A2/A2/A2/A2/c1 ;
 wire \A2/A2/A2/A2/c2 ;
 wire \A2/A2/A2/A2/c3 ;
 wire \A2/A2/A2/A2/M1/c1 ;
 wire \A2/A2/A2/A2/M1/c2 ;
 wire \A2/A2/A2/A2/M1/s1 ;
 wire \A2/A2/A2/A2/M2/c1 ;
 wire \A2/A2/A2/A2/M2/c2 ;
 wire \A2/A2/A2/A2/M2/s1 ;
 wire \A2/A2/A2/A2/M3/c1 ;
 wire \A2/A2/A2/A2/M3/c2 ;
 wire \A2/A2/A2/A2/M3/s1 ;
 wire \A2/A2/A2/A2/M4/c1 ;
 wire \A2/A2/A2/A2/M4/c2 ;
 wire \A2/A2/A2/A2/M4/s1 ;
 wire \A3/c1 ;
 wire \A3/A1/c1 ;
 wire \A3/A1/A1/c1 ;
 wire \A3/A1/A1/A1/c1 ;
 wire \A3/A1/A1/A1/c2 ;
 wire \A3/A1/A1/A1/c3 ;
 wire \A3/A1/A1/A1/M1/c1 ;
 wire \A3/A1/A1/A1/M1/c2 ;
 wire \A3/A1/A1/A1/M1/s1 ;
 wire \A3/A1/A1/A1/M2/c1 ;
 wire \A3/A1/A1/A1/M2/c2 ;
 wire \A3/A1/A1/A1/M2/s1 ;
 wire \A3/A1/A1/A1/M3/c1 ;
 wire \A3/A1/A1/A1/M3/c2 ;
 wire \A3/A1/A1/A1/M3/s1 ;
 wire \A3/A1/A1/A1/M4/c1 ;
 wire \A3/A1/A1/A1/M4/c2 ;
 wire \A3/A1/A1/A1/M4/s1 ;
 wire \A3/A1/A1/A2/c1 ;
 wire \A3/A1/A1/A2/c2 ;
 wire \A3/A1/A1/A2/c3 ;
 wire \A3/A1/A1/A2/M1/c1 ;
 wire \A3/A1/A1/A2/M1/c2 ;
 wire \A3/A1/A1/A2/M1/s1 ;
 wire \A3/A1/A1/A2/M2/c1 ;
 wire \A3/A1/A1/A2/M2/c2 ;
 wire \A3/A1/A1/A2/M2/s1 ;
 wire \A3/A1/A1/A2/M3/c1 ;
 wire \A3/A1/A1/A2/M3/c2 ;
 wire \A3/A1/A1/A2/M3/s1 ;
 wire \A3/A1/A1/A2/M4/c1 ;
 wire \A3/A1/A1/A2/M4/c2 ;
 wire \A3/A1/A1/A2/M4/s1 ;
 wire \A3/A1/A2/c1 ;
 wire \A3/A1/A2/A1/c1 ;
 wire \A3/A1/A2/A1/c2 ;
 wire \A3/A1/A2/A1/c3 ;
 wire \A3/A1/A2/A1/M1/c1 ;
 wire \A3/A1/A2/A1/M1/c2 ;
 wire \A3/A1/A2/A1/M1/s1 ;
 wire \A3/A1/A2/A1/M2/c1 ;
 wire \A3/A1/A2/A1/M2/c2 ;
 wire \A3/A1/A2/A1/M2/s1 ;
 wire \A3/A1/A2/A1/M3/c1 ;
 wire \A3/A1/A2/A1/M3/c2 ;
 wire \A3/A1/A2/A1/M3/s1 ;
 wire \A3/A1/A2/A1/M4/c1 ;
 wire \A3/A1/A2/A1/M4/c2 ;
 wire \A3/A1/A2/A1/M4/s1 ;
 wire \A3/A1/A2/A2/c1 ;
 wire \A3/A1/A2/A2/c2 ;
 wire \A3/A1/A2/A2/c3 ;
 wire \A3/A1/A2/A2/M1/c1 ;
 wire \A3/A1/A2/A2/M1/c2 ;
 wire \A3/A1/A2/A2/M1/s1 ;
 wire \A3/A1/A2/A2/M2/c1 ;
 wire \A3/A1/A2/A2/M2/c2 ;
 wire \A3/A1/A2/A2/M2/s1 ;
 wire \A3/A1/A2/A2/M3/c1 ;
 wire \A3/A1/A2/A2/M3/c2 ;
 wire \A3/A1/A2/A2/M3/s1 ;
 wire \A3/A1/A2/A2/M4/c1 ;
 wire \A3/A1/A2/A2/M4/c2 ;
 wire \A3/A1/A2/A2/M4/s1 ;
 wire \A3/A2/c1 ;
 wire \A3/A2/A1/c1 ;
 wire \A3/A2/A1/A1/c1 ;
 wire \A3/A2/A1/A1/c2 ;
 wire \A3/A2/A1/A1/c3 ;
 wire \A3/A2/A1/A1/M1/c1 ;
 wire \A3/A2/A1/A1/M1/c2 ;
 wire \A3/A2/A1/A1/M1/s1 ;
 wire \A3/A2/A1/A1/M2/c1 ;
 wire \A3/A2/A1/A1/M2/c2 ;
 wire \A3/A2/A1/A1/M2/s1 ;
 wire \A3/A2/A1/A1/M3/c1 ;
 wire \A3/A2/A1/A1/M3/c2 ;
 wire \A3/A2/A1/A1/M3/s1 ;
 wire \A3/A2/A1/A1/M4/c1 ;
 wire \A3/A2/A1/A1/M4/c2 ;
 wire \A3/A2/A1/A1/M4/s1 ;
 wire \A3/A2/A1/A2/c1 ;
 wire \A3/A2/A1/A2/c2 ;
 wire \A3/A2/A1/A2/c3 ;
 wire \A3/A2/A1/A2/M1/c1 ;
 wire \A3/A2/A1/A2/M1/c2 ;
 wire \A3/A2/A1/A2/M1/s1 ;
 wire \A3/A2/A1/A2/M2/c1 ;
 wire \A3/A2/A1/A2/M2/c2 ;
 wire \A3/A2/A1/A2/M2/s1 ;
 wire \A3/A2/A1/A2/M3/c1 ;
 wire \A3/A2/A1/A2/M3/c2 ;
 wire \A3/A2/A1/A2/M3/s1 ;
 wire \A3/A2/A1/A2/M4/c1 ;
 wire \A3/A2/A1/A2/M4/c2 ;
 wire \A3/A2/A1/A2/M4/s1 ;
 wire \A3/A2/A2/c1 ;
 wire \A3/A2/A2/A1/c1 ;
 wire \A3/A2/A2/A1/c2 ;
 wire \A3/A2/A2/A1/c3 ;
 wire \A3/A2/A2/A1/M1/c1 ;
 wire \A3/A2/A2/A1/M1/c2 ;
 wire \A3/A2/A2/A1/M1/s1 ;
 wire \A3/A2/A2/A1/M2/c1 ;
 wire \A3/A2/A2/A1/M2/c2 ;
 wire \A3/A2/A2/A1/M2/s1 ;
 wire \A3/A2/A2/A1/M3/c1 ;
 wire \A3/A2/A2/A1/M3/c2 ;
 wire \A3/A2/A2/A1/M3/s1 ;
 wire \A3/A2/A2/A1/M4/c1 ;
 wire \A3/A2/A2/A1/M4/c2 ;
 wire \A3/A2/A2/A1/M4/s1 ;
 wire \A3/A2/A2/A2/c1 ;
 wire \A3/A2/A2/A2/c2 ;
 wire \A3/A2/A2/A2/c3 ;
 wire \A3/A2/A2/A2/M1/c1 ;
 wire \A3/A2/A2/A2/M1/c2 ;
 wire \A3/A2/A2/A2/M1/s1 ;
 wire \A3/A2/A2/A2/M2/c1 ;
 wire \A3/A2/A2/A2/M2/c2 ;
 wire \A3/A2/A2/A2/M2/s1 ;
 wire \A3/A2/A2/A2/M3/c1 ;
 wire \A3/A2/A2/A2/M3/c2 ;
 wire \A3/A2/A2/A2/M3/s1 ;
 wire \A3/A2/A2/A2/M4/c1 ;
 wire \A3/A2/A2/A2/M4/c2 ;
 wire \A3/A2/A2/A2/M4/s1 ;
 wire \V1/c1 ;
 wire \V1/c2 ;
 wire \V1/c3 ;
 wire \V1/overflow ;
 wire \V1/A1/c1 ;
 wire \V1/A1/A1/c1 ;
 wire \V1/A1/A1/A1/c1 ;
 wire \V1/A1/A1/A1/c2 ;
 wire \V1/A1/A1/A1/c3 ;
 wire \V1/A1/A1/A1/M1/c1 ;
 wire \V1/A1/A1/A1/M1/c2 ;
 wire \V1/A1/A1/A1/M1/s1 ;
 wire \V1/A1/A1/A1/M2/c1 ;
 wire \V1/A1/A1/A1/M2/c2 ;
 wire \V1/A1/A1/A1/M2/s1 ;
 wire \V1/A1/A1/A1/M3/c1 ;
 wire \V1/A1/A1/A1/M3/c2 ;
 wire \V1/A1/A1/A1/M3/s1 ;
 wire \V1/A1/A1/A1/M4/c1 ;
 wire \V1/A1/A1/A1/M4/c2 ;
 wire \V1/A1/A1/A1/M4/s1 ;
 wire \V1/A1/A1/A2/c1 ;
 wire \V1/A1/A1/A2/c2 ;
 wire \V1/A1/A1/A2/c3 ;
 wire \V1/A1/A1/A2/M1/c1 ;
 wire \V1/A1/A1/A2/M1/c2 ;
 wire \V1/A1/A1/A2/M1/s1 ;
 wire \V1/A1/A1/A2/M2/c1 ;
 wire \V1/A1/A1/A2/M2/c2 ;
 wire \V1/A1/A1/A2/M2/s1 ;
 wire \V1/A1/A1/A2/M3/c1 ;
 wire \V1/A1/A1/A2/M3/c2 ;
 wire \V1/A1/A1/A2/M3/s1 ;
 wire \V1/A1/A1/A2/M4/c1 ;
 wire \V1/A1/A1/A2/M4/c2 ;
 wire \V1/A1/A1/A2/M4/s1 ;
 wire \V1/A1/A2/c1 ;
 wire \V1/A1/A2/A1/c1 ;
 wire \V1/A1/A2/A1/c2 ;
 wire \V1/A1/A2/A1/c3 ;
 wire \V1/A1/A2/A1/M1/c1 ;
 wire \V1/A1/A2/A1/M1/c2 ;
 wire \V1/A1/A2/A1/M1/s1 ;
 wire \V1/A1/A2/A1/M2/c1 ;
 wire \V1/A1/A2/A1/M2/c2 ;
 wire \V1/A1/A2/A1/M2/s1 ;
 wire \V1/A1/A2/A1/M3/c1 ;
 wire \V1/A1/A2/A1/M3/c2 ;
 wire \V1/A1/A2/A1/M3/s1 ;
 wire \V1/A1/A2/A1/M4/c1 ;
 wire \V1/A1/A2/A1/M4/c2 ;
 wire \V1/A1/A2/A1/M4/s1 ;
 wire \V1/A1/A2/A2/c1 ;
 wire \V1/A1/A2/A2/c2 ;
 wire \V1/A1/A2/A2/c3 ;
 wire \V1/A1/A2/A2/M1/c1 ;
 wire \V1/A1/A2/A2/M1/c2 ;
 wire \V1/A1/A2/A2/M1/s1 ;
 wire \V1/A1/A2/A2/M2/c1 ;
 wire \V1/A1/A2/A2/M2/c2 ;
 wire \V1/A1/A2/A2/M2/s1 ;
 wire \V1/A1/A2/A2/M3/c1 ;
 wire \V1/A1/A2/A2/M3/c2 ;
 wire \V1/A1/A2/A2/M3/s1 ;
 wire \V1/A1/A2/A2/M4/c1 ;
 wire \V1/A1/A2/A2/M4/c2 ;
 wire \V1/A1/A2/A2/M4/s1 ;
 wire \V1/A2/c1 ;
 wire \V1/A2/A1/c1 ;
 wire \V1/A2/A1/A1/c1 ;
 wire \V1/A2/A1/A1/c2 ;
 wire \V1/A2/A1/A1/c3 ;
 wire \V1/A2/A1/A1/M1/c1 ;
 wire \V1/A2/A1/A1/M1/c2 ;
 wire \V1/A2/A1/A1/M1/s1 ;
 wire \V1/A2/A1/A1/M2/c1 ;
 wire \V1/A2/A1/A1/M2/c2 ;
 wire \V1/A2/A1/A1/M2/s1 ;
 wire \V1/A2/A1/A1/M3/c1 ;
 wire \V1/A2/A1/A1/M3/c2 ;
 wire \V1/A2/A1/A1/M3/s1 ;
 wire \V1/A2/A1/A1/M4/c1 ;
 wire \V1/A2/A1/A1/M4/c2 ;
 wire \V1/A2/A1/A1/M4/s1 ;
 wire \V1/A2/A1/A2/c1 ;
 wire \V1/A2/A1/A2/c2 ;
 wire \V1/A2/A1/A2/c3 ;
 wire \V1/A2/A1/A2/M1/c1 ;
 wire \V1/A2/A1/A2/M1/c2 ;
 wire \V1/A2/A1/A2/M1/s1 ;
 wire \V1/A2/A1/A2/M2/c1 ;
 wire \V1/A2/A1/A2/M2/c2 ;
 wire \V1/A2/A1/A2/M2/s1 ;
 wire \V1/A2/A1/A2/M3/c1 ;
 wire \V1/A2/A1/A2/M3/c2 ;
 wire \V1/A2/A1/A2/M3/s1 ;
 wire \V1/A2/A1/A2/M4/c1 ;
 wire \V1/A2/A1/A2/M4/c2 ;
 wire \V1/A2/A1/A2/M4/s1 ;
 wire \V1/A2/A2/c1 ;
 wire \V1/A2/A2/A1/c1 ;
 wire \V1/A2/A2/A1/c2 ;
 wire \V1/A2/A2/A1/c3 ;
 wire \V1/A2/A2/A1/M1/c1 ;
 wire \V1/A2/A2/A1/M1/c2 ;
 wire \V1/A2/A2/A1/M1/s1 ;
 wire \V1/A2/A2/A1/M2/c1 ;
 wire \V1/A2/A2/A1/M2/c2 ;
 wire \V1/A2/A2/A1/M2/s1 ;
 wire \V1/A2/A2/A1/M3/c1 ;
 wire \V1/A2/A2/A1/M3/c2 ;
 wire \V1/A2/A2/A1/M3/s1 ;
 wire \V1/A2/A2/A1/M4/c1 ;
 wire \V1/A2/A2/A1/M4/c2 ;
 wire \V1/A2/A2/A1/M4/s1 ;
 wire \V1/A2/A2/A2/c1 ;
 wire \V1/A2/A2/A2/c2 ;
 wire \V1/A2/A2/A2/c3 ;
 wire \V1/A2/A2/A2/M1/c1 ;
 wire \V1/A2/A2/A2/M1/c2 ;
 wire \V1/A2/A2/A2/M1/s1 ;
 wire \V1/A2/A2/A2/M2/c1 ;
 wire \V1/A2/A2/A2/M2/c2 ;
 wire \V1/A2/A2/A2/M2/s1 ;
 wire \V1/A2/A2/A2/M3/c1 ;
 wire \V1/A2/A2/A2/M3/c2 ;
 wire \V1/A2/A2/A2/M3/s1 ;
 wire \V1/A2/A2/A2/M4/c1 ;
 wire \V1/A2/A2/A2/M4/c2 ;
 wire \V1/A2/A2/A2/M4/s1 ;
 wire \V1/A3/c1 ;
 wire \V1/A3/A1/c1 ;
 wire \V1/A3/A1/A1/c1 ;
 wire \V1/A3/A1/A1/c2 ;
 wire \V1/A3/A1/A1/c3 ;
 wire \V1/A3/A1/A1/M1/c1 ;
 wire \V1/A3/A1/A1/M1/c2 ;
 wire \V1/A3/A1/A1/M1/s1 ;
 wire \V1/A3/A1/A1/M2/c1 ;
 wire \V1/A3/A1/A1/M2/c2 ;
 wire \V1/A3/A1/A1/M2/s1 ;
 wire \V1/A3/A1/A1/M3/c1 ;
 wire \V1/A3/A1/A1/M3/c2 ;
 wire \V1/A3/A1/A1/M3/s1 ;
 wire \V1/A3/A1/A1/M4/c1 ;
 wire \V1/A3/A1/A1/M4/c2 ;
 wire \V1/A3/A1/A1/M4/s1 ;
 wire \V1/A3/A1/A2/c1 ;
 wire \V1/A3/A1/A2/c2 ;
 wire \V1/A3/A1/A2/c3 ;
 wire \V1/A3/A1/A2/M1/c1 ;
 wire \V1/A3/A1/A2/M1/c2 ;
 wire \V1/A3/A1/A2/M1/s1 ;
 wire \V1/A3/A1/A2/M2/c1 ;
 wire \V1/A3/A1/A2/M2/c2 ;
 wire \V1/A3/A1/A2/M2/s1 ;
 wire \V1/A3/A1/A2/M3/c1 ;
 wire \V1/A3/A1/A2/M3/c2 ;
 wire \V1/A3/A1/A2/M3/s1 ;
 wire \V1/A3/A1/A2/M4/c1 ;
 wire \V1/A3/A1/A2/M4/c2 ;
 wire \V1/A3/A1/A2/M4/s1 ;
 wire \V1/A3/A2/c1 ;
 wire \V1/A3/A2/A1/c1 ;
 wire \V1/A3/A2/A1/c2 ;
 wire \V1/A3/A2/A1/c3 ;
 wire \V1/A3/A2/A1/M1/c1 ;
 wire \V1/A3/A2/A1/M1/c2 ;
 wire \V1/A3/A2/A1/M1/s1 ;
 wire \V1/A3/A2/A1/M2/c1 ;
 wire \V1/A3/A2/A1/M2/c2 ;
 wire \V1/A3/A2/A1/M2/s1 ;
 wire \V1/A3/A2/A1/M3/c1 ;
 wire \V1/A3/A2/A1/M3/c2 ;
 wire \V1/A3/A2/A1/M3/s1 ;
 wire \V1/A3/A2/A1/M4/c1 ;
 wire \V1/A3/A2/A1/M4/c2 ;
 wire \V1/A3/A2/A1/M4/s1 ;
 wire \V1/A3/A2/A2/c1 ;
 wire \V1/A3/A2/A2/c2 ;
 wire \V1/A3/A2/A2/c3 ;
 wire \V1/A3/A2/A2/M1/c1 ;
 wire \V1/A3/A2/A2/M1/c2 ;
 wire \V1/A3/A2/A2/M1/s1 ;
 wire \V1/A3/A2/A2/M2/c1 ;
 wire \V1/A3/A2/A2/M2/c2 ;
 wire \V1/A3/A2/A2/M2/s1 ;
 wire \V1/A3/A2/A2/M3/c1 ;
 wire \V1/A3/A2/A2/M3/c2 ;
 wire \V1/A3/A2/A2/M3/s1 ;
 wire \V1/A3/A2/A2/M4/c1 ;
 wire \V1/A3/A2/A2/M4/c2 ;
 wire \V1/A3/A2/A2/M4/s1 ;
 wire \V1/V1/c1 ;
 wire \V1/V1/c2 ;
 wire \V1/V1/c3 ;
 wire \V1/V1/overflow ;
 wire \V1/V1/A1/c1 ;
 wire \V1/V1/A1/A1/c1 ;
 wire \V1/V1/A1/A1/c2 ;
 wire \V1/V1/A1/A1/c3 ;
 wire \V1/V1/A1/A1/M1/c1 ;
 wire \V1/V1/A1/A1/M1/c2 ;
 wire \V1/V1/A1/A1/M1/s1 ;
 wire \V1/V1/A1/A1/M2/c1 ;
 wire \V1/V1/A1/A1/M2/c2 ;
 wire \V1/V1/A1/A1/M2/s1 ;
 wire \V1/V1/A1/A1/M3/c1 ;
 wire \V1/V1/A1/A1/M3/c2 ;
 wire \V1/V1/A1/A1/M3/s1 ;
 wire \V1/V1/A1/A1/M4/c1 ;
 wire \V1/V1/A1/A1/M4/c2 ;
 wire \V1/V1/A1/A1/M4/s1 ;
 wire \V1/V1/A1/A2/c1 ;
 wire \V1/V1/A1/A2/c2 ;
 wire \V1/V1/A1/A2/c3 ;
 wire \V1/V1/A1/A2/M1/c1 ;
 wire \V1/V1/A1/A2/M1/c2 ;
 wire \V1/V1/A1/A2/M1/s1 ;
 wire \V1/V1/A1/A2/M2/c1 ;
 wire \V1/V1/A1/A2/M2/c2 ;
 wire \V1/V1/A1/A2/M2/s1 ;
 wire \V1/V1/A1/A2/M3/c1 ;
 wire \V1/V1/A1/A2/M3/c2 ;
 wire \V1/V1/A1/A2/M3/s1 ;
 wire \V1/V1/A1/A2/M4/c1 ;
 wire \V1/V1/A1/A2/M4/c2 ;
 wire \V1/V1/A1/A2/M4/s1 ;
 wire \V1/V1/A2/c1 ;
 wire \V1/V1/A2/A1/c1 ;
 wire \V1/V1/A2/A1/c2 ;
 wire \V1/V1/A2/A1/c3 ;
 wire \V1/V1/A2/A1/M1/c1 ;
 wire \V1/V1/A2/A1/M1/c2 ;
 wire \V1/V1/A2/A1/M1/s1 ;
 wire \V1/V1/A2/A1/M2/c1 ;
 wire \V1/V1/A2/A1/M2/c2 ;
 wire \V1/V1/A2/A1/M2/s1 ;
 wire \V1/V1/A2/A1/M3/c1 ;
 wire \V1/V1/A2/A1/M3/c2 ;
 wire \V1/V1/A2/A1/M3/s1 ;
 wire \V1/V1/A2/A1/M4/c1 ;
 wire \V1/V1/A2/A1/M4/c2 ;
 wire \V1/V1/A2/A1/M4/s1 ;
 wire \V1/V1/A2/A2/c1 ;
 wire \V1/V1/A2/A2/c2 ;
 wire \V1/V1/A2/A2/c3 ;
 wire \V1/V1/A2/A2/M1/c1 ;
 wire \V1/V1/A2/A2/M1/c2 ;
 wire \V1/V1/A2/A2/M1/s1 ;
 wire \V1/V1/A2/A2/M2/c1 ;
 wire \V1/V1/A2/A2/M2/c2 ;
 wire \V1/V1/A2/A2/M2/s1 ;
 wire \V1/V1/A2/A2/M3/c1 ;
 wire \V1/V1/A2/A2/M3/c2 ;
 wire \V1/V1/A2/A2/M3/s1 ;
 wire \V1/V1/A2/A2/M4/c1 ;
 wire \V1/V1/A2/A2/M4/c2 ;
 wire \V1/V1/A2/A2/M4/s1 ;
 wire \V1/V1/A3/c1 ;
 wire \V1/V1/A3/A1/c1 ;
 wire \V1/V1/A3/A1/c2 ;
 wire \V1/V1/A3/A1/c3 ;
 wire \V1/V1/A3/A1/M1/c1 ;
 wire \V1/V1/A3/A1/M1/c2 ;
 wire \V1/V1/A3/A1/M1/s1 ;
 wire \V1/V1/A3/A1/M2/c1 ;
 wire \V1/V1/A3/A1/M2/c2 ;
 wire \V1/V1/A3/A1/M2/s1 ;
 wire \V1/V1/A3/A1/M3/c1 ;
 wire \V1/V1/A3/A1/M3/c2 ;
 wire \V1/V1/A3/A1/M3/s1 ;
 wire \V1/V1/A3/A1/M4/c1 ;
 wire \V1/V1/A3/A1/M4/c2 ;
 wire \V1/V1/A3/A1/M4/s1 ;
 wire \V1/V1/A3/A2/c1 ;
 wire \V1/V1/A3/A2/c2 ;
 wire \V1/V1/A3/A2/c3 ;
 wire \V1/V1/A3/A2/M1/c1 ;
 wire \V1/V1/A3/A2/M1/c2 ;
 wire \V1/V1/A3/A2/M1/s1 ;
 wire \V1/V1/A3/A2/M2/c1 ;
 wire \V1/V1/A3/A2/M2/c2 ;
 wire \V1/V1/A3/A2/M2/s1 ;
 wire \V1/V1/A3/A2/M3/c1 ;
 wire \V1/V1/A3/A2/M3/c2 ;
 wire \V1/V1/A3/A2/M3/s1 ;
 wire \V1/V1/A3/A2/M4/c1 ;
 wire \V1/V1/A3/A2/M4/c2 ;
 wire \V1/V1/A3/A2/M4/s1 ;
 wire \V1/V1/V1/c1 ;
 wire \V1/V1/V1/c2 ;
 wire \V1/V1/V1/c3 ;
 wire \V1/V1/V1/overflow ;
 wire \V1/V1/V1/A1/c1 ;
 wire \V1/V1/V1/A1/c2 ;
 wire \V1/V1/V1/A1/c3 ;
 wire \V1/V1/V1/A1/M1/c1 ;
 wire \V1/V1/V1/A1/M1/c2 ;
 wire \V1/V1/V1/A1/M1/s1 ;
 wire \V1/V1/V1/A1/M2/c1 ;
 wire \V1/V1/V1/A1/M2/c2 ;
 wire \V1/V1/V1/A1/M2/s1 ;
 wire \V1/V1/V1/A1/M3/c1 ;
 wire \V1/V1/V1/A1/M3/c2 ;
 wire \V1/V1/V1/A1/M3/s1 ;
 wire \V1/V1/V1/A1/M4/c1 ;
 wire \V1/V1/V1/A1/M4/c2 ;
 wire \V1/V1/V1/A1/M4/s1 ;
 wire \V1/V1/V1/A2/c1 ;
 wire \V1/V1/V1/A2/c2 ;
 wire \V1/V1/V1/A2/c3 ;
 wire \V1/V1/V1/A2/M1/c1 ;
 wire \V1/V1/V1/A2/M1/c2 ;
 wire \V1/V1/V1/A2/M1/s1 ;
 wire \V1/V1/V1/A2/M2/c1 ;
 wire \V1/V1/V1/A2/M2/c2 ;
 wire \V1/V1/V1/A2/M2/s1 ;
 wire \V1/V1/V1/A2/M3/c1 ;
 wire \V1/V1/V1/A2/M3/c2 ;
 wire \V1/V1/V1/A2/M3/s1 ;
 wire \V1/V1/V1/A2/M4/c1 ;
 wire \V1/V1/V1/A2/M4/c2 ;
 wire \V1/V1/V1/A2/M4/s1 ;
 wire \V1/V1/V1/A3/c1 ;
 wire \V1/V1/V1/A3/c2 ;
 wire \V1/V1/V1/A3/c3 ;
 wire \V1/V1/V1/A3/M1/c1 ;
 wire \V1/V1/V1/A3/M1/c2 ;
 wire \V1/V1/V1/A3/M1/s1 ;
 wire \V1/V1/V1/A3/M2/c1 ;
 wire \V1/V1/V1/A3/M2/c2 ;
 wire \V1/V1/V1/A3/M2/s1 ;
 wire \V1/V1/V1/A3/M3/c1 ;
 wire \V1/V1/V1/A3/M3/c2 ;
 wire \V1/V1/V1/A3/M3/s1 ;
 wire \V1/V1/V1/A3/M4/c1 ;
 wire \V1/V1/V1/A3/M4/c2 ;
 wire \V1/V1/V1/A3/M4/s1 ;
 wire \V1/V1/V1/V1/w1 ;
 wire \V1/V1/V1/V1/w2 ;
 wire \V1/V1/V1/V1/w3 ;
 wire \V1/V1/V1/V1/w4 ;
 wire \V1/V1/V1/V2/w1 ;
 wire \V1/V1/V1/V2/w2 ;
 wire \V1/V1/V1/V2/w3 ;
 wire \V1/V1/V1/V2/w4 ;
 wire \V1/V1/V1/V3/w1 ;
 wire \V1/V1/V1/V3/w2 ;
 wire \V1/V1/V1/V3/w3 ;
 wire \V1/V1/V1/V3/w4 ;
 wire \V1/V1/V1/V4/w1 ;
 wire \V1/V1/V1/V4/w2 ;
 wire \V1/V1/V1/V4/w3 ;
 wire \V1/V1/V1/V4/w4 ;
 wire \V1/V1/V2/c1 ;
 wire \V1/V1/V2/c2 ;
 wire \V1/V1/V2/c3 ;
 wire \V1/V1/V2/overflow ;
 wire \V1/V1/V2/A1/c1 ;
 wire \V1/V1/V2/A1/c2 ;
 wire \V1/V1/V2/A1/c3 ;
 wire \V1/V1/V2/A1/M1/c1 ;
 wire \V1/V1/V2/A1/M1/c2 ;
 wire \V1/V1/V2/A1/M1/s1 ;
 wire \V1/V1/V2/A1/M2/c1 ;
 wire \V1/V1/V2/A1/M2/c2 ;
 wire \V1/V1/V2/A1/M2/s1 ;
 wire \V1/V1/V2/A1/M3/c1 ;
 wire \V1/V1/V2/A1/M3/c2 ;
 wire \V1/V1/V2/A1/M3/s1 ;
 wire \V1/V1/V2/A1/M4/c1 ;
 wire \V1/V1/V2/A1/M4/c2 ;
 wire \V1/V1/V2/A1/M4/s1 ;
 wire \V1/V1/V2/A2/c1 ;
 wire \V1/V1/V2/A2/c2 ;
 wire \V1/V1/V2/A2/c3 ;
 wire \V1/V1/V2/A2/M1/c1 ;
 wire \V1/V1/V2/A2/M1/c2 ;
 wire \V1/V1/V2/A2/M1/s1 ;
 wire \V1/V1/V2/A2/M2/c1 ;
 wire \V1/V1/V2/A2/M2/c2 ;
 wire \V1/V1/V2/A2/M2/s1 ;
 wire \V1/V1/V2/A2/M3/c1 ;
 wire \V1/V1/V2/A2/M3/c2 ;
 wire \V1/V1/V2/A2/M3/s1 ;
 wire \V1/V1/V2/A2/M4/c1 ;
 wire \V1/V1/V2/A2/M4/c2 ;
 wire \V1/V1/V2/A2/M4/s1 ;
 wire \V1/V1/V2/A3/c1 ;
 wire \V1/V1/V2/A3/c2 ;
 wire \V1/V1/V2/A3/c3 ;
 wire \V1/V1/V2/A3/M1/c1 ;
 wire \V1/V1/V2/A3/M1/c2 ;
 wire \V1/V1/V2/A3/M1/s1 ;
 wire \V1/V1/V2/A3/M2/c1 ;
 wire \V1/V1/V2/A3/M2/c2 ;
 wire \V1/V1/V2/A3/M2/s1 ;
 wire \V1/V1/V2/A3/M3/c1 ;
 wire \V1/V1/V2/A3/M3/c2 ;
 wire \V1/V1/V2/A3/M3/s1 ;
 wire \V1/V1/V2/A3/M4/c1 ;
 wire \V1/V1/V2/A3/M4/c2 ;
 wire \V1/V1/V2/A3/M4/s1 ;
 wire \V1/V1/V2/V1/w1 ;
 wire \V1/V1/V2/V1/w2 ;
 wire \V1/V1/V2/V1/w3 ;
 wire \V1/V1/V2/V1/w4 ;
 wire \V1/V1/V2/V2/w1 ;
 wire \V1/V1/V2/V2/w2 ;
 wire \V1/V1/V2/V2/w3 ;
 wire \V1/V1/V2/V2/w4 ;
 wire \V1/V1/V2/V3/w1 ;
 wire \V1/V1/V2/V3/w2 ;
 wire \V1/V1/V2/V3/w3 ;
 wire \V1/V1/V2/V3/w4 ;
 wire \V1/V1/V2/V4/w1 ;
 wire \V1/V1/V2/V4/w2 ;
 wire \V1/V1/V2/V4/w3 ;
 wire \V1/V1/V2/V4/w4 ;
 wire \V1/V1/V3/c1 ;
 wire \V1/V1/V3/c2 ;
 wire \V1/V1/V3/c3 ;
 wire \V1/V1/V3/overflow ;
 wire \V1/V1/V3/A1/c1 ;
 wire \V1/V1/V3/A1/c2 ;
 wire \V1/V1/V3/A1/c3 ;
 wire \V1/V1/V3/A1/M1/c1 ;
 wire \V1/V1/V3/A1/M1/c2 ;
 wire \V1/V1/V3/A1/M1/s1 ;
 wire \V1/V1/V3/A1/M2/c1 ;
 wire \V1/V1/V3/A1/M2/c2 ;
 wire \V1/V1/V3/A1/M2/s1 ;
 wire \V1/V1/V3/A1/M3/c1 ;
 wire \V1/V1/V3/A1/M3/c2 ;
 wire \V1/V1/V3/A1/M3/s1 ;
 wire \V1/V1/V3/A1/M4/c1 ;
 wire \V1/V1/V3/A1/M4/c2 ;
 wire \V1/V1/V3/A1/M4/s1 ;
 wire \V1/V1/V3/A2/c1 ;
 wire \V1/V1/V3/A2/c2 ;
 wire \V1/V1/V3/A2/c3 ;
 wire \V1/V1/V3/A2/M1/c1 ;
 wire \V1/V1/V3/A2/M1/c2 ;
 wire \V1/V1/V3/A2/M1/s1 ;
 wire \V1/V1/V3/A2/M2/c1 ;
 wire \V1/V1/V3/A2/M2/c2 ;
 wire \V1/V1/V3/A2/M2/s1 ;
 wire \V1/V1/V3/A2/M3/c1 ;
 wire \V1/V1/V3/A2/M3/c2 ;
 wire \V1/V1/V3/A2/M3/s1 ;
 wire \V1/V1/V3/A2/M4/c1 ;
 wire \V1/V1/V3/A2/M4/c2 ;
 wire \V1/V1/V3/A2/M4/s1 ;
 wire \V1/V1/V3/A3/c1 ;
 wire \V1/V1/V3/A3/c2 ;
 wire \V1/V1/V3/A3/c3 ;
 wire \V1/V1/V3/A3/M1/c1 ;
 wire \V1/V1/V3/A3/M1/c2 ;
 wire \V1/V1/V3/A3/M1/s1 ;
 wire \V1/V1/V3/A3/M2/c1 ;
 wire \V1/V1/V3/A3/M2/c2 ;
 wire \V1/V1/V3/A3/M2/s1 ;
 wire \V1/V1/V3/A3/M3/c1 ;
 wire \V1/V1/V3/A3/M3/c2 ;
 wire \V1/V1/V3/A3/M3/s1 ;
 wire \V1/V1/V3/A3/M4/c1 ;
 wire \V1/V1/V3/A3/M4/c2 ;
 wire \V1/V1/V3/A3/M4/s1 ;
 wire \V1/V1/V3/V1/w1 ;
 wire \V1/V1/V3/V1/w2 ;
 wire \V1/V1/V3/V1/w3 ;
 wire \V1/V1/V3/V1/w4 ;
 wire \V1/V1/V3/V2/w1 ;
 wire \V1/V1/V3/V2/w2 ;
 wire \V1/V1/V3/V2/w3 ;
 wire \V1/V1/V3/V2/w4 ;
 wire \V1/V1/V3/V3/w1 ;
 wire \V1/V1/V3/V3/w2 ;
 wire \V1/V1/V3/V3/w3 ;
 wire \V1/V1/V3/V3/w4 ;
 wire \V1/V1/V3/V4/w1 ;
 wire \V1/V1/V3/V4/w2 ;
 wire \V1/V1/V3/V4/w3 ;
 wire \V1/V1/V3/V4/w4 ;
 wire \V1/V1/V4/c1 ;
 wire \V1/V1/V4/c2 ;
 wire \V1/V1/V4/c3 ;
 wire \V1/V1/V4/overflow ;
 wire \V1/V1/V4/A1/c1 ;
 wire \V1/V1/V4/A1/c2 ;
 wire \V1/V1/V4/A1/c3 ;
 wire \V1/V1/V4/A1/M1/c1 ;
 wire \V1/V1/V4/A1/M1/c2 ;
 wire \V1/V1/V4/A1/M1/s1 ;
 wire \V1/V1/V4/A1/M2/c1 ;
 wire \V1/V1/V4/A1/M2/c2 ;
 wire \V1/V1/V4/A1/M2/s1 ;
 wire \V1/V1/V4/A1/M3/c1 ;
 wire \V1/V1/V4/A1/M3/c2 ;
 wire \V1/V1/V4/A1/M3/s1 ;
 wire \V1/V1/V4/A1/M4/c1 ;
 wire \V1/V1/V4/A1/M4/c2 ;
 wire \V1/V1/V4/A1/M4/s1 ;
 wire \V1/V1/V4/A2/c1 ;
 wire \V1/V1/V4/A2/c2 ;
 wire \V1/V1/V4/A2/c3 ;
 wire \V1/V1/V4/A2/M1/c1 ;
 wire \V1/V1/V4/A2/M1/c2 ;
 wire \V1/V1/V4/A2/M1/s1 ;
 wire \V1/V1/V4/A2/M2/c1 ;
 wire \V1/V1/V4/A2/M2/c2 ;
 wire \V1/V1/V4/A2/M2/s1 ;
 wire \V1/V1/V4/A2/M3/c1 ;
 wire \V1/V1/V4/A2/M3/c2 ;
 wire \V1/V1/V4/A2/M3/s1 ;
 wire \V1/V1/V4/A2/M4/c1 ;
 wire \V1/V1/V4/A2/M4/c2 ;
 wire \V1/V1/V4/A2/M4/s1 ;
 wire \V1/V1/V4/A3/c1 ;
 wire \V1/V1/V4/A3/c2 ;
 wire \V1/V1/V4/A3/c3 ;
 wire \V1/V1/V4/A3/M1/c1 ;
 wire \V1/V1/V4/A3/M1/c2 ;
 wire \V1/V1/V4/A3/M1/s1 ;
 wire \V1/V1/V4/A3/M2/c1 ;
 wire \V1/V1/V4/A3/M2/c2 ;
 wire \V1/V1/V4/A3/M2/s1 ;
 wire \V1/V1/V4/A3/M3/c1 ;
 wire \V1/V1/V4/A3/M3/c2 ;
 wire \V1/V1/V4/A3/M3/s1 ;
 wire \V1/V1/V4/A3/M4/c1 ;
 wire \V1/V1/V4/A3/M4/c2 ;
 wire \V1/V1/V4/A3/M4/s1 ;
 wire \V1/V1/V4/V1/w1 ;
 wire \V1/V1/V4/V1/w2 ;
 wire \V1/V1/V4/V1/w3 ;
 wire \V1/V1/V4/V1/w4 ;
 wire \V1/V1/V4/V2/w1 ;
 wire \V1/V1/V4/V2/w2 ;
 wire \V1/V1/V4/V2/w3 ;
 wire \V1/V1/V4/V2/w4 ;
 wire \V1/V1/V4/V3/w1 ;
 wire \V1/V1/V4/V3/w2 ;
 wire \V1/V1/V4/V3/w3 ;
 wire \V1/V1/V4/V3/w4 ;
 wire \V1/V1/V4/V4/w1 ;
 wire \V1/V1/V4/V4/w2 ;
 wire \V1/V1/V4/V4/w3 ;
 wire \V1/V1/V4/V4/w4 ;
 wire \V1/V2/c1 ;
 wire \V1/V2/c2 ;
 wire \V1/V2/c3 ;
 wire \V1/V2/overflow ;
 wire \V1/V2/A1/c1 ;
 wire \V1/V2/A1/A1/c1 ;
 wire \V1/V2/A1/A1/c2 ;
 wire \V1/V2/A1/A1/c3 ;
 wire \V1/V2/A1/A1/M1/c1 ;
 wire \V1/V2/A1/A1/M1/c2 ;
 wire \V1/V2/A1/A1/M1/s1 ;
 wire \V1/V2/A1/A1/M2/c1 ;
 wire \V1/V2/A1/A1/M2/c2 ;
 wire \V1/V2/A1/A1/M2/s1 ;
 wire \V1/V2/A1/A1/M3/c1 ;
 wire \V1/V2/A1/A1/M3/c2 ;
 wire \V1/V2/A1/A1/M3/s1 ;
 wire \V1/V2/A1/A1/M4/c1 ;
 wire \V1/V2/A1/A1/M4/c2 ;
 wire \V1/V2/A1/A1/M4/s1 ;
 wire \V1/V2/A1/A2/c1 ;
 wire \V1/V2/A1/A2/c2 ;
 wire \V1/V2/A1/A2/c3 ;
 wire \V1/V2/A1/A2/M1/c1 ;
 wire \V1/V2/A1/A2/M1/c2 ;
 wire \V1/V2/A1/A2/M1/s1 ;
 wire \V1/V2/A1/A2/M2/c1 ;
 wire \V1/V2/A1/A2/M2/c2 ;
 wire \V1/V2/A1/A2/M2/s1 ;
 wire \V1/V2/A1/A2/M3/c1 ;
 wire \V1/V2/A1/A2/M3/c2 ;
 wire \V1/V2/A1/A2/M3/s1 ;
 wire \V1/V2/A1/A2/M4/c1 ;
 wire \V1/V2/A1/A2/M4/c2 ;
 wire \V1/V2/A1/A2/M4/s1 ;
 wire \V1/V2/A2/c1 ;
 wire \V1/V2/A2/A1/c1 ;
 wire \V1/V2/A2/A1/c2 ;
 wire \V1/V2/A2/A1/c3 ;
 wire \V1/V2/A2/A1/M1/c1 ;
 wire \V1/V2/A2/A1/M1/c2 ;
 wire \V1/V2/A2/A1/M1/s1 ;
 wire \V1/V2/A2/A1/M2/c1 ;
 wire \V1/V2/A2/A1/M2/c2 ;
 wire \V1/V2/A2/A1/M2/s1 ;
 wire \V1/V2/A2/A1/M3/c1 ;
 wire \V1/V2/A2/A1/M3/c2 ;
 wire \V1/V2/A2/A1/M3/s1 ;
 wire \V1/V2/A2/A1/M4/c1 ;
 wire \V1/V2/A2/A1/M4/c2 ;
 wire \V1/V2/A2/A1/M4/s1 ;
 wire \V1/V2/A2/A2/c1 ;
 wire \V1/V2/A2/A2/c2 ;
 wire \V1/V2/A2/A2/c3 ;
 wire \V1/V2/A2/A2/M1/c1 ;
 wire \V1/V2/A2/A2/M1/c2 ;
 wire \V1/V2/A2/A2/M1/s1 ;
 wire \V1/V2/A2/A2/M2/c1 ;
 wire \V1/V2/A2/A2/M2/c2 ;
 wire \V1/V2/A2/A2/M2/s1 ;
 wire \V1/V2/A2/A2/M3/c1 ;
 wire \V1/V2/A2/A2/M3/c2 ;
 wire \V1/V2/A2/A2/M3/s1 ;
 wire \V1/V2/A2/A2/M4/c1 ;
 wire \V1/V2/A2/A2/M4/c2 ;
 wire \V1/V2/A2/A2/M4/s1 ;
 wire \V1/V2/A3/c1 ;
 wire \V1/V2/A3/A1/c1 ;
 wire \V1/V2/A3/A1/c2 ;
 wire \V1/V2/A3/A1/c3 ;
 wire \V1/V2/A3/A1/M1/c1 ;
 wire \V1/V2/A3/A1/M1/c2 ;
 wire \V1/V2/A3/A1/M1/s1 ;
 wire \V1/V2/A3/A1/M2/c1 ;
 wire \V1/V2/A3/A1/M2/c2 ;
 wire \V1/V2/A3/A1/M2/s1 ;
 wire \V1/V2/A3/A1/M3/c1 ;
 wire \V1/V2/A3/A1/M3/c2 ;
 wire \V1/V2/A3/A1/M3/s1 ;
 wire \V1/V2/A3/A1/M4/c1 ;
 wire \V1/V2/A3/A1/M4/c2 ;
 wire \V1/V2/A3/A1/M4/s1 ;
 wire \V1/V2/A3/A2/c1 ;
 wire \V1/V2/A3/A2/c2 ;
 wire \V1/V2/A3/A2/c3 ;
 wire \V1/V2/A3/A2/M1/c1 ;
 wire \V1/V2/A3/A2/M1/c2 ;
 wire \V1/V2/A3/A2/M1/s1 ;
 wire \V1/V2/A3/A2/M2/c1 ;
 wire \V1/V2/A3/A2/M2/c2 ;
 wire \V1/V2/A3/A2/M2/s1 ;
 wire \V1/V2/A3/A2/M3/c1 ;
 wire \V1/V2/A3/A2/M3/c2 ;
 wire \V1/V2/A3/A2/M3/s1 ;
 wire \V1/V2/A3/A2/M4/c1 ;
 wire \V1/V2/A3/A2/M4/c2 ;
 wire \V1/V2/A3/A2/M4/s1 ;
 wire \V1/V2/V1/c1 ;
 wire \V1/V2/V1/c2 ;
 wire \V1/V2/V1/c3 ;
 wire \V1/V2/V1/overflow ;
 wire \V1/V2/V1/A1/c1 ;
 wire \V1/V2/V1/A1/c2 ;
 wire \V1/V2/V1/A1/c3 ;
 wire \V1/V2/V1/A1/M1/c1 ;
 wire \V1/V2/V1/A1/M1/c2 ;
 wire \V1/V2/V1/A1/M1/s1 ;
 wire \V1/V2/V1/A1/M2/c1 ;
 wire \V1/V2/V1/A1/M2/c2 ;
 wire \V1/V2/V1/A1/M2/s1 ;
 wire \V1/V2/V1/A1/M3/c1 ;
 wire \V1/V2/V1/A1/M3/c2 ;
 wire \V1/V2/V1/A1/M3/s1 ;
 wire \V1/V2/V1/A1/M4/c1 ;
 wire \V1/V2/V1/A1/M4/c2 ;
 wire \V1/V2/V1/A1/M4/s1 ;
 wire \V1/V2/V1/A2/c1 ;
 wire \V1/V2/V1/A2/c2 ;
 wire \V1/V2/V1/A2/c3 ;
 wire \V1/V2/V1/A2/M1/c1 ;
 wire \V1/V2/V1/A2/M1/c2 ;
 wire \V1/V2/V1/A2/M1/s1 ;
 wire \V1/V2/V1/A2/M2/c1 ;
 wire \V1/V2/V1/A2/M2/c2 ;
 wire \V1/V2/V1/A2/M2/s1 ;
 wire \V1/V2/V1/A2/M3/c1 ;
 wire \V1/V2/V1/A2/M3/c2 ;
 wire \V1/V2/V1/A2/M3/s1 ;
 wire \V1/V2/V1/A2/M4/c1 ;
 wire \V1/V2/V1/A2/M4/c2 ;
 wire \V1/V2/V1/A2/M4/s1 ;
 wire \V1/V2/V1/A3/c1 ;
 wire \V1/V2/V1/A3/c2 ;
 wire \V1/V2/V1/A3/c3 ;
 wire \V1/V2/V1/A3/M1/c1 ;
 wire \V1/V2/V1/A3/M1/c2 ;
 wire \V1/V2/V1/A3/M1/s1 ;
 wire \V1/V2/V1/A3/M2/c1 ;
 wire \V1/V2/V1/A3/M2/c2 ;
 wire \V1/V2/V1/A3/M2/s1 ;
 wire \V1/V2/V1/A3/M3/c1 ;
 wire \V1/V2/V1/A3/M3/c2 ;
 wire \V1/V2/V1/A3/M3/s1 ;
 wire \V1/V2/V1/A3/M4/c1 ;
 wire \V1/V2/V1/A3/M4/c2 ;
 wire \V1/V2/V1/A3/M4/s1 ;
 wire \V1/V2/V1/V1/w1 ;
 wire \V1/V2/V1/V1/w2 ;
 wire \V1/V2/V1/V1/w3 ;
 wire \V1/V2/V1/V1/w4 ;
 wire \V1/V2/V1/V2/w1 ;
 wire \V1/V2/V1/V2/w2 ;
 wire \V1/V2/V1/V2/w3 ;
 wire \V1/V2/V1/V2/w4 ;
 wire \V1/V2/V1/V3/w1 ;
 wire \V1/V2/V1/V3/w2 ;
 wire \V1/V2/V1/V3/w3 ;
 wire \V1/V2/V1/V3/w4 ;
 wire \V1/V2/V1/V4/w1 ;
 wire \V1/V2/V1/V4/w2 ;
 wire \V1/V2/V1/V4/w3 ;
 wire \V1/V2/V1/V4/w4 ;
 wire \V1/V2/V2/c1 ;
 wire \V1/V2/V2/c2 ;
 wire \V1/V2/V2/c3 ;
 wire \V1/V2/V2/overflow ;
 wire \V1/V2/V2/A1/c1 ;
 wire \V1/V2/V2/A1/c2 ;
 wire \V1/V2/V2/A1/c3 ;
 wire \V1/V2/V2/A1/M1/c1 ;
 wire \V1/V2/V2/A1/M1/c2 ;
 wire \V1/V2/V2/A1/M1/s1 ;
 wire \V1/V2/V2/A1/M2/c1 ;
 wire \V1/V2/V2/A1/M2/c2 ;
 wire \V1/V2/V2/A1/M2/s1 ;
 wire \V1/V2/V2/A1/M3/c1 ;
 wire \V1/V2/V2/A1/M3/c2 ;
 wire \V1/V2/V2/A1/M3/s1 ;
 wire \V1/V2/V2/A1/M4/c1 ;
 wire \V1/V2/V2/A1/M4/c2 ;
 wire \V1/V2/V2/A1/M4/s1 ;
 wire \V1/V2/V2/A2/c1 ;
 wire \V1/V2/V2/A2/c2 ;
 wire \V1/V2/V2/A2/c3 ;
 wire \V1/V2/V2/A2/M1/c1 ;
 wire \V1/V2/V2/A2/M1/c2 ;
 wire \V1/V2/V2/A2/M1/s1 ;
 wire \V1/V2/V2/A2/M2/c1 ;
 wire \V1/V2/V2/A2/M2/c2 ;
 wire \V1/V2/V2/A2/M2/s1 ;
 wire \V1/V2/V2/A2/M3/c1 ;
 wire \V1/V2/V2/A2/M3/c2 ;
 wire \V1/V2/V2/A2/M3/s1 ;
 wire \V1/V2/V2/A2/M4/c1 ;
 wire \V1/V2/V2/A2/M4/c2 ;
 wire \V1/V2/V2/A2/M4/s1 ;
 wire \V1/V2/V2/A3/c1 ;
 wire \V1/V2/V2/A3/c2 ;
 wire \V1/V2/V2/A3/c3 ;
 wire \V1/V2/V2/A3/M1/c1 ;
 wire \V1/V2/V2/A3/M1/c2 ;
 wire \V1/V2/V2/A3/M1/s1 ;
 wire \V1/V2/V2/A3/M2/c1 ;
 wire \V1/V2/V2/A3/M2/c2 ;
 wire \V1/V2/V2/A3/M2/s1 ;
 wire \V1/V2/V2/A3/M3/c1 ;
 wire \V1/V2/V2/A3/M3/c2 ;
 wire \V1/V2/V2/A3/M3/s1 ;
 wire \V1/V2/V2/A3/M4/c1 ;
 wire \V1/V2/V2/A3/M4/c2 ;
 wire \V1/V2/V2/A3/M4/s1 ;
 wire \V1/V2/V2/V1/w1 ;
 wire \V1/V2/V2/V1/w2 ;
 wire \V1/V2/V2/V1/w3 ;
 wire \V1/V2/V2/V1/w4 ;
 wire \V1/V2/V2/V2/w1 ;
 wire \V1/V2/V2/V2/w2 ;
 wire \V1/V2/V2/V2/w3 ;
 wire \V1/V2/V2/V2/w4 ;
 wire \V1/V2/V2/V3/w1 ;
 wire \V1/V2/V2/V3/w2 ;
 wire \V1/V2/V2/V3/w3 ;
 wire \V1/V2/V2/V3/w4 ;
 wire \V1/V2/V2/V4/w1 ;
 wire \V1/V2/V2/V4/w2 ;
 wire \V1/V2/V2/V4/w3 ;
 wire \V1/V2/V2/V4/w4 ;
 wire \V1/V2/V3/c1 ;
 wire \V1/V2/V3/c2 ;
 wire \V1/V2/V3/c3 ;
 wire \V1/V2/V3/overflow ;
 wire \V1/V2/V3/A1/c1 ;
 wire \V1/V2/V3/A1/c2 ;
 wire \V1/V2/V3/A1/c3 ;
 wire \V1/V2/V3/A1/M1/c1 ;
 wire \V1/V2/V3/A1/M1/c2 ;
 wire \V1/V2/V3/A1/M1/s1 ;
 wire \V1/V2/V3/A1/M2/c1 ;
 wire \V1/V2/V3/A1/M2/c2 ;
 wire \V1/V2/V3/A1/M2/s1 ;
 wire \V1/V2/V3/A1/M3/c1 ;
 wire \V1/V2/V3/A1/M3/c2 ;
 wire \V1/V2/V3/A1/M3/s1 ;
 wire \V1/V2/V3/A1/M4/c1 ;
 wire \V1/V2/V3/A1/M4/c2 ;
 wire \V1/V2/V3/A1/M4/s1 ;
 wire \V1/V2/V3/A2/c1 ;
 wire \V1/V2/V3/A2/c2 ;
 wire \V1/V2/V3/A2/c3 ;
 wire \V1/V2/V3/A2/M1/c1 ;
 wire \V1/V2/V3/A2/M1/c2 ;
 wire \V1/V2/V3/A2/M1/s1 ;
 wire \V1/V2/V3/A2/M2/c1 ;
 wire \V1/V2/V3/A2/M2/c2 ;
 wire \V1/V2/V3/A2/M2/s1 ;
 wire \V1/V2/V3/A2/M3/c1 ;
 wire \V1/V2/V3/A2/M3/c2 ;
 wire \V1/V2/V3/A2/M3/s1 ;
 wire \V1/V2/V3/A2/M4/c1 ;
 wire \V1/V2/V3/A2/M4/c2 ;
 wire \V1/V2/V3/A2/M4/s1 ;
 wire \V1/V2/V3/A3/c1 ;
 wire \V1/V2/V3/A3/c2 ;
 wire \V1/V2/V3/A3/c3 ;
 wire \V1/V2/V3/A3/M1/c1 ;
 wire \V1/V2/V3/A3/M1/c2 ;
 wire \V1/V2/V3/A3/M1/s1 ;
 wire \V1/V2/V3/A3/M2/c1 ;
 wire \V1/V2/V3/A3/M2/c2 ;
 wire \V1/V2/V3/A3/M2/s1 ;
 wire \V1/V2/V3/A3/M3/c1 ;
 wire \V1/V2/V3/A3/M3/c2 ;
 wire \V1/V2/V3/A3/M3/s1 ;
 wire \V1/V2/V3/A3/M4/c1 ;
 wire \V1/V2/V3/A3/M4/c2 ;
 wire \V1/V2/V3/A3/M4/s1 ;
 wire \V1/V2/V3/V1/w1 ;
 wire \V1/V2/V3/V1/w2 ;
 wire \V1/V2/V3/V1/w3 ;
 wire \V1/V2/V3/V1/w4 ;
 wire \V1/V2/V3/V2/w1 ;
 wire \V1/V2/V3/V2/w2 ;
 wire \V1/V2/V3/V2/w3 ;
 wire \V1/V2/V3/V2/w4 ;
 wire \V1/V2/V3/V3/w1 ;
 wire \V1/V2/V3/V3/w2 ;
 wire \V1/V2/V3/V3/w3 ;
 wire \V1/V2/V3/V3/w4 ;
 wire \V1/V2/V3/V4/w1 ;
 wire \V1/V2/V3/V4/w2 ;
 wire \V1/V2/V3/V4/w3 ;
 wire \V1/V2/V3/V4/w4 ;
 wire \V1/V2/V4/c1 ;
 wire \V1/V2/V4/c2 ;
 wire \V1/V2/V4/c3 ;
 wire \V1/V2/V4/overflow ;
 wire \V1/V2/V4/A1/c1 ;
 wire \V1/V2/V4/A1/c2 ;
 wire \V1/V2/V4/A1/c3 ;
 wire \V1/V2/V4/A1/M1/c1 ;
 wire \V1/V2/V4/A1/M1/c2 ;
 wire \V1/V2/V4/A1/M1/s1 ;
 wire \V1/V2/V4/A1/M2/c1 ;
 wire \V1/V2/V4/A1/M2/c2 ;
 wire \V1/V2/V4/A1/M2/s1 ;
 wire \V1/V2/V4/A1/M3/c1 ;
 wire \V1/V2/V4/A1/M3/c2 ;
 wire \V1/V2/V4/A1/M3/s1 ;
 wire \V1/V2/V4/A1/M4/c1 ;
 wire \V1/V2/V4/A1/M4/c2 ;
 wire \V1/V2/V4/A1/M4/s1 ;
 wire \V1/V2/V4/A2/c1 ;
 wire \V1/V2/V4/A2/c2 ;
 wire \V1/V2/V4/A2/c3 ;
 wire \V1/V2/V4/A2/M1/c1 ;
 wire \V1/V2/V4/A2/M1/c2 ;
 wire \V1/V2/V4/A2/M1/s1 ;
 wire \V1/V2/V4/A2/M2/c1 ;
 wire \V1/V2/V4/A2/M2/c2 ;
 wire \V1/V2/V4/A2/M2/s1 ;
 wire \V1/V2/V4/A2/M3/c1 ;
 wire \V1/V2/V4/A2/M3/c2 ;
 wire \V1/V2/V4/A2/M3/s1 ;
 wire \V1/V2/V4/A2/M4/c1 ;
 wire \V1/V2/V4/A2/M4/c2 ;
 wire \V1/V2/V4/A2/M4/s1 ;
 wire \V1/V2/V4/A3/c1 ;
 wire \V1/V2/V4/A3/c2 ;
 wire \V1/V2/V4/A3/c3 ;
 wire \V1/V2/V4/A3/M1/c1 ;
 wire \V1/V2/V4/A3/M1/c2 ;
 wire \V1/V2/V4/A3/M1/s1 ;
 wire \V1/V2/V4/A3/M2/c1 ;
 wire \V1/V2/V4/A3/M2/c2 ;
 wire \V1/V2/V4/A3/M2/s1 ;
 wire \V1/V2/V4/A3/M3/c1 ;
 wire \V1/V2/V4/A3/M3/c2 ;
 wire \V1/V2/V4/A3/M3/s1 ;
 wire \V1/V2/V4/A3/M4/c1 ;
 wire \V1/V2/V4/A3/M4/c2 ;
 wire \V1/V2/V4/A3/M4/s1 ;
 wire \V1/V2/V4/V1/w1 ;
 wire \V1/V2/V4/V1/w2 ;
 wire \V1/V2/V4/V1/w3 ;
 wire \V1/V2/V4/V1/w4 ;
 wire \V1/V2/V4/V2/w1 ;
 wire \V1/V2/V4/V2/w2 ;
 wire \V1/V2/V4/V2/w3 ;
 wire \V1/V2/V4/V2/w4 ;
 wire \V1/V2/V4/V3/w1 ;
 wire \V1/V2/V4/V3/w2 ;
 wire \V1/V2/V4/V3/w3 ;
 wire \V1/V2/V4/V3/w4 ;
 wire \V1/V2/V4/V4/w1 ;
 wire \V1/V2/V4/V4/w2 ;
 wire \V1/V2/V4/V4/w3 ;
 wire \V1/V2/V4/V4/w4 ;
 wire \V1/V3/c1 ;
 wire \V1/V3/c2 ;
 wire \V1/V3/c3 ;
 wire \V1/V3/overflow ;
 wire \V1/V3/A1/c1 ;
 wire \V1/V3/A1/A1/c1 ;
 wire \V1/V3/A1/A1/c2 ;
 wire \V1/V3/A1/A1/c3 ;
 wire \V1/V3/A1/A1/M1/c1 ;
 wire \V1/V3/A1/A1/M1/c2 ;
 wire \V1/V3/A1/A1/M1/s1 ;
 wire \V1/V3/A1/A1/M2/c1 ;
 wire \V1/V3/A1/A1/M2/c2 ;
 wire \V1/V3/A1/A1/M2/s1 ;
 wire \V1/V3/A1/A1/M3/c1 ;
 wire \V1/V3/A1/A1/M3/c2 ;
 wire \V1/V3/A1/A1/M3/s1 ;
 wire \V1/V3/A1/A1/M4/c1 ;
 wire \V1/V3/A1/A1/M4/c2 ;
 wire \V1/V3/A1/A1/M4/s1 ;
 wire \V1/V3/A1/A2/c1 ;
 wire \V1/V3/A1/A2/c2 ;
 wire \V1/V3/A1/A2/c3 ;
 wire \V1/V3/A1/A2/M1/c1 ;
 wire \V1/V3/A1/A2/M1/c2 ;
 wire \V1/V3/A1/A2/M1/s1 ;
 wire \V1/V3/A1/A2/M2/c1 ;
 wire \V1/V3/A1/A2/M2/c2 ;
 wire \V1/V3/A1/A2/M2/s1 ;
 wire \V1/V3/A1/A2/M3/c1 ;
 wire \V1/V3/A1/A2/M3/c2 ;
 wire \V1/V3/A1/A2/M3/s1 ;
 wire \V1/V3/A1/A2/M4/c1 ;
 wire \V1/V3/A1/A2/M4/c2 ;
 wire \V1/V3/A1/A2/M4/s1 ;
 wire \V1/V3/A2/c1 ;
 wire \V1/V3/A2/A1/c1 ;
 wire \V1/V3/A2/A1/c2 ;
 wire \V1/V3/A2/A1/c3 ;
 wire \V1/V3/A2/A1/M1/c1 ;
 wire \V1/V3/A2/A1/M1/c2 ;
 wire \V1/V3/A2/A1/M1/s1 ;
 wire \V1/V3/A2/A1/M2/c1 ;
 wire \V1/V3/A2/A1/M2/c2 ;
 wire \V1/V3/A2/A1/M2/s1 ;
 wire \V1/V3/A2/A1/M3/c1 ;
 wire \V1/V3/A2/A1/M3/c2 ;
 wire \V1/V3/A2/A1/M3/s1 ;
 wire \V1/V3/A2/A1/M4/c1 ;
 wire \V1/V3/A2/A1/M4/c2 ;
 wire \V1/V3/A2/A1/M4/s1 ;
 wire \V1/V3/A2/A2/c1 ;
 wire \V1/V3/A2/A2/c2 ;
 wire \V1/V3/A2/A2/c3 ;
 wire \V1/V3/A2/A2/M1/c1 ;
 wire \V1/V3/A2/A2/M1/c2 ;
 wire \V1/V3/A2/A2/M1/s1 ;
 wire \V1/V3/A2/A2/M2/c1 ;
 wire \V1/V3/A2/A2/M2/c2 ;
 wire \V1/V3/A2/A2/M2/s1 ;
 wire \V1/V3/A2/A2/M3/c1 ;
 wire \V1/V3/A2/A2/M3/c2 ;
 wire \V1/V3/A2/A2/M3/s1 ;
 wire \V1/V3/A2/A2/M4/c1 ;
 wire \V1/V3/A2/A2/M4/c2 ;
 wire \V1/V3/A2/A2/M4/s1 ;
 wire \V1/V3/A3/c1 ;
 wire \V1/V3/A3/A1/c1 ;
 wire \V1/V3/A3/A1/c2 ;
 wire \V1/V3/A3/A1/c3 ;
 wire \V1/V3/A3/A1/M1/c1 ;
 wire \V1/V3/A3/A1/M1/c2 ;
 wire \V1/V3/A3/A1/M1/s1 ;
 wire \V1/V3/A3/A1/M2/c1 ;
 wire \V1/V3/A3/A1/M2/c2 ;
 wire \V1/V3/A3/A1/M2/s1 ;
 wire \V1/V3/A3/A1/M3/c1 ;
 wire \V1/V3/A3/A1/M3/c2 ;
 wire \V1/V3/A3/A1/M3/s1 ;
 wire \V1/V3/A3/A1/M4/c1 ;
 wire \V1/V3/A3/A1/M4/c2 ;
 wire \V1/V3/A3/A1/M4/s1 ;
 wire \V1/V3/A3/A2/c1 ;
 wire \V1/V3/A3/A2/c2 ;
 wire \V1/V3/A3/A2/c3 ;
 wire \V1/V3/A3/A2/M1/c1 ;
 wire \V1/V3/A3/A2/M1/c2 ;
 wire \V1/V3/A3/A2/M1/s1 ;
 wire \V1/V3/A3/A2/M2/c1 ;
 wire \V1/V3/A3/A2/M2/c2 ;
 wire \V1/V3/A3/A2/M2/s1 ;
 wire \V1/V3/A3/A2/M3/c1 ;
 wire \V1/V3/A3/A2/M3/c2 ;
 wire \V1/V3/A3/A2/M3/s1 ;
 wire \V1/V3/A3/A2/M4/c1 ;
 wire \V1/V3/A3/A2/M4/c2 ;
 wire \V1/V3/A3/A2/M4/s1 ;
 wire \V1/V3/V1/c1 ;
 wire \V1/V3/V1/c2 ;
 wire \V1/V3/V1/c3 ;
 wire \V1/V3/V1/overflow ;
 wire \V1/V3/V1/A1/c1 ;
 wire \V1/V3/V1/A1/c2 ;
 wire \V1/V3/V1/A1/c3 ;
 wire \V1/V3/V1/A1/M1/c1 ;
 wire \V1/V3/V1/A1/M1/c2 ;
 wire \V1/V3/V1/A1/M1/s1 ;
 wire \V1/V3/V1/A1/M2/c1 ;
 wire \V1/V3/V1/A1/M2/c2 ;
 wire \V1/V3/V1/A1/M2/s1 ;
 wire \V1/V3/V1/A1/M3/c1 ;
 wire \V1/V3/V1/A1/M3/c2 ;
 wire \V1/V3/V1/A1/M3/s1 ;
 wire \V1/V3/V1/A1/M4/c1 ;
 wire \V1/V3/V1/A1/M4/c2 ;
 wire \V1/V3/V1/A1/M4/s1 ;
 wire \V1/V3/V1/A2/c1 ;
 wire \V1/V3/V1/A2/c2 ;
 wire \V1/V3/V1/A2/c3 ;
 wire \V1/V3/V1/A2/M1/c1 ;
 wire \V1/V3/V1/A2/M1/c2 ;
 wire \V1/V3/V1/A2/M1/s1 ;
 wire \V1/V3/V1/A2/M2/c1 ;
 wire \V1/V3/V1/A2/M2/c2 ;
 wire \V1/V3/V1/A2/M2/s1 ;
 wire \V1/V3/V1/A2/M3/c1 ;
 wire \V1/V3/V1/A2/M3/c2 ;
 wire \V1/V3/V1/A2/M3/s1 ;
 wire \V1/V3/V1/A2/M4/c1 ;
 wire \V1/V3/V1/A2/M4/c2 ;
 wire \V1/V3/V1/A2/M4/s1 ;
 wire \V1/V3/V1/A3/c1 ;
 wire \V1/V3/V1/A3/c2 ;
 wire \V1/V3/V1/A3/c3 ;
 wire \V1/V3/V1/A3/M1/c1 ;
 wire \V1/V3/V1/A3/M1/c2 ;
 wire \V1/V3/V1/A3/M1/s1 ;
 wire \V1/V3/V1/A3/M2/c1 ;
 wire \V1/V3/V1/A3/M2/c2 ;
 wire \V1/V3/V1/A3/M2/s1 ;
 wire \V1/V3/V1/A3/M3/c1 ;
 wire \V1/V3/V1/A3/M3/c2 ;
 wire \V1/V3/V1/A3/M3/s1 ;
 wire \V1/V3/V1/A3/M4/c1 ;
 wire \V1/V3/V1/A3/M4/c2 ;
 wire \V1/V3/V1/A3/M4/s1 ;
 wire \V1/V3/V1/V1/w1 ;
 wire \V1/V3/V1/V1/w2 ;
 wire \V1/V3/V1/V1/w3 ;
 wire \V1/V3/V1/V1/w4 ;
 wire \V1/V3/V1/V2/w1 ;
 wire \V1/V3/V1/V2/w2 ;
 wire \V1/V3/V1/V2/w3 ;
 wire \V1/V3/V1/V2/w4 ;
 wire \V1/V3/V1/V3/w1 ;
 wire \V1/V3/V1/V3/w2 ;
 wire \V1/V3/V1/V3/w3 ;
 wire \V1/V3/V1/V3/w4 ;
 wire \V1/V3/V1/V4/w1 ;
 wire \V1/V3/V1/V4/w2 ;
 wire \V1/V3/V1/V4/w3 ;
 wire \V1/V3/V1/V4/w4 ;
 wire \V1/V3/V2/c1 ;
 wire \V1/V3/V2/c2 ;
 wire \V1/V3/V2/c3 ;
 wire \V1/V3/V2/overflow ;
 wire \V1/V3/V2/A1/c1 ;
 wire \V1/V3/V2/A1/c2 ;
 wire \V1/V3/V2/A1/c3 ;
 wire \V1/V3/V2/A1/M1/c1 ;
 wire \V1/V3/V2/A1/M1/c2 ;
 wire \V1/V3/V2/A1/M1/s1 ;
 wire \V1/V3/V2/A1/M2/c1 ;
 wire \V1/V3/V2/A1/M2/c2 ;
 wire \V1/V3/V2/A1/M2/s1 ;
 wire \V1/V3/V2/A1/M3/c1 ;
 wire \V1/V3/V2/A1/M3/c2 ;
 wire \V1/V3/V2/A1/M3/s1 ;
 wire \V1/V3/V2/A1/M4/c1 ;
 wire \V1/V3/V2/A1/M4/c2 ;
 wire \V1/V3/V2/A1/M4/s1 ;
 wire \V1/V3/V2/A2/c1 ;
 wire \V1/V3/V2/A2/c2 ;
 wire \V1/V3/V2/A2/c3 ;
 wire \V1/V3/V2/A2/M1/c1 ;
 wire \V1/V3/V2/A2/M1/c2 ;
 wire \V1/V3/V2/A2/M1/s1 ;
 wire \V1/V3/V2/A2/M2/c1 ;
 wire \V1/V3/V2/A2/M2/c2 ;
 wire \V1/V3/V2/A2/M2/s1 ;
 wire \V1/V3/V2/A2/M3/c1 ;
 wire \V1/V3/V2/A2/M3/c2 ;
 wire \V1/V3/V2/A2/M3/s1 ;
 wire \V1/V3/V2/A2/M4/c1 ;
 wire \V1/V3/V2/A2/M4/c2 ;
 wire \V1/V3/V2/A2/M4/s1 ;
 wire \V1/V3/V2/A3/c1 ;
 wire \V1/V3/V2/A3/c2 ;
 wire \V1/V3/V2/A3/c3 ;
 wire \V1/V3/V2/A3/M1/c1 ;
 wire \V1/V3/V2/A3/M1/c2 ;
 wire \V1/V3/V2/A3/M1/s1 ;
 wire \V1/V3/V2/A3/M2/c1 ;
 wire \V1/V3/V2/A3/M2/c2 ;
 wire \V1/V3/V2/A3/M2/s1 ;
 wire \V1/V3/V2/A3/M3/c1 ;
 wire \V1/V3/V2/A3/M3/c2 ;
 wire \V1/V3/V2/A3/M3/s1 ;
 wire \V1/V3/V2/A3/M4/c1 ;
 wire \V1/V3/V2/A3/M4/c2 ;
 wire \V1/V3/V2/A3/M4/s1 ;
 wire \V1/V3/V2/V1/w1 ;
 wire \V1/V3/V2/V1/w2 ;
 wire \V1/V3/V2/V1/w3 ;
 wire \V1/V3/V2/V1/w4 ;
 wire \V1/V3/V2/V2/w1 ;
 wire \V1/V3/V2/V2/w2 ;
 wire \V1/V3/V2/V2/w3 ;
 wire \V1/V3/V2/V2/w4 ;
 wire \V1/V3/V2/V3/w1 ;
 wire \V1/V3/V2/V3/w2 ;
 wire \V1/V3/V2/V3/w3 ;
 wire \V1/V3/V2/V3/w4 ;
 wire \V1/V3/V2/V4/w1 ;
 wire \V1/V3/V2/V4/w2 ;
 wire \V1/V3/V2/V4/w3 ;
 wire \V1/V3/V2/V4/w4 ;
 wire \V1/V3/V3/c1 ;
 wire \V1/V3/V3/c2 ;
 wire \V1/V3/V3/c3 ;
 wire \V1/V3/V3/overflow ;
 wire \V1/V3/V3/A1/c1 ;
 wire \V1/V3/V3/A1/c2 ;
 wire \V1/V3/V3/A1/c3 ;
 wire \V1/V3/V3/A1/M1/c1 ;
 wire \V1/V3/V3/A1/M1/c2 ;
 wire \V1/V3/V3/A1/M1/s1 ;
 wire \V1/V3/V3/A1/M2/c1 ;
 wire \V1/V3/V3/A1/M2/c2 ;
 wire \V1/V3/V3/A1/M2/s1 ;
 wire \V1/V3/V3/A1/M3/c1 ;
 wire \V1/V3/V3/A1/M3/c2 ;
 wire \V1/V3/V3/A1/M3/s1 ;
 wire \V1/V3/V3/A1/M4/c1 ;
 wire \V1/V3/V3/A1/M4/c2 ;
 wire \V1/V3/V3/A1/M4/s1 ;
 wire \V1/V3/V3/A2/c1 ;
 wire \V1/V3/V3/A2/c2 ;
 wire \V1/V3/V3/A2/c3 ;
 wire \V1/V3/V3/A2/M1/c1 ;
 wire \V1/V3/V3/A2/M1/c2 ;
 wire \V1/V3/V3/A2/M1/s1 ;
 wire \V1/V3/V3/A2/M2/c1 ;
 wire \V1/V3/V3/A2/M2/c2 ;
 wire \V1/V3/V3/A2/M2/s1 ;
 wire \V1/V3/V3/A2/M3/c1 ;
 wire \V1/V3/V3/A2/M3/c2 ;
 wire \V1/V3/V3/A2/M3/s1 ;
 wire \V1/V3/V3/A2/M4/c1 ;
 wire \V1/V3/V3/A2/M4/c2 ;
 wire \V1/V3/V3/A2/M4/s1 ;
 wire \V1/V3/V3/A3/c1 ;
 wire \V1/V3/V3/A3/c2 ;
 wire \V1/V3/V3/A3/c3 ;
 wire \V1/V3/V3/A3/M1/c1 ;
 wire \V1/V3/V3/A3/M1/c2 ;
 wire \V1/V3/V3/A3/M1/s1 ;
 wire \V1/V3/V3/A3/M2/c1 ;
 wire \V1/V3/V3/A3/M2/c2 ;
 wire \V1/V3/V3/A3/M2/s1 ;
 wire \V1/V3/V3/A3/M3/c1 ;
 wire \V1/V3/V3/A3/M3/c2 ;
 wire \V1/V3/V3/A3/M3/s1 ;
 wire \V1/V3/V3/A3/M4/c1 ;
 wire \V1/V3/V3/A3/M4/c2 ;
 wire \V1/V3/V3/A3/M4/s1 ;
 wire \V1/V3/V3/V1/w1 ;
 wire \V1/V3/V3/V1/w2 ;
 wire \V1/V3/V3/V1/w3 ;
 wire \V1/V3/V3/V1/w4 ;
 wire \V1/V3/V3/V2/w1 ;
 wire \V1/V3/V3/V2/w2 ;
 wire \V1/V3/V3/V2/w3 ;
 wire \V1/V3/V3/V2/w4 ;
 wire \V1/V3/V3/V3/w1 ;
 wire \V1/V3/V3/V3/w2 ;
 wire \V1/V3/V3/V3/w3 ;
 wire \V1/V3/V3/V3/w4 ;
 wire \V1/V3/V3/V4/w1 ;
 wire \V1/V3/V3/V4/w2 ;
 wire \V1/V3/V3/V4/w3 ;
 wire \V1/V3/V3/V4/w4 ;
 wire \V1/V3/V4/c1 ;
 wire \V1/V3/V4/c2 ;
 wire \V1/V3/V4/c3 ;
 wire \V1/V3/V4/overflow ;
 wire \V1/V3/V4/A1/c1 ;
 wire \V1/V3/V4/A1/c2 ;
 wire \V1/V3/V4/A1/c3 ;
 wire \V1/V3/V4/A1/M1/c1 ;
 wire \V1/V3/V4/A1/M1/c2 ;
 wire \V1/V3/V4/A1/M1/s1 ;
 wire \V1/V3/V4/A1/M2/c1 ;
 wire \V1/V3/V4/A1/M2/c2 ;
 wire \V1/V3/V4/A1/M2/s1 ;
 wire \V1/V3/V4/A1/M3/c1 ;
 wire \V1/V3/V4/A1/M3/c2 ;
 wire \V1/V3/V4/A1/M3/s1 ;
 wire \V1/V3/V4/A1/M4/c1 ;
 wire \V1/V3/V4/A1/M4/c2 ;
 wire \V1/V3/V4/A1/M4/s1 ;
 wire \V1/V3/V4/A2/c1 ;
 wire \V1/V3/V4/A2/c2 ;
 wire \V1/V3/V4/A2/c3 ;
 wire \V1/V3/V4/A2/M1/c1 ;
 wire \V1/V3/V4/A2/M1/c2 ;
 wire \V1/V3/V4/A2/M1/s1 ;
 wire \V1/V3/V4/A2/M2/c1 ;
 wire \V1/V3/V4/A2/M2/c2 ;
 wire \V1/V3/V4/A2/M2/s1 ;
 wire \V1/V3/V4/A2/M3/c1 ;
 wire \V1/V3/V4/A2/M3/c2 ;
 wire \V1/V3/V4/A2/M3/s1 ;
 wire \V1/V3/V4/A2/M4/c1 ;
 wire \V1/V3/V4/A2/M4/c2 ;
 wire \V1/V3/V4/A2/M4/s1 ;
 wire \V1/V3/V4/A3/c1 ;
 wire \V1/V3/V4/A3/c2 ;
 wire \V1/V3/V4/A3/c3 ;
 wire \V1/V3/V4/A3/M1/c1 ;
 wire \V1/V3/V4/A3/M1/c2 ;
 wire \V1/V3/V4/A3/M1/s1 ;
 wire \V1/V3/V4/A3/M2/c1 ;
 wire \V1/V3/V4/A3/M2/c2 ;
 wire \V1/V3/V4/A3/M2/s1 ;
 wire \V1/V3/V4/A3/M3/c1 ;
 wire \V1/V3/V4/A3/M3/c2 ;
 wire \V1/V3/V4/A3/M3/s1 ;
 wire \V1/V3/V4/A3/M4/c1 ;
 wire \V1/V3/V4/A3/M4/c2 ;
 wire \V1/V3/V4/A3/M4/s1 ;
 wire \V1/V3/V4/V1/w1 ;
 wire \V1/V3/V4/V1/w2 ;
 wire \V1/V3/V4/V1/w3 ;
 wire \V1/V3/V4/V1/w4 ;
 wire \V1/V3/V4/V2/w1 ;
 wire \V1/V3/V4/V2/w2 ;
 wire \V1/V3/V4/V2/w3 ;
 wire \V1/V3/V4/V2/w4 ;
 wire \V1/V3/V4/V3/w1 ;
 wire \V1/V3/V4/V3/w2 ;
 wire \V1/V3/V4/V3/w3 ;
 wire \V1/V3/V4/V3/w4 ;
 wire \V1/V3/V4/V4/w1 ;
 wire \V1/V3/V4/V4/w2 ;
 wire \V1/V3/V4/V4/w3 ;
 wire \V1/V3/V4/V4/w4 ;
 wire \V1/V4/c1 ;
 wire \V1/V4/c2 ;
 wire \V1/V4/c3 ;
 wire \V1/V4/overflow ;
 wire \V1/V4/A1/c1 ;
 wire \V1/V4/A1/A1/c1 ;
 wire \V1/V4/A1/A1/c2 ;
 wire \V1/V4/A1/A1/c3 ;
 wire \V1/V4/A1/A1/M1/c1 ;
 wire \V1/V4/A1/A1/M1/c2 ;
 wire \V1/V4/A1/A1/M1/s1 ;
 wire \V1/V4/A1/A1/M2/c1 ;
 wire \V1/V4/A1/A1/M2/c2 ;
 wire \V1/V4/A1/A1/M2/s1 ;
 wire \V1/V4/A1/A1/M3/c1 ;
 wire \V1/V4/A1/A1/M3/c2 ;
 wire \V1/V4/A1/A1/M3/s1 ;
 wire \V1/V4/A1/A1/M4/c1 ;
 wire \V1/V4/A1/A1/M4/c2 ;
 wire \V1/V4/A1/A1/M4/s1 ;
 wire \V1/V4/A1/A2/c1 ;
 wire \V1/V4/A1/A2/c2 ;
 wire \V1/V4/A1/A2/c3 ;
 wire \V1/V4/A1/A2/M1/c1 ;
 wire \V1/V4/A1/A2/M1/c2 ;
 wire \V1/V4/A1/A2/M1/s1 ;
 wire \V1/V4/A1/A2/M2/c1 ;
 wire \V1/V4/A1/A2/M2/c2 ;
 wire \V1/V4/A1/A2/M2/s1 ;
 wire \V1/V4/A1/A2/M3/c1 ;
 wire \V1/V4/A1/A2/M3/c2 ;
 wire \V1/V4/A1/A2/M3/s1 ;
 wire \V1/V4/A1/A2/M4/c1 ;
 wire \V1/V4/A1/A2/M4/c2 ;
 wire \V1/V4/A1/A2/M4/s1 ;
 wire \V1/V4/A2/c1 ;
 wire \V1/V4/A2/A1/c1 ;
 wire \V1/V4/A2/A1/c2 ;
 wire \V1/V4/A2/A1/c3 ;
 wire \V1/V4/A2/A1/M1/c1 ;
 wire \V1/V4/A2/A1/M1/c2 ;
 wire \V1/V4/A2/A1/M1/s1 ;
 wire \V1/V4/A2/A1/M2/c1 ;
 wire \V1/V4/A2/A1/M2/c2 ;
 wire \V1/V4/A2/A1/M2/s1 ;
 wire \V1/V4/A2/A1/M3/c1 ;
 wire \V1/V4/A2/A1/M3/c2 ;
 wire \V1/V4/A2/A1/M3/s1 ;
 wire \V1/V4/A2/A1/M4/c1 ;
 wire \V1/V4/A2/A1/M4/c2 ;
 wire \V1/V4/A2/A1/M4/s1 ;
 wire \V1/V4/A2/A2/c1 ;
 wire \V1/V4/A2/A2/c2 ;
 wire \V1/V4/A2/A2/c3 ;
 wire \V1/V4/A2/A2/M1/c1 ;
 wire \V1/V4/A2/A2/M1/c2 ;
 wire \V1/V4/A2/A2/M1/s1 ;
 wire \V1/V4/A2/A2/M2/c1 ;
 wire \V1/V4/A2/A2/M2/c2 ;
 wire \V1/V4/A2/A2/M2/s1 ;
 wire \V1/V4/A2/A2/M3/c1 ;
 wire \V1/V4/A2/A2/M3/c2 ;
 wire \V1/V4/A2/A2/M3/s1 ;
 wire \V1/V4/A2/A2/M4/c1 ;
 wire \V1/V4/A2/A2/M4/c2 ;
 wire \V1/V4/A2/A2/M4/s1 ;
 wire \V1/V4/A3/c1 ;
 wire \V1/V4/A3/A1/c1 ;
 wire \V1/V4/A3/A1/c2 ;
 wire \V1/V4/A3/A1/c3 ;
 wire \V1/V4/A3/A1/M1/c1 ;
 wire \V1/V4/A3/A1/M1/c2 ;
 wire \V1/V4/A3/A1/M1/s1 ;
 wire \V1/V4/A3/A1/M2/c1 ;
 wire \V1/V4/A3/A1/M2/c2 ;
 wire \V1/V4/A3/A1/M2/s1 ;
 wire \V1/V4/A3/A1/M3/c1 ;
 wire \V1/V4/A3/A1/M3/c2 ;
 wire \V1/V4/A3/A1/M3/s1 ;
 wire \V1/V4/A3/A1/M4/c1 ;
 wire \V1/V4/A3/A1/M4/c2 ;
 wire \V1/V4/A3/A1/M4/s1 ;
 wire \V1/V4/A3/A2/c1 ;
 wire \V1/V4/A3/A2/c2 ;
 wire \V1/V4/A3/A2/c3 ;
 wire \V1/V4/A3/A2/M1/c1 ;
 wire \V1/V4/A3/A2/M1/c2 ;
 wire \V1/V4/A3/A2/M1/s1 ;
 wire \V1/V4/A3/A2/M2/c1 ;
 wire \V1/V4/A3/A2/M2/c2 ;
 wire \V1/V4/A3/A2/M2/s1 ;
 wire \V1/V4/A3/A2/M3/c1 ;
 wire \V1/V4/A3/A2/M3/c2 ;
 wire \V1/V4/A3/A2/M3/s1 ;
 wire \V1/V4/A3/A2/M4/c1 ;
 wire \V1/V4/A3/A2/M4/c2 ;
 wire \V1/V4/A3/A2/M4/s1 ;
 wire \V1/V4/V1/c1 ;
 wire \V1/V4/V1/c2 ;
 wire \V1/V4/V1/c3 ;
 wire \V1/V4/V1/overflow ;
 wire \V1/V4/V1/A1/c1 ;
 wire \V1/V4/V1/A1/c2 ;
 wire \V1/V4/V1/A1/c3 ;
 wire \V1/V4/V1/A1/M1/c1 ;
 wire \V1/V4/V1/A1/M1/c2 ;
 wire \V1/V4/V1/A1/M1/s1 ;
 wire \V1/V4/V1/A1/M2/c1 ;
 wire \V1/V4/V1/A1/M2/c2 ;
 wire \V1/V4/V1/A1/M2/s1 ;
 wire \V1/V4/V1/A1/M3/c1 ;
 wire \V1/V4/V1/A1/M3/c2 ;
 wire \V1/V4/V1/A1/M3/s1 ;
 wire \V1/V4/V1/A1/M4/c1 ;
 wire \V1/V4/V1/A1/M4/c2 ;
 wire \V1/V4/V1/A1/M4/s1 ;
 wire \V1/V4/V1/A2/c1 ;
 wire \V1/V4/V1/A2/c2 ;
 wire \V1/V4/V1/A2/c3 ;
 wire \V1/V4/V1/A2/M1/c1 ;
 wire \V1/V4/V1/A2/M1/c2 ;
 wire \V1/V4/V1/A2/M1/s1 ;
 wire \V1/V4/V1/A2/M2/c1 ;
 wire \V1/V4/V1/A2/M2/c2 ;
 wire \V1/V4/V1/A2/M2/s1 ;
 wire \V1/V4/V1/A2/M3/c1 ;
 wire \V1/V4/V1/A2/M3/c2 ;
 wire \V1/V4/V1/A2/M3/s1 ;
 wire \V1/V4/V1/A2/M4/c1 ;
 wire \V1/V4/V1/A2/M4/c2 ;
 wire \V1/V4/V1/A2/M4/s1 ;
 wire \V1/V4/V1/A3/c1 ;
 wire \V1/V4/V1/A3/c2 ;
 wire \V1/V4/V1/A3/c3 ;
 wire \V1/V4/V1/A3/M1/c1 ;
 wire \V1/V4/V1/A3/M1/c2 ;
 wire \V1/V4/V1/A3/M1/s1 ;
 wire \V1/V4/V1/A3/M2/c1 ;
 wire \V1/V4/V1/A3/M2/c2 ;
 wire \V1/V4/V1/A3/M2/s1 ;
 wire \V1/V4/V1/A3/M3/c1 ;
 wire \V1/V4/V1/A3/M3/c2 ;
 wire \V1/V4/V1/A3/M3/s1 ;
 wire \V1/V4/V1/A3/M4/c1 ;
 wire \V1/V4/V1/A3/M4/c2 ;
 wire \V1/V4/V1/A3/M4/s1 ;
 wire \V1/V4/V1/V1/w1 ;
 wire \V1/V4/V1/V1/w2 ;
 wire \V1/V4/V1/V1/w3 ;
 wire \V1/V4/V1/V1/w4 ;
 wire \V1/V4/V1/V2/w1 ;
 wire \V1/V4/V1/V2/w2 ;
 wire \V1/V4/V1/V2/w3 ;
 wire \V1/V4/V1/V2/w4 ;
 wire \V1/V4/V1/V3/w1 ;
 wire \V1/V4/V1/V3/w2 ;
 wire \V1/V4/V1/V3/w3 ;
 wire \V1/V4/V1/V3/w4 ;
 wire \V1/V4/V1/V4/w1 ;
 wire \V1/V4/V1/V4/w2 ;
 wire \V1/V4/V1/V4/w3 ;
 wire \V1/V4/V1/V4/w4 ;
 wire \V1/V4/V2/c1 ;
 wire \V1/V4/V2/c2 ;
 wire \V1/V4/V2/c3 ;
 wire \V1/V4/V2/overflow ;
 wire \V1/V4/V2/A1/c1 ;
 wire \V1/V4/V2/A1/c2 ;
 wire \V1/V4/V2/A1/c3 ;
 wire \V1/V4/V2/A1/M1/c1 ;
 wire \V1/V4/V2/A1/M1/c2 ;
 wire \V1/V4/V2/A1/M1/s1 ;
 wire \V1/V4/V2/A1/M2/c1 ;
 wire \V1/V4/V2/A1/M2/c2 ;
 wire \V1/V4/V2/A1/M2/s1 ;
 wire \V1/V4/V2/A1/M3/c1 ;
 wire \V1/V4/V2/A1/M3/c2 ;
 wire \V1/V4/V2/A1/M3/s1 ;
 wire \V1/V4/V2/A1/M4/c1 ;
 wire \V1/V4/V2/A1/M4/c2 ;
 wire \V1/V4/V2/A1/M4/s1 ;
 wire \V1/V4/V2/A2/c1 ;
 wire \V1/V4/V2/A2/c2 ;
 wire \V1/V4/V2/A2/c3 ;
 wire \V1/V4/V2/A2/M1/c1 ;
 wire \V1/V4/V2/A2/M1/c2 ;
 wire \V1/V4/V2/A2/M1/s1 ;
 wire \V1/V4/V2/A2/M2/c1 ;
 wire \V1/V4/V2/A2/M2/c2 ;
 wire \V1/V4/V2/A2/M2/s1 ;
 wire \V1/V4/V2/A2/M3/c1 ;
 wire \V1/V4/V2/A2/M3/c2 ;
 wire \V1/V4/V2/A2/M3/s1 ;
 wire \V1/V4/V2/A2/M4/c1 ;
 wire \V1/V4/V2/A2/M4/c2 ;
 wire \V1/V4/V2/A2/M4/s1 ;
 wire \V1/V4/V2/A3/c1 ;
 wire \V1/V4/V2/A3/c2 ;
 wire \V1/V4/V2/A3/c3 ;
 wire \V1/V4/V2/A3/M1/c1 ;
 wire \V1/V4/V2/A3/M1/c2 ;
 wire \V1/V4/V2/A3/M1/s1 ;
 wire \V1/V4/V2/A3/M2/c1 ;
 wire \V1/V4/V2/A3/M2/c2 ;
 wire \V1/V4/V2/A3/M2/s1 ;
 wire \V1/V4/V2/A3/M3/c1 ;
 wire \V1/V4/V2/A3/M3/c2 ;
 wire \V1/V4/V2/A3/M3/s1 ;
 wire \V1/V4/V2/A3/M4/c1 ;
 wire \V1/V4/V2/A3/M4/c2 ;
 wire \V1/V4/V2/A3/M4/s1 ;
 wire \V1/V4/V2/V1/w1 ;
 wire \V1/V4/V2/V1/w2 ;
 wire \V1/V4/V2/V1/w3 ;
 wire \V1/V4/V2/V1/w4 ;
 wire \V1/V4/V2/V2/w1 ;
 wire \V1/V4/V2/V2/w2 ;
 wire \V1/V4/V2/V2/w3 ;
 wire \V1/V4/V2/V2/w4 ;
 wire \V1/V4/V2/V3/w1 ;
 wire \V1/V4/V2/V3/w2 ;
 wire \V1/V4/V2/V3/w3 ;
 wire \V1/V4/V2/V3/w4 ;
 wire \V1/V4/V2/V4/w1 ;
 wire \V1/V4/V2/V4/w2 ;
 wire \V1/V4/V2/V4/w3 ;
 wire \V1/V4/V2/V4/w4 ;
 wire \V1/V4/V3/c1 ;
 wire \V1/V4/V3/c2 ;
 wire \V1/V4/V3/c3 ;
 wire \V1/V4/V3/overflow ;
 wire \V1/V4/V3/A1/c1 ;
 wire \V1/V4/V3/A1/c2 ;
 wire \V1/V4/V3/A1/c3 ;
 wire \V1/V4/V3/A1/M1/c1 ;
 wire \V1/V4/V3/A1/M1/c2 ;
 wire \V1/V4/V3/A1/M1/s1 ;
 wire \V1/V4/V3/A1/M2/c1 ;
 wire \V1/V4/V3/A1/M2/c2 ;
 wire \V1/V4/V3/A1/M2/s1 ;
 wire \V1/V4/V3/A1/M3/c1 ;
 wire \V1/V4/V3/A1/M3/c2 ;
 wire \V1/V4/V3/A1/M3/s1 ;
 wire \V1/V4/V3/A1/M4/c1 ;
 wire \V1/V4/V3/A1/M4/c2 ;
 wire \V1/V4/V3/A1/M4/s1 ;
 wire \V1/V4/V3/A2/c1 ;
 wire \V1/V4/V3/A2/c2 ;
 wire \V1/V4/V3/A2/c3 ;
 wire \V1/V4/V3/A2/M1/c1 ;
 wire \V1/V4/V3/A2/M1/c2 ;
 wire \V1/V4/V3/A2/M1/s1 ;
 wire \V1/V4/V3/A2/M2/c1 ;
 wire \V1/V4/V3/A2/M2/c2 ;
 wire \V1/V4/V3/A2/M2/s1 ;
 wire \V1/V4/V3/A2/M3/c1 ;
 wire \V1/V4/V3/A2/M3/c2 ;
 wire \V1/V4/V3/A2/M3/s1 ;
 wire \V1/V4/V3/A2/M4/c1 ;
 wire \V1/V4/V3/A2/M4/c2 ;
 wire \V1/V4/V3/A2/M4/s1 ;
 wire \V1/V4/V3/A3/c1 ;
 wire \V1/V4/V3/A3/c2 ;
 wire \V1/V4/V3/A3/c3 ;
 wire \V1/V4/V3/A3/M1/c1 ;
 wire \V1/V4/V3/A3/M1/c2 ;
 wire \V1/V4/V3/A3/M1/s1 ;
 wire \V1/V4/V3/A3/M2/c1 ;
 wire \V1/V4/V3/A3/M2/c2 ;
 wire \V1/V4/V3/A3/M2/s1 ;
 wire \V1/V4/V3/A3/M3/c1 ;
 wire \V1/V4/V3/A3/M3/c2 ;
 wire \V1/V4/V3/A3/M3/s1 ;
 wire \V1/V4/V3/A3/M4/c1 ;
 wire \V1/V4/V3/A3/M4/c2 ;
 wire \V1/V4/V3/A3/M4/s1 ;
 wire \V1/V4/V3/V1/w1 ;
 wire \V1/V4/V3/V1/w2 ;
 wire \V1/V4/V3/V1/w3 ;
 wire \V1/V4/V3/V1/w4 ;
 wire \V1/V4/V3/V2/w1 ;
 wire \V1/V4/V3/V2/w2 ;
 wire \V1/V4/V3/V2/w3 ;
 wire \V1/V4/V3/V2/w4 ;
 wire \V1/V4/V3/V3/w1 ;
 wire \V1/V4/V3/V3/w2 ;
 wire \V1/V4/V3/V3/w3 ;
 wire \V1/V4/V3/V3/w4 ;
 wire \V1/V4/V3/V4/w1 ;
 wire \V1/V4/V3/V4/w2 ;
 wire \V1/V4/V3/V4/w3 ;
 wire \V1/V4/V3/V4/w4 ;
 wire \V1/V4/V4/c1 ;
 wire \V1/V4/V4/c2 ;
 wire \V1/V4/V4/c3 ;
 wire \V1/V4/V4/overflow ;
 wire \V1/V4/V4/A1/c1 ;
 wire \V1/V4/V4/A1/c2 ;
 wire \V1/V4/V4/A1/c3 ;
 wire \V1/V4/V4/A1/M1/c1 ;
 wire \V1/V4/V4/A1/M1/c2 ;
 wire \V1/V4/V4/A1/M1/s1 ;
 wire \V1/V4/V4/A1/M2/c1 ;
 wire \V1/V4/V4/A1/M2/c2 ;
 wire \V1/V4/V4/A1/M2/s1 ;
 wire \V1/V4/V4/A1/M3/c1 ;
 wire \V1/V4/V4/A1/M3/c2 ;
 wire \V1/V4/V4/A1/M3/s1 ;
 wire \V1/V4/V4/A1/M4/c1 ;
 wire \V1/V4/V4/A1/M4/c2 ;
 wire \V1/V4/V4/A1/M4/s1 ;
 wire \V1/V4/V4/A2/c1 ;
 wire \V1/V4/V4/A2/c2 ;
 wire \V1/V4/V4/A2/c3 ;
 wire \V1/V4/V4/A2/M1/c1 ;
 wire \V1/V4/V4/A2/M1/c2 ;
 wire \V1/V4/V4/A2/M1/s1 ;
 wire \V1/V4/V4/A2/M2/c1 ;
 wire \V1/V4/V4/A2/M2/c2 ;
 wire \V1/V4/V4/A2/M2/s1 ;
 wire \V1/V4/V4/A2/M3/c1 ;
 wire \V1/V4/V4/A2/M3/c2 ;
 wire \V1/V4/V4/A2/M3/s1 ;
 wire \V1/V4/V4/A2/M4/c1 ;
 wire \V1/V4/V4/A2/M4/c2 ;
 wire \V1/V4/V4/A2/M4/s1 ;
 wire \V1/V4/V4/A3/c1 ;
 wire \V1/V4/V4/A3/c2 ;
 wire \V1/V4/V4/A3/c3 ;
 wire \V1/V4/V4/A3/M1/c1 ;
 wire \V1/V4/V4/A3/M1/c2 ;
 wire \V1/V4/V4/A3/M1/s1 ;
 wire \V1/V4/V4/A3/M2/c1 ;
 wire \V1/V4/V4/A3/M2/c2 ;
 wire \V1/V4/V4/A3/M2/s1 ;
 wire \V1/V4/V4/A3/M3/c1 ;
 wire \V1/V4/V4/A3/M3/c2 ;
 wire \V1/V4/V4/A3/M3/s1 ;
 wire \V1/V4/V4/A3/M4/c1 ;
 wire \V1/V4/V4/A3/M4/c2 ;
 wire \V1/V4/V4/A3/M4/s1 ;
 wire \V1/V4/V4/V1/w1 ;
 wire \V1/V4/V4/V1/w2 ;
 wire \V1/V4/V4/V1/w3 ;
 wire \V1/V4/V4/V1/w4 ;
 wire \V1/V4/V4/V2/w1 ;
 wire \V1/V4/V4/V2/w2 ;
 wire \V1/V4/V4/V2/w3 ;
 wire \V1/V4/V4/V2/w4 ;
 wire \V1/V4/V4/V3/w1 ;
 wire \V1/V4/V4/V3/w2 ;
 wire \V1/V4/V4/V3/w3 ;
 wire \V1/V4/V4/V3/w4 ;
 wire \V1/V4/V4/V4/w1 ;
 wire \V1/V4/V4/V4/w2 ;
 wire \V1/V4/V4/V4/w3 ;
 wire \V1/V4/V4/V4/w4 ;
 wire \V2/c1 ;
 wire \V2/c2 ;
 wire \V2/c3 ;
 wire \V2/overflow ;
 wire \V2/A1/c1 ;
 wire \V2/A1/A1/c1 ;
 wire \V2/A1/A1/A1/c1 ;
 wire \V2/A1/A1/A1/c2 ;
 wire \V2/A1/A1/A1/c3 ;
 wire \V2/A1/A1/A1/M1/c1 ;
 wire \V2/A1/A1/A1/M1/c2 ;
 wire \V2/A1/A1/A1/M1/s1 ;
 wire \V2/A1/A1/A1/M2/c1 ;
 wire \V2/A1/A1/A1/M2/c2 ;
 wire \V2/A1/A1/A1/M2/s1 ;
 wire \V2/A1/A1/A1/M3/c1 ;
 wire \V2/A1/A1/A1/M3/c2 ;
 wire \V2/A1/A1/A1/M3/s1 ;
 wire \V2/A1/A1/A1/M4/c1 ;
 wire \V2/A1/A1/A1/M4/c2 ;
 wire \V2/A1/A1/A1/M4/s1 ;
 wire \V2/A1/A1/A2/c1 ;
 wire \V2/A1/A1/A2/c2 ;
 wire \V2/A1/A1/A2/c3 ;
 wire \V2/A1/A1/A2/M1/c1 ;
 wire \V2/A1/A1/A2/M1/c2 ;
 wire \V2/A1/A1/A2/M1/s1 ;
 wire \V2/A1/A1/A2/M2/c1 ;
 wire \V2/A1/A1/A2/M2/c2 ;
 wire \V2/A1/A1/A2/M2/s1 ;
 wire \V2/A1/A1/A2/M3/c1 ;
 wire \V2/A1/A1/A2/M3/c2 ;
 wire \V2/A1/A1/A2/M3/s1 ;
 wire \V2/A1/A1/A2/M4/c1 ;
 wire \V2/A1/A1/A2/M4/c2 ;
 wire \V2/A1/A1/A2/M4/s1 ;
 wire \V2/A1/A2/c1 ;
 wire \V2/A1/A2/A1/c1 ;
 wire \V2/A1/A2/A1/c2 ;
 wire \V2/A1/A2/A1/c3 ;
 wire \V2/A1/A2/A1/M1/c1 ;
 wire \V2/A1/A2/A1/M1/c2 ;
 wire \V2/A1/A2/A1/M1/s1 ;
 wire \V2/A1/A2/A1/M2/c1 ;
 wire \V2/A1/A2/A1/M2/c2 ;
 wire \V2/A1/A2/A1/M2/s1 ;
 wire \V2/A1/A2/A1/M3/c1 ;
 wire \V2/A1/A2/A1/M3/c2 ;
 wire \V2/A1/A2/A1/M3/s1 ;
 wire \V2/A1/A2/A1/M4/c1 ;
 wire \V2/A1/A2/A1/M4/c2 ;
 wire \V2/A1/A2/A1/M4/s1 ;
 wire \V2/A1/A2/A2/c1 ;
 wire \V2/A1/A2/A2/c2 ;
 wire \V2/A1/A2/A2/c3 ;
 wire \V2/A1/A2/A2/M1/c1 ;
 wire \V2/A1/A2/A2/M1/c2 ;
 wire \V2/A1/A2/A2/M1/s1 ;
 wire \V2/A1/A2/A2/M2/c1 ;
 wire \V2/A1/A2/A2/M2/c2 ;
 wire \V2/A1/A2/A2/M2/s1 ;
 wire \V2/A1/A2/A2/M3/c1 ;
 wire \V2/A1/A2/A2/M3/c2 ;
 wire \V2/A1/A2/A2/M3/s1 ;
 wire \V2/A1/A2/A2/M4/c1 ;
 wire \V2/A1/A2/A2/M4/c2 ;
 wire \V2/A1/A2/A2/M4/s1 ;
 wire \V2/A2/c1 ;
 wire \V2/A2/A1/c1 ;
 wire \V2/A2/A1/A1/c1 ;
 wire \V2/A2/A1/A1/c2 ;
 wire \V2/A2/A1/A1/c3 ;
 wire \V2/A2/A1/A1/M1/c1 ;
 wire \V2/A2/A1/A1/M1/c2 ;
 wire \V2/A2/A1/A1/M1/s1 ;
 wire \V2/A2/A1/A1/M2/c1 ;
 wire \V2/A2/A1/A1/M2/c2 ;
 wire \V2/A2/A1/A1/M2/s1 ;
 wire \V2/A2/A1/A1/M3/c1 ;
 wire \V2/A2/A1/A1/M3/c2 ;
 wire \V2/A2/A1/A1/M3/s1 ;
 wire \V2/A2/A1/A1/M4/c1 ;
 wire \V2/A2/A1/A1/M4/c2 ;
 wire \V2/A2/A1/A1/M4/s1 ;
 wire \V2/A2/A1/A2/c1 ;
 wire \V2/A2/A1/A2/c2 ;
 wire \V2/A2/A1/A2/c3 ;
 wire \V2/A2/A1/A2/M1/c1 ;
 wire \V2/A2/A1/A2/M1/c2 ;
 wire \V2/A2/A1/A2/M1/s1 ;
 wire \V2/A2/A1/A2/M2/c1 ;
 wire \V2/A2/A1/A2/M2/c2 ;
 wire \V2/A2/A1/A2/M2/s1 ;
 wire \V2/A2/A1/A2/M3/c1 ;
 wire \V2/A2/A1/A2/M3/c2 ;
 wire \V2/A2/A1/A2/M3/s1 ;
 wire \V2/A2/A1/A2/M4/c1 ;
 wire \V2/A2/A1/A2/M4/c2 ;
 wire \V2/A2/A1/A2/M4/s1 ;
 wire \V2/A2/A2/c1 ;
 wire \V2/A2/A2/A1/c1 ;
 wire \V2/A2/A2/A1/c2 ;
 wire \V2/A2/A2/A1/c3 ;
 wire \V2/A2/A2/A1/M1/c1 ;
 wire \V2/A2/A2/A1/M1/c2 ;
 wire \V2/A2/A2/A1/M1/s1 ;
 wire \V2/A2/A2/A1/M2/c1 ;
 wire \V2/A2/A2/A1/M2/c2 ;
 wire \V2/A2/A2/A1/M2/s1 ;
 wire \V2/A2/A2/A1/M3/c1 ;
 wire \V2/A2/A2/A1/M3/c2 ;
 wire \V2/A2/A2/A1/M3/s1 ;
 wire \V2/A2/A2/A1/M4/c1 ;
 wire \V2/A2/A2/A1/M4/c2 ;
 wire \V2/A2/A2/A1/M4/s1 ;
 wire \V2/A2/A2/A2/c1 ;
 wire \V2/A2/A2/A2/c2 ;
 wire \V2/A2/A2/A2/c3 ;
 wire \V2/A2/A2/A2/M1/c1 ;
 wire \V2/A2/A2/A2/M1/c2 ;
 wire \V2/A2/A2/A2/M1/s1 ;
 wire \V2/A2/A2/A2/M2/c1 ;
 wire \V2/A2/A2/A2/M2/c2 ;
 wire \V2/A2/A2/A2/M2/s1 ;
 wire \V2/A2/A2/A2/M3/c1 ;
 wire \V2/A2/A2/A2/M3/c2 ;
 wire \V2/A2/A2/A2/M3/s1 ;
 wire \V2/A2/A2/A2/M4/c1 ;
 wire \V2/A2/A2/A2/M4/c2 ;
 wire \V2/A2/A2/A2/M4/s1 ;
 wire \V2/A3/c1 ;
 wire \V2/A3/A1/c1 ;
 wire \V2/A3/A1/A1/c1 ;
 wire \V2/A3/A1/A1/c2 ;
 wire \V2/A3/A1/A1/c3 ;
 wire \V2/A3/A1/A1/M1/c1 ;
 wire \V2/A3/A1/A1/M1/c2 ;
 wire \V2/A3/A1/A1/M1/s1 ;
 wire \V2/A3/A1/A1/M2/c1 ;
 wire \V2/A3/A1/A1/M2/c2 ;
 wire \V2/A3/A1/A1/M2/s1 ;
 wire \V2/A3/A1/A1/M3/c1 ;
 wire \V2/A3/A1/A1/M3/c2 ;
 wire \V2/A3/A1/A1/M3/s1 ;
 wire \V2/A3/A1/A1/M4/c1 ;
 wire \V2/A3/A1/A1/M4/c2 ;
 wire \V2/A3/A1/A1/M4/s1 ;
 wire \V2/A3/A1/A2/c1 ;
 wire \V2/A3/A1/A2/c2 ;
 wire \V2/A3/A1/A2/c3 ;
 wire \V2/A3/A1/A2/M1/c1 ;
 wire \V2/A3/A1/A2/M1/c2 ;
 wire \V2/A3/A1/A2/M1/s1 ;
 wire \V2/A3/A1/A2/M2/c1 ;
 wire \V2/A3/A1/A2/M2/c2 ;
 wire \V2/A3/A1/A2/M2/s1 ;
 wire \V2/A3/A1/A2/M3/c1 ;
 wire \V2/A3/A1/A2/M3/c2 ;
 wire \V2/A3/A1/A2/M3/s1 ;
 wire \V2/A3/A1/A2/M4/c1 ;
 wire \V2/A3/A1/A2/M4/c2 ;
 wire \V2/A3/A1/A2/M4/s1 ;
 wire \V2/A3/A2/c1 ;
 wire \V2/A3/A2/A1/c1 ;
 wire \V2/A3/A2/A1/c2 ;
 wire \V2/A3/A2/A1/c3 ;
 wire \V2/A3/A2/A1/M1/c1 ;
 wire \V2/A3/A2/A1/M1/c2 ;
 wire \V2/A3/A2/A1/M1/s1 ;
 wire \V2/A3/A2/A1/M2/c1 ;
 wire \V2/A3/A2/A1/M2/c2 ;
 wire \V2/A3/A2/A1/M2/s1 ;
 wire \V2/A3/A2/A1/M3/c1 ;
 wire \V2/A3/A2/A1/M3/c2 ;
 wire \V2/A3/A2/A1/M3/s1 ;
 wire \V2/A3/A2/A1/M4/c1 ;
 wire \V2/A3/A2/A1/M4/c2 ;
 wire \V2/A3/A2/A1/M4/s1 ;
 wire \V2/A3/A2/A2/c1 ;
 wire \V2/A3/A2/A2/c2 ;
 wire \V2/A3/A2/A2/c3 ;
 wire \V2/A3/A2/A2/M1/c1 ;
 wire \V2/A3/A2/A2/M1/c2 ;
 wire \V2/A3/A2/A2/M1/s1 ;
 wire \V2/A3/A2/A2/M2/c1 ;
 wire \V2/A3/A2/A2/M2/c2 ;
 wire \V2/A3/A2/A2/M2/s1 ;
 wire \V2/A3/A2/A2/M3/c1 ;
 wire \V2/A3/A2/A2/M3/c2 ;
 wire \V2/A3/A2/A2/M3/s1 ;
 wire \V2/A3/A2/A2/M4/c1 ;
 wire \V2/A3/A2/A2/M4/c2 ;
 wire \V2/A3/A2/A2/M4/s1 ;
 wire \V2/V1/c1 ;
 wire \V2/V1/c2 ;
 wire \V2/V1/c3 ;
 wire \V2/V1/overflow ;
 wire \V2/V1/A1/c1 ;
 wire \V2/V1/A1/A1/c1 ;
 wire \V2/V1/A1/A1/c2 ;
 wire \V2/V1/A1/A1/c3 ;
 wire \V2/V1/A1/A1/M1/c1 ;
 wire \V2/V1/A1/A1/M1/c2 ;
 wire \V2/V1/A1/A1/M1/s1 ;
 wire \V2/V1/A1/A1/M2/c1 ;
 wire \V2/V1/A1/A1/M2/c2 ;
 wire \V2/V1/A1/A1/M2/s1 ;
 wire \V2/V1/A1/A1/M3/c1 ;
 wire \V2/V1/A1/A1/M3/c2 ;
 wire \V2/V1/A1/A1/M3/s1 ;
 wire \V2/V1/A1/A1/M4/c1 ;
 wire \V2/V1/A1/A1/M4/c2 ;
 wire \V2/V1/A1/A1/M4/s1 ;
 wire \V2/V1/A1/A2/c1 ;
 wire \V2/V1/A1/A2/c2 ;
 wire \V2/V1/A1/A2/c3 ;
 wire \V2/V1/A1/A2/M1/c1 ;
 wire \V2/V1/A1/A2/M1/c2 ;
 wire \V2/V1/A1/A2/M1/s1 ;
 wire \V2/V1/A1/A2/M2/c1 ;
 wire \V2/V1/A1/A2/M2/c2 ;
 wire \V2/V1/A1/A2/M2/s1 ;
 wire \V2/V1/A1/A2/M3/c1 ;
 wire \V2/V1/A1/A2/M3/c2 ;
 wire \V2/V1/A1/A2/M3/s1 ;
 wire \V2/V1/A1/A2/M4/c1 ;
 wire \V2/V1/A1/A2/M4/c2 ;
 wire \V2/V1/A1/A2/M4/s1 ;
 wire \V2/V1/A2/c1 ;
 wire \V2/V1/A2/A1/c1 ;
 wire \V2/V1/A2/A1/c2 ;
 wire \V2/V1/A2/A1/c3 ;
 wire \V2/V1/A2/A1/M1/c1 ;
 wire \V2/V1/A2/A1/M1/c2 ;
 wire \V2/V1/A2/A1/M1/s1 ;
 wire \V2/V1/A2/A1/M2/c1 ;
 wire \V2/V1/A2/A1/M2/c2 ;
 wire \V2/V1/A2/A1/M2/s1 ;
 wire \V2/V1/A2/A1/M3/c1 ;
 wire \V2/V1/A2/A1/M3/c2 ;
 wire \V2/V1/A2/A1/M3/s1 ;
 wire \V2/V1/A2/A1/M4/c1 ;
 wire \V2/V1/A2/A1/M4/c2 ;
 wire \V2/V1/A2/A1/M4/s1 ;
 wire \V2/V1/A2/A2/c1 ;
 wire \V2/V1/A2/A2/c2 ;
 wire \V2/V1/A2/A2/c3 ;
 wire \V2/V1/A2/A2/M1/c1 ;
 wire \V2/V1/A2/A2/M1/c2 ;
 wire \V2/V1/A2/A2/M1/s1 ;
 wire \V2/V1/A2/A2/M2/c1 ;
 wire \V2/V1/A2/A2/M2/c2 ;
 wire \V2/V1/A2/A2/M2/s1 ;
 wire \V2/V1/A2/A2/M3/c1 ;
 wire \V2/V1/A2/A2/M3/c2 ;
 wire \V2/V1/A2/A2/M3/s1 ;
 wire \V2/V1/A2/A2/M4/c1 ;
 wire \V2/V1/A2/A2/M4/c2 ;
 wire \V2/V1/A2/A2/M4/s1 ;
 wire \V2/V1/A3/c1 ;
 wire \V2/V1/A3/A1/c1 ;
 wire \V2/V1/A3/A1/c2 ;
 wire \V2/V1/A3/A1/c3 ;
 wire \V2/V1/A3/A1/M1/c1 ;
 wire \V2/V1/A3/A1/M1/c2 ;
 wire \V2/V1/A3/A1/M1/s1 ;
 wire \V2/V1/A3/A1/M2/c1 ;
 wire \V2/V1/A3/A1/M2/c2 ;
 wire \V2/V1/A3/A1/M2/s1 ;
 wire \V2/V1/A3/A1/M3/c1 ;
 wire \V2/V1/A3/A1/M3/c2 ;
 wire \V2/V1/A3/A1/M3/s1 ;
 wire \V2/V1/A3/A1/M4/c1 ;
 wire \V2/V1/A3/A1/M4/c2 ;
 wire \V2/V1/A3/A1/M4/s1 ;
 wire \V2/V1/A3/A2/c1 ;
 wire \V2/V1/A3/A2/c2 ;
 wire \V2/V1/A3/A2/c3 ;
 wire \V2/V1/A3/A2/M1/c1 ;
 wire \V2/V1/A3/A2/M1/c2 ;
 wire \V2/V1/A3/A2/M1/s1 ;
 wire \V2/V1/A3/A2/M2/c1 ;
 wire \V2/V1/A3/A2/M2/c2 ;
 wire \V2/V1/A3/A2/M2/s1 ;
 wire \V2/V1/A3/A2/M3/c1 ;
 wire \V2/V1/A3/A2/M3/c2 ;
 wire \V2/V1/A3/A2/M3/s1 ;
 wire \V2/V1/A3/A2/M4/c1 ;
 wire \V2/V1/A3/A2/M4/c2 ;
 wire \V2/V1/A3/A2/M4/s1 ;
 wire \V2/V1/V1/c1 ;
 wire \V2/V1/V1/c2 ;
 wire \V2/V1/V1/c3 ;
 wire \V2/V1/V1/overflow ;
 wire \V2/V1/V1/A1/c1 ;
 wire \V2/V1/V1/A1/c2 ;
 wire \V2/V1/V1/A1/c3 ;
 wire \V2/V1/V1/A1/M1/c1 ;
 wire \V2/V1/V1/A1/M1/c2 ;
 wire \V2/V1/V1/A1/M1/s1 ;
 wire \V2/V1/V1/A1/M2/c1 ;
 wire \V2/V1/V1/A1/M2/c2 ;
 wire \V2/V1/V1/A1/M2/s1 ;
 wire \V2/V1/V1/A1/M3/c1 ;
 wire \V2/V1/V1/A1/M3/c2 ;
 wire \V2/V1/V1/A1/M3/s1 ;
 wire \V2/V1/V1/A1/M4/c1 ;
 wire \V2/V1/V1/A1/M4/c2 ;
 wire \V2/V1/V1/A1/M4/s1 ;
 wire \V2/V1/V1/A2/c1 ;
 wire \V2/V1/V1/A2/c2 ;
 wire \V2/V1/V1/A2/c3 ;
 wire \V2/V1/V1/A2/M1/c1 ;
 wire \V2/V1/V1/A2/M1/c2 ;
 wire \V2/V1/V1/A2/M1/s1 ;
 wire \V2/V1/V1/A2/M2/c1 ;
 wire \V2/V1/V1/A2/M2/c2 ;
 wire \V2/V1/V1/A2/M2/s1 ;
 wire \V2/V1/V1/A2/M3/c1 ;
 wire \V2/V1/V1/A2/M3/c2 ;
 wire \V2/V1/V1/A2/M3/s1 ;
 wire \V2/V1/V1/A2/M4/c1 ;
 wire \V2/V1/V1/A2/M4/c2 ;
 wire \V2/V1/V1/A2/M4/s1 ;
 wire \V2/V1/V1/A3/c1 ;
 wire \V2/V1/V1/A3/c2 ;
 wire \V2/V1/V1/A3/c3 ;
 wire \V2/V1/V1/A3/M1/c1 ;
 wire \V2/V1/V1/A3/M1/c2 ;
 wire \V2/V1/V1/A3/M1/s1 ;
 wire \V2/V1/V1/A3/M2/c1 ;
 wire \V2/V1/V1/A3/M2/c2 ;
 wire \V2/V1/V1/A3/M2/s1 ;
 wire \V2/V1/V1/A3/M3/c1 ;
 wire \V2/V1/V1/A3/M3/c2 ;
 wire \V2/V1/V1/A3/M3/s1 ;
 wire \V2/V1/V1/A3/M4/c1 ;
 wire \V2/V1/V1/A3/M4/c2 ;
 wire \V2/V1/V1/A3/M4/s1 ;
 wire \V2/V1/V1/V1/w1 ;
 wire \V2/V1/V1/V1/w2 ;
 wire \V2/V1/V1/V1/w3 ;
 wire \V2/V1/V1/V1/w4 ;
 wire \V2/V1/V1/V2/w1 ;
 wire \V2/V1/V1/V2/w2 ;
 wire \V2/V1/V1/V2/w3 ;
 wire \V2/V1/V1/V2/w4 ;
 wire \V2/V1/V1/V3/w1 ;
 wire \V2/V1/V1/V3/w2 ;
 wire \V2/V1/V1/V3/w3 ;
 wire \V2/V1/V1/V3/w4 ;
 wire \V2/V1/V1/V4/w1 ;
 wire \V2/V1/V1/V4/w2 ;
 wire \V2/V1/V1/V4/w3 ;
 wire \V2/V1/V1/V4/w4 ;
 wire \V2/V1/V2/c1 ;
 wire \V2/V1/V2/c2 ;
 wire \V2/V1/V2/c3 ;
 wire \V2/V1/V2/overflow ;
 wire \V2/V1/V2/A1/c1 ;
 wire \V2/V1/V2/A1/c2 ;
 wire \V2/V1/V2/A1/c3 ;
 wire \V2/V1/V2/A1/M1/c1 ;
 wire \V2/V1/V2/A1/M1/c2 ;
 wire \V2/V1/V2/A1/M1/s1 ;
 wire \V2/V1/V2/A1/M2/c1 ;
 wire \V2/V1/V2/A1/M2/c2 ;
 wire \V2/V1/V2/A1/M2/s1 ;
 wire \V2/V1/V2/A1/M3/c1 ;
 wire \V2/V1/V2/A1/M3/c2 ;
 wire \V2/V1/V2/A1/M3/s1 ;
 wire \V2/V1/V2/A1/M4/c1 ;
 wire \V2/V1/V2/A1/M4/c2 ;
 wire \V2/V1/V2/A1/M4/s1 ;
 wire \V2/V1/V2/A2/c1 ;
 wire \V2/V1/V2/A2/c2 ;
 wire \V2/V1/V2/A2/c3 ;
 wire \V2/V1/V2/A2/M1/c1 ;
 wire \V2/V1/V2/A2/M1/c2 ;
 wire \V2/V1/V2/A2/M1/s1 ;
 wire \V2/V1/V2/A2/M2/c1 ;
 wire \V2/V1/V2/A2/M2/c2 ;
 wire \V2/V1/V2/A2/M2/s1 ;
 wire \V2/V1/V2/A2/M3/c1 ;
 wire \V2/V1/V2/A2/M3/c2 ;
 wire \V2/V1/V2/A2/M3/s1 ;
 wire \V2/V1/V2/A2/M4/c1 ;
 wire \V2/V1/V2/A2/M4/c2 ;
 wire \V2/V1/V2/A2/M4/s1 ;
 wire \V2/V1/V2/A3/c1 ;
 wire \V2/V1/V2/A3/c2 ;
 wire \V2/V1/V2/A3/c3 ;
 wire \V2/V1/V2/A3/M1/c1 ;
 wire \V2/V1/V2/A3/M1/c2 ;
 wire \V2/V1/V2/A3/M1/s1 ;
 wire \V2/V1/V2/A3/M2/c1 ;
 wire \V2/V1/V2/A3/M2/c2 ;
 wire \V2/V1/V2/A3/M2/s1 ;
 wire \V2/V1/V2/A3/M3/c1 ;
 wire \V2/V1/V2/A3/M3/c2 ;
 wire \V2/V1/V2/A3/M3/s1 ;
 wire \V2/V1/V2/A3/M4/c1 ;
 wire \V2/V1/V2/A3/M4/c2 ;
 wire \V2/V1/V2/A3/M4/s1 ;
 wire \V2/V1/V2/V1/w1 ;
 wire \V2/V1/V2/V1/w2 ;
 wire \V2/V1/V2/V1/w3 ;
 wire \V2/V1/V2/V1/w4 ;
 wire \V2/V1/V2/V2/w1 ;
 wire \V2/V1/V2/V2/w2 ;
 wire \V2/V1/V2/V2/w3 ;
 wire \V2/V1/V2/V2/w4 ;
 wire \V2/V1/V2/V3/w1 ;
 wire \V2/V1/V2/V3/w2 ;
 wire \V2/V1/V2/V3/w3 ;
 wire \V2/V1/V2/V3/w4 ;
 wire \V2/V1/V2/V4/w1 ;
 wire \V2/V1/V2/V4/w2 ;
 wire \V2/V1/V2/V4/w3 ;
 wire \V2/V1/V2/V4/w4 ;
 wire \V2/V1/V3/c1 ;
 wire \V2/V1/V3/c2 ;
 wire \V2/V1/V3/c3 ;
 wire \V2/V1/V3/overflow ;
 wire \V2/V1/V3/A1/c1 ;
 wire \V2/V1/V3/A1/c2 ;
 wire \V2/V1/V3/A1/c3 ;
 wire \V2/V1/V3/A1/M1/c1 ;
 wire \V2/V1/V3/A1/M1/c2 ;
 wire \V2/V1/V3/A1/M1/s1 ;
 wire \V2/V1/V3/A1/M2/c1 ;
 wire \V2/V1/V3/A1/M2/c2 ;
 wire \V2/V1/V3/A1/M2/s1 ;
 wire \V2/V1/V3/A1/M3/c1 ;
 wire \V2/V1/V3/A1/M3/c2 ;
 wire \V2/V1/V3/A1/M3/s1 ;
 wire \V2/V1/V3/A1/M4/c1 ;
 wire \V2/V1/V3/A1/M4/c2 ;
 wire \V2/V1/V3/A1/M4/s1 ;
 wire \V2/V1/V3/A2/c1 ;
 wire \V2/V1/V3/A2/c2 ;
 wire \V2/V1/V3/A2/c3 ;
 wire \V2/V1/V3/A2/M1/c1 ;
 wire \V2/V1/V3/A2/M1/c2 ;
 wire \V2/V1/V3/A2/M1/s1 ;
 wire \V2/V1/V3/A2/M2/c1 ;
 wire \V2/V1/V3/A2/M2/c2 ;
 wire \V2/V1/V3/A2/M2/s1 ;
 wire \V2/V1/V3/A2/M3/c1 ;
 wire \V2/V1/V3/A2/M3/c2 ;
 wire \V2/V1/V3/A2/M3/s1 ;
 wire \V2/V1/V3/A2/M4/c1 ;
 wire \V2/V1/V3/A2/M4/c2 ;
 wire \V2/V1/V3/A2/M4/s1 ;
 wire \V2/V1/V3/A3/c1 ;
 wire \V2/V1/V3/A3/c2 ;
 wire \V2/V1/V3/A3/c3 ;
 wire \V2/V1/V3/A3/M1/c1 ;
 wire \V2/V1/V3/A3/M1/c2 ;
 wire \V2/V1/V3/A3/M1/s1 ;
 wire \V2/V1/V3/A3/M2/c1 ;
 wire \V2/V1/V3/A3/M2/c2 ;
 wire \V2/V1/V3/A3/M2/s1 ;
 wire \V2/V1/V3/A3/M3/c1 ;
 wire \V2/V1/V3/A3/M3/c2 ;
 wire \V2/V1/V3/A3/M3/s1 ;
 wire \V2/V1/V3/A3/M4/c1 ;
 wire \V2/V1/V3/A3/M4/c2 ;
 wire \V2/V1/V3/A3/M4/s1 ;
 wire \V2/V1/V3/V1/w1 ;
 wire \V2/V1/V3/V1/w2 ;
 wire \V2/V1/V3/V1/w3 ;
 wire \V2/V1/V3/V1/w4 ;
 wire \V2/V1/V3/V2/w1 ;
 wire \V2/V1/V3/V2/w2 ;
 wire \V2/V1/V3/V2/w3 ;
 wire \V2/V1/V3/V2/w4 ;
 wire \V2/V1/V3/V3/w1 ;
 wire \V2/V1/V3/V3/w2 ;
 wire \V2/V1/V3/V3/w3 ;
 wire \V2/V1/V3/V3/w4 ;
 wire \V2/V1/V3/V4/w1 ;
 wire \V2/V1/V3/V4/w2 ;
 wire \V2/V1/V3/V4/w3 ;
 wire \V2/V1/V3/V4/w4 ;
 wire \V2/V1/V4/c1 ;
 wire \V2/V1/V4/c2 ;
 wire \V2/V1/V4/c3 ;
 wire \V2/V1/V4/overflow ;
 wire \V2/V1/V4/A1/c1 ;
 wire \V2/V1/V4/A1/c2 ;
 wire \V2/V1/V4/A1/c3 ;
 wire \V2/V1/V4/A1/M1/c1 ;
 wire \V2/V1/V4/A1/M1/c2 ;
 wire \V2/V1/V4/A1/M1/s1 ;
 wire \V2/V1/V4/A1/M2/c1 ;
 wire \V2/V1/V4/A1/M2/c2 ;
 wire \V2/V1/V4/A1/M2/s1 ;
 wire \V2/V1/V4/A1/M3/c1 ;
 wire \V2/V1/V4/A1/M3/c2 ;
 wire \V2/V1/V4/A1/M3/s1 ;
 wire \V2/V1/V4/A1/M4/c1 ;
 wire \V2/V1/V4/A1/M4/c2 ;
 wire \V2/V1/V4/A1/M4/s1 ;
 wire \V2/V1/V4/A2/c1 ;
 wire \V2/V1/V4/A2/c2 ;
 wire \V2/V1/V4/A2/c3 ;
 wire \V2/V1/V4/A2/M1/c1 ;
 wire \V2/V1/V4/A2/M1/c2 ;
 wire \V2/V1/V4/A2/M1/s1 ;
 wire \V2/V1/V4/A2/M2/c1 ;
 wire \V2/V1/V4/A2/M2/c2 ;
 wire \V2/V1/V4/A2/M2/s1 ;
 wire \V2/V1/V4/A2/M3/c1 ;
 wire \V2/V1/V4/A2/M3/c2 ;
 wire \V2/V1/V4/A2/M3/s1 ;
 wire \V2/V1/V4/A2/M4/c1 ;
 wire \V2/V1/V4/A2/M4/c2 ;
 wire \V2/V1/V4/A2/M4/s1 ;
 wire \V2/V1/V4/A3/c1 ;
 wire \V2/V1/V4/A3/c2 ;
 wire \V2/V1/V4/A3/c3 ;
 wire \V2/V1/V4/A3/M1/c1 ;
 wire \V2/V1/V4/A3/M1/c2 ;
 wire \V2/V1/V4/A3/M1/s1 ;
 wire \V2/V1/V4/A3/M2/c1 ;
 wire \V2/V1/V4/A3/M2/c2 ;
 wire \V2/V1/V4/A3/M2/s1 ;
 wire \V2/V1/V4/A3/M3/c1 ;
 wire \V2/V1/V4/A3/M3/c2 ;
 wire \V2/V1/V4/A3/M3/s1 ;
 wire \V2/V1/V4/A3/M4/c1 ;
 wire \V2/V1/V4/A3/M4/c2 ;
 wire \V2/V1/V4/A3/M4/s1 ;
 wire \V2/V1/V4/V1/w1 ;
 wire \V2/V1/V4/V1/w2 ;
 wire \V2/V1/V4/V1/w3 ;
 wire \V2/V1/V4/V1/w4 ;
 wire \V2/V1/V4/V2/w1 ;
 wire \V2/V1/V4/V2/w2 ;
 wire \V2/V1/V4/V2/w3 ;
 wire \V2/V1/V4/V2/w4 ;
 wire \V2/V1/V4/V3/w1 ;
 wire \V2/V1/V4/V3/w2 ;
 wire \V2/V1/V4/V3/w3 ;
 wire \V2/V1/V4/V3/w4 ;
 wire \V2/V1/V4/V4/w1 ;
 wire \V2/V1/V4/V4/w2 ;
 wire \V2/V1/V4/V4/w3 ;
 wire \V2/V1/V4/V4/w4 ;
 wire \V2/V2/c1 ;
 wire \V2/V2/c2 ;
 wire \V2/V2/c3 ;
 wire \V2/V2/overflow ;
 wire \V2/V2/A1/c1 ;
 wire \V2/V2/A1/A1/c1 ;
 wire \V2/V2/A1/A1/c2 ;
 wire \V2/V2/A1/A1/c3 ;
 wire \V2/V2/A1/A1/M1/c1 ;
 wire \V2/V2/A1/A1/M1/c2 ;
 wire \V2/V2/A1/A1/M1/s1 ;
 wire \V2/V2/A1/A1/M2/c1 ;
 wire \V2/V2/A1/A1/M2/c2 ;
 wire \V2/V2/A1/A1/M2/s1 ;
 wire \V2/V2/A1/A1/M3/c1 ;
 wire \V2/V2/A1/A1/M3/c2 ;
 wire \V2/V2/A1/A1/M3/s1 ;
 wire \V2/V2/A1/A1/M4/c1 ;
 wire \V2/V2/A1/A1/M4/c2 ;
 wire \V2/V2/A1/A1/M4/s1 ;
 wire \V2/V2/A1/A2/c1 ;
 wire \V2/V2/A1/A2/c2 ;
 wire \V2/V2/A1/A2/c3 ;
 wire \V2/V2/A1/A2/M1/c1 ;
 wire \V2/V2/A1/A2/M1/c2 ;
 wire \V2/V2/A1/A2/M1/s1 ;
 wire \V2/V2/A1/A2/M2/c1 ;
 wire \V2/V2/A1/A2/M2/c2 ;
 wire \V2/V2/A1/A2/M2/s1 ;
 wire \V2/V2/A1/A2/M3/c1 ;
 wire \V2/V2/A1/A2/M3/c2 ;
 wire \V2/V2/A1/A2/M3/s1 ;
 wire \V2/V2/A1/A2/M4/c1 ;
 wire \V2/V2/A1/A2/M4/c2 ;
 wire \V2/V2/A1/A2/M4/s1 ;
 wire \V2/V2/A2/c1 ;
 wire \V2/V2/A2/A1/c1 ;
 wire \V2/V2/A2/A1/c2 ;
 wire \V2/V2/A2/A1/c3 ;
 wire \V2/V2/A2/A1/M1/c1 ;
 wire \V2/V2/A2/A1/M1/c2 ;
 wire \V2/V2/A2/A1/M1/s1 ;
 wire \V2/V2/A2/A1/M2/c1 ;
 wire \V2/V2/A2/A1/M2/c2 ;
 wire \V2/V2/A2/A1/M2/s1 ;
 wire \V2/V2/A2/A1/M3/c1 ;
 wire \V2/V2/A2/A1/M3/c2 ;
 wire \V2/V2/A2/A1/M3/s1 ;
 wire \V2/V2/A2/A1/M4/c1 ;
 wire \V2/V2/A2/A1/M4/c2 ;
 wire \V2/V2/A2/A1/M4/s1 ;
 wire \V2/V2/A2/A2/c1 ;
 wire \V2/V2/A2/A2/c2 ;
 wire \V2/V2/A2/A2/c3 ;
 wire \V2/V2/A2/A2/M1/c1 ;
 wire \V2/V2/A2/A2/M1/c2 ;
 wire \V2/V2/A2/A2/M1/s1 ;
 wire \V2/V2/A2/A2/M2/c1 ;
 wire \V2/V2/A2/A2/M2/c2 ;
 wire \V2/V2/A2/A2/M2/s1 ;
 wire \V2/V2/A2/A2/M3/c1 ;
 wire \V2/V2/A2/A2/M3/c2 ;
 wire \V2/V2/A2/A2/M3/s1 ;
 wire \V2/V2/A2/A2/M4/c1 ;
 wire \V2/V2/A2/A2/M4/c2 ;
 wire \V2/V2/A2/A2/M4/s1 ;
 wire \V2/V2/A3/c1 ;
 wire \V2/V2/A3/A1/c1 ;
 wire \V2/V2/A3/A1/c2 ;
 wire \V2/V2/A3/A1/c3 ;
 wire \V2/V2/A3/A1/M1/c1 ;
 wire \V2/V2/A3/A1/M1/c2 ;
 wire \V2/V2/A3/A1/M1/s1 ;
 wire \V2/V2/A3/A1/M2/c1 ;
 wire \V2/V2/A3/A1/M2/c2 ;
 wire \V2/V2/A3/A1/M2/s1 ;
 wire \V2/V2/A3/A1/M3/c1 ;
 wire \V2/V2/A3/A1/M3/c2 ;
 wire \V2/V2/A3/A1/M3/s1 ;
 wire \V2/V2/A3/A1/M4/c1 ;
 wire \V2/V2/A3/A1/M4/c2 ;
 wire \V2/V2/A3/A1/M4/s1 ;
 wire \V2/V2/A3/A2/c1 ;
 wire \V2/V2/A3/A2/c2 ;
 wire \V2/V2/A3/A2/c3 ;
 wire \V2/V2/A3/A2/M1/c1 ;
 wire \V2/V2/A3/A2/M1/c2 ;
 wire \V2/V2/A3/A2/M1/s1 ;
 wire \V2/V2/A3/A2/M2/c1 ;
 wire \V2/V2/A3/A2/M2/c2 ;
 wire \V2/V2/A3/A2/M2/s1 ;
 wire \V2/V2/A3/A2/M3/c1 ;
 wire \V2/V2/A3/A2/M3/c2 ;
 wire \V2/V2/A3/A2/M3/s1 ;
 wire \V2/V2/A3/A2/M4/c1 ;
 wire \V2/V2/A3/A2/M4/c2 ;
 wire \V2/V2/A3/A2/M4/s1 ;
 wire \V2/V2/V1/c1 ;
 wire \V2/V2/V1/c2 ;
 wire \V2/V2/V1/c3 ;
 wire \V2/V2/V1/overflow ;
 wire \V2/V2/V1/A1/c1 ;
 wire \V2/V2/V1/A1/c2 ;
 wire \V2/V2/V1/A1/c3 ;
 wire \V2/V2/V1/A1/M1/c1 ;
 wire \V2/V2/V1/A1/M1/c2 ;
 wire \V2/V2/V1/A1/M1/s1 ;
 wire \V2/V2/V1/A1/M2/c1 ;
 wire \V2/V2/V1/A1/M2/c2 ;
 wire \V2/V2/V1/A1/M2/s1 ;
 wire \V2/V2/V1/A1/M3/c1 ;
 wire \V2/V2/V1/A1/M3/c2 ;
 wire \V2/V2/V1/A1/M3/s1 ;
 wire \V2/V2/V1/A1/M4/c1 ;
 wire \V2/V2/V1/A1/M4/c2 ;
 wire \V2/V2/V1/A1/M4/s1 ;
 wire \V2/V2/V1/A2/c1 ;
 wire \V2/V2/V1/A2/c2 ;
 wire \V2/V2/V1/A2/c3 ;
 wire \V2/V2/V1/A2/M1/c1 ;
 wire \V2/V2/V1/A2/M1/c2 ;
 wire \V2/V2/V1/A2/M1/s1 ;
 wire \V2/V2/V1/A2/M2/c1 ;
 wire \V2/V2/V1/A2/M2/c2 ;
 wire \V2/V2/V1/A2/M2/s1 ;
 wire \V2/V2/V1/A2/M3/c1 ;
 wire \V2/V2/V1/A2/M3/c2 ;
 wire \V2/V2/V1/A2/M3/s1 ;
 wire \V2/V2/V1/A2/M4/c1 ;
 wire \V2/V2/V1/A2/M4/c2 ;
 wire \V2/V2/V1/A2/M4/s1 ;
 wire \V2/V2/V1/A3/c1 ;
 wire \V2/V2/V1/A3/c2 ;
 wire \V2/V2/V1/A3/c3 ;
 wire \V2/V2/V1/A3/M1/c1 ;
 wire \V2/V2/V1/A3/M1/c2 ;
 wire \V2/V2/V1/A3/M1/s1 ;
 wire \V2/V2/V1/A3/M2/c1 ;
 wire \V2/V2/V1/A3/M2/c2 ;
 wire \V2/V2/V1/A3/M2/s1 ;
 wire \V2/V2/V1/A3/M3/c1 ;
 wire \V2/V2/V1/A3/M3/c2 ;
 wire \V2/V2/V1/A3/M3/s1 ;
 wire \V2/V2/V1/A3/M4/c1 ;
 wire \V2/V2/V1/A3/M4/c2 ;
 wire \V2/V2/V1/A3/M4/s1 ;
 wire \V2/V2/V1/V1/w1 ;
 wire \V2/V2/V1/V1/w2 ;
 wire \V2/V2/V1/V1/w3 ;
 wire \V2/V2/V1/V1/w4 ;
 wire \V2/V2/V1/V2/w1 ;
 wire \V2/V2/V1/V2/w2 ;
 wire \V2/V2/V1/V2/w3 ;
 wire \V2/V2/V1/V2/w4 ;
 wire \V2/V2/V1/V3/w1 ;
 wire \V2/V2/V1/V3/w2 ;
 wire \V2/V2/V1/V3/w3 ;
 wire \V2/V2/V1/V3/w4 ;
 wire \V2/V2/V1/V4/w1 ;
 wire \V2/V2/V1/V4/w2 ;
 wire \V2/V2/V1/V4/w3 ;
 wire \V2/V2/V1/V4/w4 ;
 wire \V2/V2/V2/c1 ;
 wire \V2/V2/V2/c2 ;
 wire \V2/V2/V2/c3 ;
 wire \V2/V2/V2/overflow ;
 wire \V2/V2/V2/A1/c1 ;
 wire \V2/V2/V2/A1/c2 ;
 wire \V2/V2/V2/A1/c3 ;
 wire \V2/V2/V2/A1/M1/c1 ;
 wire \V2/V2/V2/A1/M1/c2 ;
 wire \V2/V2/V2/A1/M1/s1 ;
 wire \V2/V2/V2/A1/M2/c1 ;
 wire \V2/V2/V2/A1/M2/c2 ;
 wire \V2/V2/V2/A1/M2/s1 ;
 wire \V2/V2/V2/A1/M3/c1 ;
 wire \V2/V2/V2/A1/M3/c2 ;
 wire \V2/V2/V2/A1/M3/s1 ;
 wire \V2/V2/V2/A1/M4/c1 ;
 wire \V2/V2/V2/A1/M4/c2 ;
 wire \V2/V2/V2/A1/M4/s1 ;
 wire \V2/V2/V2/A2/c1 ;
 wire \V2/V2/V2/A2/c2 ;
 wire \V2/V2/V2/A2/c3 ;
 wire \V2/V2/V2/A2/M1/c1 ;
 wire \V2/V2/V2/A2/M1/c2 ;
 wire \V2/V2/V2/A2/M1/s1 ;
 wire \V2/V2/V2/A2/M2/c1 ;
 wire \V2/V2/V2/A2/M2/c2 ;
 wire \V2/V2/V2/A2/M2/s1 ;
 wire \V2/V2/V2/A2/M3/c1 ;
 wire \V2/V2/V2/A2/M3/c2 ;
 wire \V2/V2/V2/A2/M3/s1 ;
 wire \V2/V2/V2/A2/M4/c1 ;
 wire \V2/V2/V2/A2/M4/c2 ;
 wire \V2/V2/V2/A2/M4/s1 ;
 wire \V2/V2/V2/A3/c1 ;
 wire \V2/V2/V2/A3/c2 ;
 wire \V2/V2/V2/A3/c3 ;
 wire \V2/V2/V2/A3/M1/c1 ;
 wire \V2/V2/V2/A3/M1/c2 ;
 wire \V2/V2/V2/A3/M1/s1 ;
 wire \V2/V2/V2/A3/M2/c1 ;
 wire \V2/V2/V2/A3/M2/c2 ;
 wire \V2/V2/V2/A3/M2/s1 ;
 wire \V2/V2/V2/A3/M3/c1 ;
 wire \V2/V2/V2/A3/M3/c2 ;
 wire \V2/V2/V2/A3/M3/s1 ;
 wire \V2/V2/V2/A3/M4/c1 ;
 wire \V2/V2/V2/A3/M4/c2 ;
 wire \V2/V2/V2/A3/M4/s1 ;
 wire \V2/V2/V2/V1/w1 ;
 wire \V2/V2/V2/V1/w2 ;
 wire \V2/V2/V2/V1/w3 ;
 wire \V2/V2/V2/V1/w4 ;
 wire \V2/V2/V2/V2/w1 ;
 wire \V2/V2/V2/V2/w2 ;
 wire \V2/V2/V2/V2/w3 ;
 wire \V2/V2/V2/V2/w4 ;
 wire \V2/V2/V2/V3/w1 ;
 wire \V2/V2/V2/V3/w2 ;
 wire \V2/V2/V2/V3/w3 ;
 wire \V2/V2/V2/V3/w4 ;
 wire \V2/V2/V2/V4/w1 ;
 wire \V2/V2/V2/V4/w2 ;
 wire \V2/V2/V2/V4/w3 ;
 wire \V2/V2/V2/V4/w4 ;
 wire \V2/V2/V3/c1 ;
 wire \V2/V2/V3/c2 ;
 wire \V2/V2/V3/c3 ;
 wire \V2/V2/V3/overflow ;
 wire \V2/V2/V3/A1/c1 ;
 wire \V2/V2/V3/A1/c2 ;
 wire \V2/V2/V3/A1/c3 ;
 wire \V2/V2/V3/A1/M1/c1 ;
 wire \V2/V2/V3/A1/M1/c2 ;
 wire \V2/V2/V3/A1/M1/s1 ;
 wire \V2/V2/V3/A1/M2/c1 ;
 wire \V2/V2/V3/A1/M2/c2 ;
 wire \V2/V2/V3/A1/M2/s1 ;
 wire \V2/V2/V3/A1/M3/c1 ;
 wire \V2/V2/V3/A1/M3/c2 ;
 wire \V2/V2/V3/A1/M3/s1 ;
 wire \V2/V2/V3/A1/M4/c1 ;
 wire \V2/V2/V3/A1/M4/c2 ;
 wire \V2/V2/V3/A1/M4/s1 ;
 wire \V2/V2/V3/A2/c1 ;
 wire \V2/V2/V3/A2/c2 ;
 wire \V2/V2/V3/A2/c3 ;
 wire \V2/V2/V3/A2/M1/c1 ;
 wire \V2/V2/V3/A2/M1/c2 ;
 wire \V2/V2/V3/A2/M1/s1 ;
 wire \V2/V2/V3/A2/M2/c1 ;
 wire \V2/V2/V3/A2/M2/c2 ;
 wire \V2/V2/V3/A2/M2/s1 ;
 wire \V2/V2/V3/A2/M3/c1 ;
 wire \V2/V2/V3/A2/M3/c2 ;
 wire \V2/V2/V3/A2/M3/s1 ;
 wire \V2/V2/V3/A2/M4/c1 ;
 wire \V2/V2/V3/A2/M4/c2 ;
 wire \V2/V2/V3/A2/M4/s1 ;
 wire \V2/V2/V3/A3/c1 ;
 wire \V2/V2/V3/A3/c2 ;
 wire \V2/V2/V3/A3/c3 ;
 wire \V2/V2/V3/A3/M1/c1 ;
 wire \V2/V2/V3/A3/M1/c2 ;
 wire \V2/V2/V3/A3/M1/s1 ;
 wire \V2/V2/V3/A3/M2/c1 ;
 wire \V2/V2/V3/A3/M2/c2 ;
 wire \V2/V2/V3/A3/M2/s1 ;
 wire \V2/V2/V3/A3/M3/c1 ;
 wire \V2/V2/V3/A3/M3/c2 ;
 wire \V2/V2/V3/A3/M3/s1 ;
 wire \V2/V2/V3/A3/M4/c1 ;
 wire \V2/V2/V3/A3/M4/c2 ;
 wire \V2/V2/V3/A3/M4/s1 ;
 wire \V2/V2/V3/V1/w1 ;
 wire \V2/V2/V3/V1/w2 ;
 wire \V2/V2/V3/V1/w3 ;
 wire \V2/V2/V3/V1/w4 ;
 wire \V2/V2/V3/V2/w1 ;
 wire \V2/V2/V3/V2/w2 ;
 wire \V2/V2/V3/V2/w3 ;
 wire \V2/V2/V3/V2/w4 ;
 wire \V2/V2/V3/V3/w1 ;
 wire \V2/V2/V3/V3/w2 ;
 wire \V2/V2/V3/V3/w3 ;
 wire \V2/V2/V3/V3/w4 ;
 wire \V2/V2/V3/V4/w1 ;
 wire \V2/V2/V3/V4/w2 ;
 wire \V2/V2/V3/V4/w3 ;
 wire \V2/V2/V3/V4/w4 ;
 wire \V2/V2/V4/c1 ;
 wire \V2/V2/V4/c2 ;
 wire \V2/V2/V4/c3 ;
 wire \V2/V2/V4/overflow ;
 wire \V2/V2/V4/A1/c1 ;
 wire \V2/V2/V4/A1/c2 ;
 wire \V2/V2/V4/A1/c3 ;
 wire \V2/V2/V4/A1/M1/c1 ;
 wire \V2/V2/V4/A1/M1/c2 ;
 wire \V2/V2/V4/A1/M1/s1 ;
 wire \V2/V2/V4/A1/M2/c1 ;
 wire \V2/V2/V4/A1/M2/c2 ;
 wire \V2/V2/V4/A1/M2/s1 ;
 wire \V2/V2/V4/A1/M3/c1 ;
 wire \V2/V2/V4/A1/M3/c2 ;
 wire \V2/V2/V4/A1/M3/s1 ;
 wire \V2/V2/V4/A1/M4/c1 ;
 wire \V2/V2/V4/A1/M4/c2 ;
 wire \V2/V2/V4/A1/M4/s1 ;
 wire \V2/V2/V4/A2/c1 ;
 wire \V2/V2/V4/A2/c2 ;
 wire \V2/V2/V4/A2/c3 ;
 wire \V2/V2/V4/A2/M1/c1 ;
 wire \V2/V2/V4/A2/M1/c2 ;
 wire \V2/V2/V4/A2/M1/s1 ;
 wire \V2/V2/V4/A2/M2/c1 ;
 wire \V2/V2/V4/A2/M2/c2 ;
 wire \V2/V2/V4/A2/M2/s1 ;
 wire \V2/V2/V4/A2/M3/c1 ;
 wire \V2/V2/V4/A2/M3/c2 ;
 wire \V2/V2/V4/A2/M3/s1 ;
 wire \V2/V2/V4/A2/M4/c1 ;
 wire \V2/V2/V4/A2/M4/c2 ;
 wire \V2/V2/V4/A2/M4/s1 ;
 wire \V2/V2/V4/A3/c1 ;
 wire \V2/V2/V4/A3/c2 ;
 wire \V2/V2/V4/A3/c3 ;
 wire \V2/V2/V4/A3/M1/c1 ;
 wire \V2/V2/V4/A3/M1/c2 ;
 wire \V2/V2/V4/A3/M1/s1 ;
 wire \V2/V2/V4/A3/M2/c1 ;
 wire \V2/V2/V4/A3/M2/c2 ;
 wire \V2/V2/V4/A3/M2/s1 ;
 wire \V2/V2/V4/A3/M3/c1 ;
 wire \V2/V2/V4/A3/M3/c2 ;
 wire \V2/V2/V4/A3/M3/s1 ;
 wire \V2/V2/V4/A3/M4/c1 ;
 wire \V2/V2/V4/A3/M4/c2 ;
 wire \V2/V2/V4/A3/M4/s1 ;
 wire \V2/V2/V4/V1/w1 ;
 wire \V2/V2/V4/V1/w2 ;
 wire \V2/V2/V4/V1/w3 ;
 wire \V2/V2/V4/V1/w4 ;
 wire \V2/V2/V4/V2/w1 ;
 wire \V2/V2/V4/V2/w2 ;
 wire \V2/V2/V4/V2/w3 ;
 wire \V2/V2/V4/V2/w4 ;
 wire \V2/V2/V4/V3/w1 ;
 wire \V2/V2/V4/V3/w2 ;
 wire \V2/V2/V4/V3/w3 ;
 wire \V2/V2/V4/V3/w4 ;
 wire \V2/V2/V4/V4/w1 ;
 wire \V2/V2/V4/V4/w2 ;
 wire \V2/V2/V4/V4/w3 ;
 wire \V2/V2/V4/V4/w4 ;
 wire \V2/V3/c1 ;
 wire \V2/V3/c2 ;
 wire \V2/V3/c3 ;
 wire \V2/V3/overflow ;
 wire \V2/V3/A1/c1 ;
 wire \V2/V3/A1/A1/c1 ;
 wire \V2/V3/A1/A1/c2 ;
 wire \V2/V3/A1/A1/c3 ;
 wire \V2/V3/A1/A1/M1/c1 ;
 wire \V2/V3/A1/A1/M1/c2 ;
 wire \V2/V3/A1/A1/M1/s1 ;
 wire \V2/V3/A1/A1/M2/c1 ;
 wire \V2/V3/A1/A1/M2/c2 ;
 wire \V2/V3/A1/A1/M2/s1 ;
 wire \V2/V3/A1/A1/M3/c1 ;
 wire \V2/V3/A1/A1/M3/c2 ;
 wire \V2/V3/A1/A1/M3/s1 ;
 wire \V2/V3/A1/A1/M4/c1 ;
 wire \V2/V3/A1/A1/M4/c2 ;
 wire \V2/V3/A1/A1/M4/s1 ;
 wire \V2/V3/A1/A2/c1 ;
 wire \V2/V3/A1/A2/c2 ;
 wire \V2/V3/A1/A2/c3 ;
 wire \V2/V3/A1/A2/M1/c1 ;
 wire \V2/V3/A1/A2/M1/c2 ;
 wire \V2/V3/A1/A2/M1/s1 ;
 wire \V2/V3/A1/A2/M2/c1 ;
 wire \V2/V3/A1/A2/M2/c2 ;
 wire \V2/V3/A1/A2/M2/s1 ;
 wire \V2/V3/A1/A2/M3/c1 ;
 wire \V2/V3/A1/A2/M3/c2 ;
 wire \V2/V3/A1/A2/M3/s1 ;
 wire \V2/V3/A1/A2/M4/c1 ;
 wire \V2/V3/A1/A2/M4/c2 ;
 wire \V2/V3/A1/A2/M4/s1 ;
 wire \V2/V3/A2/c1 ;
 wire \V2/V3/A2/A1/c1 ;
 wire \V2/V3/A2/A1/c2 ;
 wire \V2/V3/A2/A1/c3 ;
 wire \V2/V3/A2/A1/M1/c1 ;
 wire \V2/V3/A2/A1/M1/c2 ;
 wire \V2/V3/A2/A1/M1/s1 ;
 wire \V2/V3/A2/A1/M2/c1 ;
 wire \V2/V3/A2/A1/M2/c2 ;
 wire \V2/V3/A2/A1/M2/s1 ;
 wire \V2/V3/A2/A1/M3/c1 ;
 wire \V2/V3/A2/A1/M3/c2 ;
 wire \V2/V3/A2/A1/M3/s1 ;
 wire \V2/V3/A2/A1/M4/c1 ;
 wire \V2/V3/A2/A1/M4/c2 ;
 wire \V2/V3/A2/A1/M4/s1 ;
 wire \V2/V3/A2/A2/c1 ;
 wire \V2/V3/A2/A2/c2 ;
 wire \V2/V3/A2/A2/c3 ;
 wire \V2/V3/A2/A2/M1/c1 ;
 wire \V2/V3/A2/A2/M1/c2 ;
 wire \V2/V3/A2/A2/M1/s1 ;
 wire \V2/V3/A2/A2/M2/c1 ;
 wire \V2/V3/A2/A2/M2/c2 ;
 wire \V2/V3/A2/A2/M2/s1 ;
 wire \V2/V3/A2/A2/M3/c1 ;
 wire \V2/V3/A2/A2/M3/c2 ;
 wire \V2/V3/A2/A2/M3/s1 ;
 wire \V2/V3/A2/A2/M4/c1 ;
 wire \V2/V3/A2/A2/M4/c2 ;
 wire \V2/V3/A2/A2/M4/s1 ;
 wire \V2/V3/A3/c1 ;
 wire \V2/V3/A3/A1/c1 ;
 wire \V2/V3/A3/A1/c2 ;
 wire \V2/V3/A3/A1/c3 ;
 wire \V2/V3/A3/A1/M1/c1 ;
 wire \V2/V3/A3/A1/M1/c2 ;
 wire \V2/V3/A3/A1/M1/s1 ;
 wire \V2/V3/A3/A1/M2/c1 ;
 wire \V2/V3/A3/A1/M2/c2 ;
 wire \V2/V3/A3/A1/M2/s1 ;
 wire \V2/V3/A3/A1/M3/c1 ;
 wire \V2/V3/A3/A1/M3/c2 ;
 wire \V2/V3/A3/A1/M3/s1 ;
 wire \V2/V3/A3/A1/M4/c1 ;
 wire \V2/V3/A3/A1/M4/c2 ;
 wire \V2/V3/A3/A1/M4/s1 ;
 wire \V2/V3/A3/A2/c1 ;
 wire \V2/V3/A3/A2/c2 ;
 wire \V2/V3/A3/A2/c3 ;
 wire \V2/V3/A3/A2/M1/c1 ;
 wire \V2/V3/A3/A2/M1/c2 ;
 wire \V2/V3/A3/A2/M1/s1 ;
 wire \V2/V3/A3/A2/M2/c1 ;
 wire \V2/V3/A3/A2/M2/c2 ;
 wire \V2/V3/A3/A2/M2/s1 ;
 wire \V2/V3/A3/A2/M3/c1 ;
 wire \V2/V3/A3/A2/M3/c2 ;
 wire \V2/V3/A3/A2/M3/s1 ;
 wire \V2/V3/A3/A2/M4/c1 ;
 wire \V2/V3/A3/A2/M4/c2 ;
 wire \V2/V3/A3/A2/M4/s1 ;
 wire \V2/V3/V1/c1 ;
 wire \V2/V3/V1/c2 ;
 wire \V2/V3/V1/c3 ;
 wire \V2/V3/V1/overflow ;
 wire \V2/V3/V1/A1/c1 ;
 wire \V2/V3/V1/A1/c2 ;
 wire \V2/V3/V1/A1/c3 ;
 wire \V2/V3/V1/A1/M1/c1 ;
 wire \V2/V3/V1/A1/M1/c2 ;
 wire \V2/V3/V1/A1/M1/s1 ;
 wire \V2/V3/V1/A1/M2/c1 ;
 wire \V2/V3/V1/A1/M2/c2 ;
 wire \V2/V3/V1/A1/M2/s1 ;
 wire \V2/V3/V1/A1/M3/c1 ;
 wire \V2/V3/V1/A1/M3/c2 ;
 wire \V2/V3/V1/A1/M3/s1 ;
 wire \V2/V3/V1/A1/M4/c1 ;
 wire \V2/V3/V1/A1/M4/c2 ;
 wire \V2/V3/V1/A1/M4/s1 ;
 wire \V2/V3/V1/A2/c1 ;
 wire \V2/V3/V1/A2/c2 ;
 wire \V2/V3/V1/A2/c3 ;
 wire \V2/V3/V1/A2/M1/c1 ;
 wire \V2/V3/V1/A2/M1/c2 ;
 wire \V2/V3/V1/A2/M1/s1 ;
 wire \V2/V3/V1/A2/M2/c1 ;
 wire \V2/V3/V1/A2/M2/c2 ;
 wire \V2/V3/V1/A2/M2/s1 ;
 wire \V2/V3/V1/A2/M3/c1 ;
 wire \V2/V3/V1/A2/M3/c2 ;
 wire \V2/V3/V1/A2/M3/s1 ;
 wire \V2/V3/V1/A2/M4/c1 ;
 wire \V2/V3/V1/A2/M4/c2 ;
 wire \V2/V3/V1/A2/M4/s1 ;
 wire \V2/V3/V1/A3/c1 ;
 wire \V2/V3/V1/A3/c2 ;
 wire \V2/V3/V1/A3/c3 ;
 wire \V2/V3/V1/A3/M1/c1 ;
 wire \V2/V3/V1/A3/M1/c2 ;
 wire \V2/V3/V1/A3/M1/s1 ;
 wire \V2/V3/V1/A3/M2/c1 ;
 wire \V2/V3/V1/A3/M2/c2 ;
 wire \V2/V3/V1/A3/M2/s1 ;
 wire \V2/V3/V1/A3/M3/c1 ;
 wire \V2/V3/V1/A3/M3/c2 ;
 wire \V2/V3/V1/A3/M3/s1 ;
 wire \V2/V3/V1/A3/M4/c1 ;
 wire \V2/V3/V1/A3/M4/c2 ;
 wire \V2/V3/V1/A3/M4/s1 ;
 wire \V2/V3/V1/V1/w1 ;
 wire \V2/V3/V1/V1/w2 ;
 wire \V2/V3/V1/V1/w3 ;
 wire \V2/V3/V1/V1/w4 ;
 wire \V2/V3/V1/V2/w1 ;
 wire \V2/V3/V1/V2/w2 ;
 wire \V2/V3/V1/V2/w3 ;
 wire \V2/V3/V1/V2/w4 ;
 wire \V2/V3/V1/V3/w1 ;
 wire \V2/V3/V1/V3/w2 ;
 wire \V2/V3/V1/V3/w3 ;
 wire \V2/V3/V1/V3/w4 ;
 wire \V2/V3/V1/V4/w1 ;
 wire \V2/V3/V1/V4/w2 ;
 wire \V2/V3/V1/V4/w3 ;
 wire \V2/V3/V1/V4/w4 ;
 wire \V2/V3/V2/c1 ;
 wire \V2/V3/V2/c2 ;
 wire \V2/V3/V2/c3 ;
 wire \V2/V3/V2/overflow ;
 wire \V2/V3/V2/A1/c1 ;
 wire \V2/V3/V2/A1/c2 ;
 wire \V2/V3/V2/A1/c3 ;
 wire \V2/V3/V2/A1/M1/c1 ;
 wire \V2/V3/V2/A1/M1/c2 ;
 wire \V2/V3/V2/A1/M1/s1 ;
 wire \V2/V3/V2/A1/M2/c1 ;
 wire \V2/V3/V2/A1/M2/c2 ;
 wire \V2/V3/V2/A1/M2/s1 ;
 wire \V2/V3/V2/A1/M3/c1 ;
 wire \V2/V3/V2/A1/M3/c2 ;
 wire \V2/V3/V2/A1/M3/s1 ;
 wire \V2/V3/V2/A1/M4/c1 ;
 wire \V2/V3/V2/A1/M4/c2 ;
 wire \V2/V3/V2/A1/M4/s1 ;
 wire \V2/V3/V2/A2/c1 ;
 wire \V2/V3/V2/A2/c2 ;
 wire \V2/V3/V2/A2/c3 ;
 wire \V2/V3/V2/A2/M1/c1 ;
 wire \V2/V3/V2/A2/M1/c2 ;
 wire \V2/V3/V2/A2/M1/s1 ;
 wire \V2/V3/V2/A2/M2/c1 ;
 wire \V2/V3/V2/A2/M2/c2 ;
 wire \V2/V3/V2/A2/M2/s1 ;
 wire \V2/V3/V2/A2/M3/c1 ;
 wire \V2/V3/V2/A2/M3/c2 ;
 wire \V2/V3/V2/A2/M3/s1 ;
 wire \V2/V3/V2/A2/M4/c1 ;
 wire \V2/V3/V2/A2/M4/c2 ;
 wire \V2/V3/V2/A2/M4/s1 ;
 wire \V2/V3/V2/A3/c1 ;
 wire \V2/V3/V2/A3/c2 ;
 wire \V2/V3/V2/A3/c3 ;
 wire \V2/V3/V2/A3/M1/c1 ;
 wire \V2/V3/V2/A3/M1/c2 ;
 wire \V2/V3/V2/A3/M1/s1 ;
 wire \V2/V3/V2/A3/M2/c1 ;
 wire \V2/V3/V2/A3/M2/c2 ;
 wire \V2/V3/V2/A3/M2/s1 ;
 wire \V2/V3/V2/A3/M3/c1 ;
 wire \V2/V3/V2/A3/M3/c2 ;
 wire \V2/V3/V2/A3/M3/s1 ;
 wire \V2/V3/V2/A3/M4/c1 ;
 wire \V2/V3/V2/A3/M4/c2 ;
 wire \V2/V3/V2/A3/M4/s1 ;
 wire \V2/V3/V2/V1/w1 ;
 wire \V2/V3/V2/V1/w2 ;
 wire \V2/V3/V2/V1/w3 ;
 wire \V2/V3/V2/V1/w4 ;
 wire \V2/V3/V2/V2/w1 ;
 wire \V2/V3/V2/V2/w2 ;
 wire \V2/V3/V2/V2/w3 ;
 wire \V2/V3/V2/V2/w4 ;
 wire \V2/V3/V2/V3/w1 ;
 wire \V2/V3/V2/V3/w2 ;
 wire \V2/V3/V2/V3/w3 ;
 wire \V2/V3/V2/V3/w4 ;
 wire \V2/V3/V2/V4/w1 ;
 wire \V2/V3/V2/V4/w2 ;
 wire \V2/V3/V2/V4/w3 ;
 wire \V2/V3/V2/V4/w4 ;
 wire \V2/V3/V3/c1 ;
 wire \V2/V3/V3/c2 ;
 wire \V2/V3/V3/c3 ;
 wire \V2/V3/V3/overflow ;
 wire \V2/V3/V3/A1/c1 ;
 wire \V2/V3/V3/A1/c2 ;
 wire \V2/V3/V3/A1/c3 ;
 wire \V2/V3/V3/A1/M1/c1 ;
 wire \V2/V3/V3/A1/M1/c2 ;
 wire \V2/V3/V3/A1/M1/s1 ;
 wire \V2/V3/V3/A1/M2/c1 ;
 wire \V2/V3/V3/A1/M2/c2 ;
 wire \V2/V3/V3/A1/M2/s1 ;
 wire \V2/V3/V3/A1/M3/c1 ;
 wire \V2/V3/V3/A1/M3/c2 ;
 wire \V2/V3/V3/A1/M3/s1 ;
 wire \V2/V3/V3/A1/M4/c1 ;
 wire \V2/V3/V3/A1/M4/c2 ;
 wire \V2/V3/V3/A1/M4/s1 ;
 wire \V2/V3/V3/A2/c1 ;
 wire \V2/V3/V3/A2/c2 ;
 wire \V2/V3/V3/A2/c3 ;
 wire \V2/V3/V3/A2/M1/c1 ;
 wire \V2/V3/V3/A2/M1/c2 ;
 wire \V2/V3/V3/A2/M1/s1 ;
 wire \V2/V3/V3/A2/M2/c1 ;
 wire \V2/V3/V3/A2/M2/c2 ;
 wire \V2/V3/V3/A2/M2/s1 ;
 wire \V2/V3/V3/A2/M3/c1 ;
 wire \V2/V3/V3/A2/M3/c2 ;
 wire \V2/V3/V3/A2/M3/s1 ;
 wire \V2/V3/V3/A2/M4/c1 ;
 wire \V2/V3/V3/A2/M4/c2 ;
 wire \V2/V3/V3/A2/M4/s1 ;
 wire \V2/V3/V3/A3/c1 ;
 wire \V2/V3/V3/A3/c2 ;
 wire \V2/V3/V3/A3/c3 ;
 wire \V2/V3/V3/A3/M1/c1 ;
 wire \V2/V3/V3/A3/M1/c2 ;
 wire \V2/V3/V3/A3/M1/s1 ;
 wire \V2/V3/V3/A3/M2/c1 ;
 wire \V2/V3/V3/A3/M2/c2 ;
 wire \V2/V3/V3/A3/M2/s1 ;
 wire \V2/V3/V3/A3/M3/c1 ;
 wire \V2/V3/V3/A3/M3/c2 ;
 wire \V2/V3/V3/A3/M3/s1 ;
 wire \V2/V3/V3/A3/M4/c1 ;
 wire \V2/V3/V3/A3/M4/c2 ;
 wire \V2/V3/V3/A3/M4/s1 ;
 wire \V2/V3/V3/V1/w1 ;
 wire \V2/V3/V3/V1/w2 ;
 wire \V2/V3/V3/V1/w3 ;
 wire \V2/V3/V3/V1/w4 ;
 wire \V2/V3/V3/V2/w1 ;
 wire \V2/V3/V3/V2/w2 ;
 wire \V2/V3/V3/V2/w3 ;
 wire \V2/V3/V3/V2/w4 ;
 wire \V2/V3/V3/V3/w1 ;
 wire \V2/V3/V3/V3/w2 ;
 wire \V2/V3/V3/V3/w3 ;
 wire \V2/V3/V3/V3/w4 ;
 wire \V2/V3/V3/V4/w1 ;
 wire \V2/V3/V3/V4/w2 ;
 wire \V2/V3/V3/V4/w3 ;
 wire \V2/V3/V3/V4/w4 ;
 wire \V2/V3/V4/c1 ;
 wire \V2/V3/V4/c2 ;
 wire \V2/V3/V4/c3 ;
 wire \V2/V3/V4/overflow ;
 wire \V2/V3/V4/A1/c1 ;
 wire \V2/V3/V4/A1/c2 ;
 wire \V2/V3/V4/A1/c3 ;
 wire \V2/V3/V4/A1/M1/c1 ;
 wire \V2/V3/V4/A1/M1/c2 ;
 wire \V2/V3/V4/A1/M1/s1 ;
 wire \V2/V3/V4/A1/M2/c1 ;
 wire \V2/V3/V4/A1/M2/c2 ;
 wire \V2/V3/V4/A1/M2/s1 ;
 wire \V2/V3/V4/A1/M3/c1 ;
 wire \V2/V3/V4/A1/M3/c2 ;
 wire \V2/V3/V4/A1/M3/s1 ;
 wire \V2/V3/V4/A1/M4/c1 ;
 wire \V2/V3/V4/A1/M4/c2 ;
 wire \V2/V3/V4/A1/M4/s1 ;
 wire \V2/V3/V4/A2/c1 ;
 wire \V2/V3/V4/A2/c2 ;
 wire \V2/V3/V4/A2/c3 ;
 wire \V2/V3/V4/A2/M1/c1 ;
 wire \V2/V3/V4/A2/M1/c2 ;
 wire \V2/V3/V4/A2/M1/s1 ;
 wire \V2/V3/V4/A2/M2/c1 ;
 wire \V2/V3/V4/A2/M2/c2 ;
 wire \V2/V3/V4/A2/M2/s1 ;
 wire \V2/V3/V4/A2/M3/c1 ;
 wire \V2/V3/V4/A2/M3/c2 ;
 wire \V2/V3/V4/A2/M3/s1 ;
 wire \V2/V3/V4/A2/M4/c1 ;
 wire \V2/V3/V4/A2/M4/c2 ;
 wire \V2/V3/V4/A2/M4/s1 ;
 wire \V2/V3/V4/A3/c1 ;
 wire \V2/V3/V4/A3/c2 ;
 wire \V2/V3/V4/A3/c3 ;
 wire \V2/V3/V4/A3/M1/c1 ;
 wire \V2/V3/V4/A3/M1/c2 ;
 wire \V2/V3/V4/A3/M1/s1 ;
 wire \V2/V3/V4/A3/M2/c1 ;
 wire \V2/V3/V4/A3/M2/c2 ;
 wire \V2/V3/V4/A3/M2/s1 ;
 wire \V2/V3/V4/A3/M3/c1 ;
 wire \V2/V3/V4/A3/M3/c2 ;
 wire \V2/V3/V4/A3/M3/s1 ;
 wire \V2/V3/V4/A3/M4/c1 ;
 wire \V2/V3/V4/A3/M4/c2 ;
 wire \V2/V3/V4/A3/M4/s1 ;
 wire \V2/V3/V4/V1/w1 ;
 wire \V2/V3/V4/V1/w2 ;
 wire \V2/V3/V4/V1/w3 ;
 wire \V2/V3/V4/V1/w4 ;
 wire \V2/V3/V4/V2/w1 ;
 wire \V2/V3/V4/V2/w2 ;
 wire \V2/V3/V4/V2/w3 ;
 wire \V2/V3/V4/V2/w4 ;
 wire \V2/V3/V4/V3/w1 ;
 wire \V2/V3/V4/V3/w2 ;
 wire \V2/V3/V4/V3/w3 ;
 wire \V2/V3/V4/V3/w4 ;
 wire \V2/V3/V4/V4/w1 ;
 wire \V2/V3/V4/V4/w2 ;
 wire \V2/V3/V4/V4/w3 ;
 wire \V2/V3/V4/V4/w4 ;
 wire \V2/V4/c1 ;
 wire \V2/V4/c2 ;
 wire \V2/V4/c3 ;
 wire \V2/V4/overflow ;
 wire \V2/V4/A1/c1 ;
 wire \V2/V4/A1/A1/c1 ;
 wire \V2/V4/A1/A1/c2 ;
 wire \V2/V4/A1/A1/c3 ;
 wire \V2/V4/A1/A1/M1/c1 ;
 wire \V2/V4/A1/A1/M1/c2 ;
 wire \V2/V4/A1/A1/M1/s1 ;
 wire \V2/V4/A1/A1/M2/c1 ;
 wire \V2/V4/A1/A1/M2/c2 ;
 wire \V2/V4/A1/A1/M2/s1 ;
 wire \V2/V4/A1/A1/M3/c1 ;
 wire \V2/V4/A1/A1/M3/c2 ;
 wire \V2/V4/A1/A1/M3/s1 ;
 wire \V2/V4/A1/A1/M4/c1 ;
 wire \V2/V4/A1/A1/M4/c2 ;
 wire \V2/V4/A1/A1/M4/s1 ;
 wire \V2/V4/A1/A2/c1 ;
 wire \V2/V4/A1/A2/c2 ;
 wire \V2/V4/A1/A2/c3 ;
 wire \V2/V4/A1/A2/M1/c1 ;
 wire \V2/V4/A1/A2/M1/c2 ;
 wire \V2/V4/A1/A2/M1/s1 ;
 wire \V2/V4/A1/A2/M2/c1 ;
 wire \V2/V4/A1/A2/M2/c2 ;
 wire \V2/V4/A1/A2/M2/s1 ;
 wire \V2/V4/A1/A2/M3/c1 ;
 wire \V2/V4/A1/A2/M3/c2 ;
 wire \V2/V4/A1/A2/M3/s1 ;
 wire \V2/V4/A1/A2/M4/c1 ;
 wire \V2/V4/A1/A2/M4/c2 ;
 wire \V2/V4/A1/A2/M4/s1 ;
 wire \V2/V4/A2/c1 ;
 wire \V2/V4/A2/A1/c1 ;
 wire \V2/V4/A2/A1/c2 ;
 wire \V2/V4/A2/A1/c3 ;
 wire \V2/V4/A2/A1/M1/c1 ;
 wire \V2/V4/A2/A1/M1/c2 ;
 wire \V2/V4/A2/A1/M1/s1 ;
 wire \V2/V4/A2/A1/M2/c1 ;
 wire \V2/V4/A2/A1/M2/c2 ;
 wire \V2/V4/A2/A1/M2/s1 ;
 wire \V2/V4/A2/A1/M3/c1 ;
 wire \V2/V4/A2/A1/M3/c2 ;
 wire \V2/V4/A2/A1/M3/s1 ;
 wire \V2/V4/A2/A1/M4/c1 ;
 wire \V2/V4/A2/A1/M4/c2 ;
 wire \V2/V4/A2/A1/M4/s1 ;
 wire \V2/V4/A2/A2/c1 ;
 wire \V2/V4/A2/A2/c2 ;
 wire \V2/V4/A2/A2/c3 ;
 wire \V2/V4/A2/A2/M1/c1 ;
 wire \V2/V4/A2/A2/M1/c2 ;
 wire \V2/V4/A2/A2/M1/s1 ;
 wire \V2/V4/A2/A2/M2/c1 ;
 wire \V2/V4/A2/A2/M2/c2 ;
 wire \V2/V4/A2/A2/M2/s1 ;
 wire \V2/V4/A2/A2/M3/c1 ;
 wire \V2/V4/A2/A2/M3/c2 ;
 wire \V2/V4/A2/A2/M3/s1 ;
 wire \V2/V4/A2/A2/M4/c1 ;
 wire \V2/V4/A2/A2/M4/c2 ;
 wire \V2/V4/A2/A2/M4/s1 ;
 wire \V2/V4/A3/c1 ;
 wire \V2/V4/A3/A1/c1 ;
 wire \V2/V4/A3/A1/c2 ;
 wire \V2/V4/A3/A1/c3 ;
 wire \V2/V4/A3/A1/M1/c1 ;
 wire \V2/V4/A3/A1/M1/c2 ;
 wire \V2/V4/A3/A1/M1/s1 ;
 wire \V2/V4/A3/A1/M2/c1 ;
 wire \V2/V4/A3/A1/M2/c2 ;
 wire \V2/V4/A3/A1/M2/s1 ;
 wire \V2/V4/A3/A1/M3/c1 ;
 wire \V2/V4/A3/A1/M3/c2 ;
 wire \V2/V4/A3/A1/M3/s1 ;
 wire \V2/V4/A3/A1/M4/c1 ;
 wire \V2/V4/A3/A1/M4/c2 ;
 wire \V2/V4/A3/A1/M4/s1 ;
 wire \V2/V4/A3/A2/c1 ;
 wire \V2/V4/A3/A2/c2 ;
 wire \V2/V4/A3/A2/c3 ;
 wire \V2/V4/A3/A2/M1/c1 ;
 wire \V2/V4/A3/A2/M1/c2 ;
 wire \V2/V4/A3/A2/M1/s1 ;
 wire \V2/V4/A3/A2/M2/c1 ;
 wire \V2/V4/A3/A2/M2/c2 ;
 wire \V2/V4/A3/A2/M2/s1 ;
 wire \V2/V4/A3/A2/M3/c1 ;
 wire \V2/V4/A3/A2/M3/c2 ;
 wire \V2/V4/A3/A2/M3/s1 ;
 wire \V2/V4/A3/A2/M4/c1 ;
 wire \V2/V4/A3/A2/M4/c2 ;
 wire \V2/V4/A3/A2/M4/s1 ;
 wire \V2/V4/V1/c1 ;
 wire \V2/V4/V1/c2 ;
 wire \V2/V4/V1/c3 ;
 wire \V2/V4/V1/overflow ;
 wire \V2/V4/V1/A1/c1 ;
 wire \V2/V4/V1/A1/c2 ;
 wire \V2/V4/V1/A1/c3 ;
 wire \V2/V4/V1/A1/M1/c1 ;
 wire \V2/V4/V1/A1/M1/c2 ;
 wire \V2/V4/V1/A1/M1/s1 ;
 wire \V2/V4/V1/A1/M2/c1 ;
 wire \V2/V4/V1/A1/M2/c2 ;
 wire \V2/V4/V1/A1/M2/s1 ;
 wire \V2/V4/V1/A1/M3/c1 ;
 wire \V2/V4/V1/A1/M3/c2 ;
 wire \V2/V4/V1/A1/M3/s1 ;
 wire \V2/V4/V1/A1/M4/c1 ;
 wire \V2/V4/V1/A1/M4/c2 ;
 wire \V2/V4/V1/A1/M4/s1 ;
 wire \V2/V4/V1/A2/c1 ;
 wire \V2/V4/V1/A2/c2 ;
 wire \V2/V4/V1/A2/c3 ;
 wire \V2/V4/V1/A2/M1/c1 ;
 wire \V2/V4/V1/A2/M1/c2 ;
 wire \V2/V4/V1/A2/M1/s1 ;
 wire \V2/V4/V1/A2/M2/c1 ;
 wire \V2/V4/V1/A2/M2/c2 ;
 wire \V2/V4/V1/A2/M2/s1 ;
 wire \V2/V4/V1/A2/M3/c1 ;
 wire \V2/V4/V1/A2/M3/c2 ;
 wire \V2/V4/V1/A2/M3/s1 ;
 wire \V2/V4/V1/A2/M4/c1 ;
 wire \V2/V4/V1/A2/M4/c2 ;
 wire \V2/V4/V1/A2/M4/s1 ;
 wire \V2/V4/V1/A3/c1 ;
 wire \V2/V4/V1/A3/c2 ;
 wire \V2/V4/V1/A3/c3 ;
 wire \V2/V4/V1/A3/M1/c1 ;
 wire \V2/V4/V1/A3/M1/c2 ;
 wire \V2/V4/V1/A3/M1/s1 ;
 wire \V2/V4/V1/A3/M2/c1 ;
 wire \V2/V4/V1/A3/M2/c2 ;
 wire \V2/V4/V1/A3/M2/s1 ;
 wire \V2/V4/V1/A3/M3/c1 ;
 wire \V2/V4/V1/A3/M3/c2 ;
 wire \V2/V4/V1/A3/M3/s1 ;
 wire \V2/V4/V1/A3/M4/c1 ;
 wire \V2/V4/V1/A3/M4/c2 ;
 wire \V2/V4/V1/A3/M4/s1 ;
 wire \V2/V4/V1/V1/w1 ;
 wire \V2/V4/V1/V1/w2 ;
 wire \V2/V4/V1/V1/w3 ;
 wire \V2/V4/V1/V1/w4 ;
 wire \V2/V4/V1/V2/w1 ;
 wire \V2/V4/V1/V2/w2 ;
 wire \V2/V4/V1/V2/w3 ;
 wire \V2/V4/V1/V2/w4 ;
 wire \V2/V4/V1/V3/w1 ;
 wire \V2/V4/V1/V3/w2 ;
 wire \V2/V4/V1/V3/w3 ;
 wire \V2/V4/V1/V3/w4 ;
 wire \V2/V4/V1/V4/w1 ;
 wire \V2/V4/V1/V4/w2 ;
 wire \V2/V4/V1/V4/w3 ;
 wire \V2/V4/V1/V4/w4 ;
 wire \V2/V4/V2/c1 ;
 wire \V2/V4/V2/c2 ;
 wire \V2/V4/V2/c3 ;
 wire \V2/V4/V2/overflow ;
 wire \V2/V4/V2/A1/c1 ;
 wire \V2/V4/V2/A1/c2 ;
 wire \V2/V4/V2/A1/c3 ;
 wire \V2/V4/V2/A1/M1/c1 ;
 wire \V2/V4/V2/A1/M1/c2 ;
 wire \V2/V4/V2/A1/M1/s1 ;
 wire \V2/V4/V2/A1/M2/c1 ;
 wire \V2/V4/V2/A1/M2/c2 ;
 wire \V2/V4/V2/A1/M2/s1 ;
 wire \V2/V4/V2/A1/M3/c1 ;
 wire \V2/V4/V2/A1/M3/c2 ;
 wire \V2/V4/V2/A1/M3/s1 ;
 wire \V2/V4/V2/A1/M4/c1 ;
 wire \V2/V4/V2/A1/M4/c2 ;
 wire \V2/V4/V2/A1/M4/s1 ;
 wire \V2/V4/V2/A2/c1 ;
 wire \V2/V4/V2/A2/c2 ;
 wire \V2/V4/V2/A2/c3 ;
 wire \V2/V4/V2/A2/M1/c1 ;
 wire \V2/V4/V2/A2/M1/c2 ;
 wire \V2/V4/V2/A2/M1/s1 ;
 wire \V2/V4/V2/A2/M2/c1 ;
 wire \V2/V4/V2/A2/M2/c2 ;
 wire \V2/V4/V2/A2/M2/s1 ;
 wire \V2/V4/V2/A2/M3/c1 ;
 wire \V2/V4/V2/A2/M3/c2 ;
 wire \V2/V4/V2/A2/M3/s1 ;
 wire \V2/V4/V2/A2/M4/c1 ;
 wire \V2/V4/V2/A2/M4/c2 ;
 wire \V2/V4/V2/A2/M4/s1 ;
 wire \V2/V4/V2/A3/c1 ;
 wire \V2/V4/V2/A3/c2 ;
 wire \V2/V4/V2/A3/c3 ;
 wire \V2/V4/V2/A3/M1/c1 ;
 wire \V2/V4/V2/A3/M1/c2 ;
 wire \V2/V4/V2/A3/M1/s1 ;
 wire \V2/V4/V2/A3/M2/c1 ;
 wire \V2/V4/V2/A3/M2/c2 ;
 wire \V2/V4/V2/A3/M2/s1 ;
 wire \V2/V4/V2/A3/M3/c1 ;
 wire \V2/V4/V2/A3/M3/c2 ;
 wire \V2/V4/V2/A3/M3/s1 ;
 wire \V2/V4/V2/A3/M4/c1 ;
 wire \V2/V4/V2/A3/M4/c2 ;
 wire \V2/V4/V2/A3/M4/s1 ;
 wire \V2/V4/V2/V1/w1 ;
 wire \V2/V4/V2/V1/w2 ;
 wire \V2/V4/V2/V1/w3 ;
 wire \V2/V4/V2/V1/w4 ;
 wire \V2/V4/V2/V2/w1 ;
 wire \V2/V4/V2/V2/w2 ;
 wire \V2/V4/V2/V2/w3 ;
 wire \V2/V4/V2/V2/w4 ;
 wire \V2/V4/V2/V3/w1 ;
 wire \V2/V4/V2/V3/w2 ;
 wire \V2/V4/V2/V3/w3 ;
 wire \V2/V4/V2/V3/w4 ;
 wire \V2/V4/V2/V4/w1 ;
 wire \V2/V4/V2/V4/w2 ;
 wire \V2/V4/V2/V4/w3 ;
 wire \V2/V4/V2/V4/w4 ;
 wire \V2/V4/V3/c1 ;
 wire \V2/V4/V3/c2 ;
 wire \V2/V4/V3/c3 ;
 wire \V2/V4/V3/overflow ;
 wire \V2/V4/V3/A1/c1 ;
 wire \V2/V4/V3/A1/c2 ;
 wire \V2/V4/V3/A1/c3 ;
 wire \V2/V4/V3/A1/M1/c1 ;
 wire \V2/V4/V3/A1/M1/c2 ;
 wire \V2/V4/V3/A1/M1/s1 ;
 wire \V2/V4/V3/A1/M2/c1 ;
 wire \V2/V4/V3/A1/M2/c2 ;
 wire \V2/V4/V3/A1/M2/s1 ;
 wire \V2/V4/V3/A1/M3/c1 ;
 wire \V2/V4/V3/A1/M3/c2 ;
 wire \V2/V4/V3/A1/M3/s1 ;
 wire \V2/V4/V3/A1/M4/c1 ;
 wire \V2/V4/V3/A1/M4/c2 ;
 wire \V2/V4/V3/A1/M4/s1 ;
 wire \V2/V4/V3/A2/c1 ;
 wire \V2/V4/V3/A2/c2 ;
 wire \V2/V4/V3/A2/c3 ;
 wire \V2/V4/V3/A2/M1/c1 ;
 wire \V2/V4/V3/A2/M1/c2 ;
 wire \V2/V4/V3/A2/M1/s1 ;
 wire \V2/V4/V3/A2/M2/c1 ;
 wire \V2/V4/V3/A2/M2/c2 ;
 wire \V2/V4/V3/A2/M2/s1 ;
 wire \V2/V4/V3/A2/M3/c1 ;
 wire \V2/V4/V3/A2/M3/c2 ;
 wire \V2/V4/V3/A2/M3/s1 ;
 wire \V2/V4/V3/A2/M4/c1 ;
 wire \V2/V4/V3/A2/M4/c2 ;
 wire \V2/V4/V3/A2/M4/s1 ;
 wire \V2/V4/V3/A3/c1 ;
 wire \V2/V4/V3/A3/c2 ;
 wire \V2/V4/V3/A3/c3 ;
 wire \V2/V4/V3/A3/M1/c1 ;
 wire \V2/V4/V3/A3/M1/c2 ;
 wire \V2/V4/V3/A3/M1/s1 ;
 wire \V2/V4/V3/A3/M2/c1 ;
 wire \V2/V4/V3/A3/M2/c2 ;
 wire \V2/V4/V3/A3/M2/s1 ;
 wire \V2/V4/V3/A3/M3/c1 ;
 wire \V2/V4/V3/A3/M3/c2 ;
 wire \V2/V4/V3/A3/M3/s1 ;
 wire \V2/V4/V3/A3/M4/c1 ;
 wire \V2/V4/V3/A3/M4/c2 ;
 wire \V2/V4/V3/A3/M4/s1 ;
 wire \V2/V4/V3/V1/w1 ;
 wire \V2/V4/V3/V1/w2 ;
 wire \V2/V4/V3/V1/w3 ;
 wire \V2/V4/V3/V1/w4 ;
 wire \V2/V4/V3/V2/w1 ;
 wire \V2/V4/V3/V2/w2 ;
 wire \V2/V4/V3/V2/w3 ;
 wire \V2/V4/V3/V2/w4 ;
 wire \V2/V4/V3/V3/w1 ;
 wire \V2/V4/V3/V3/w2 ;
 wire \V2/V4/V3/V3/w3 ;
 wire \V2/V4/V3/V3/w4 ;
 wire \V2/V4/V3/V4/w1 ;
 wire \V2/V4/V3/V4/w2 ;
 wire \V2/V4/V3/V4/w3 ;
 wire \V2/V4/V3/V4/w4 ;
 wire \V2/V4/V4/c1 ;
 wire \V2/V4/V4/c2 ;
 wire \V2/V4/V4/c3 ;
 wire \V2/V4/V4/overflow ;
 wire \V2/V4/V4/A1/c1 ;
 wire \V2/V4/V4/A1/c2 ;
 wire \V2/V4/V4/A1/c3 ;
 wire \V2/V4/V4/A1/M1/c1 ;
 wire \V2/V4/V4/A1/M1/c2 ;
 wire \V2/V4/V4/A1/M1/s1 ;
 wire \V2/V4/V4/A1/M2/c1 ;
 wire \V2/V4/V4/A1/M2/c2 ;
 wire \V2/V4/V4/A1/M2/s1 ;
 wire \V2/V4/V4/A1/M3/c1 ;
 wire \V2/V4/V4/A1/M3/c2 ;
 wire \V2/V4/V4/A1/M3/s1 ;
 wire \V2/V4/V4/A1/M4/c1 ;
 wire \V2/V4/V4/A1/M4/c2 ;
 wire \V2/V4/V4/A1/M4/s1 ;
 wire \V2/V4/V4/A2/c1 ;
 wire \V2/V4/V4/A2/c2 ;
 wire \V2/V4/V4/A2/c3 ;
 wire \V2/V4/V4/A2/M1/c1 ;
 wire \V2/V4/V4/A2/M1/c2 ;
 wire \V2/V4/V4/A2/M1/s1 ;
 wire \V2/V4/V4/A2/M2/c1 ;
 wire \V2/V4/V4/A2/M2/c2 ;
 wire \V2/V4/V4/A2/M2/s1 ;
 wire \V2/V4/V4/A2/M3/c1 ;
 wire \V2/V4/V4/A2/M3/c2 ;
 wire \V2/V4/V4/A2/M3/s1 ;
 wire \V2/V4/V4/A2/M4/c1 ;
 wire \V2/V4/V4/A2/M4/c2 ;
 wire \V2/V4/V4/A2/M4/s1 ;
 wire \V2/V4/V4/A3/c1 ;
 wire \V2/V4/V4/A3/c2 ;
 wire \V2/V4/V4/A3/c3 ;
 wire \V2/V4/V4/A3/M1/c1 ;
 wire \V2/V4/V4/A3/M1/c2 ;
 wire \V2/V4/V4/A3/M1/s1 ;
 wire \V2/V4/V4/A3/M2/c1 ;
 wire \V2/V4/V4/A3/M2/c2 ;
 wire \V2/V4/V4/A3/M2/s1 ;
 wire \V2/V4/V4/A3/M3/c1 ;
 wire \V2/V4/V4/A3/M3/c2 ;
 wire \V2/V4/V4/A3/M3/s1 ;
 wire \V2/V4/V4/A3/M4/c1 ;
 wire \V2/V4/V4/A3/M4/c2 ;
 wire \V2/V4/V4/A3/M4/s1 ;
 wire \V2/V4/V4/V1/w1 ;
 wire \V2/V4/V4/V1/w2 ;
 wire \V2/V4/V4/V1/w3 ;
 wire \V2/V4/V4/V1/w4 ;
 wire \V2/V4/V4/V2/w1 ;
 wire \V2/V4/V4/V2/w2 ;
 wire \V2/V4/V4/V2/w3 ;
 wire \V2/V4/V4/V2/w4 ;
 wire \V2/V4/V4/V3/w1 ;
 wire \V2/V4/V4/V3/w2 ;
 wire \V2/V4/V4/V3/w3 ;
 wire \V2/V4/V4/V3/w4 ;
 wire \V2/V4/V4/V4/w1 ;
 wire \V2/V4/V4/V4/w2 ;
 wire \V2/V4/V4/V4/w3 ;
 wire \V2/V4/V4/V4/w4 ;
 wire \V3/c1 ;
 wire \V3/c2 ;
 wire \V3/c3 ;
 wire \V3/overflow ;
 wire \V3/A1/c1 ;
 wire \V3/A1/A1/c1 ;
 wire \V3/A1/A1/A1/c1 ;
 wire \V3/A1/A1/A1/c2 ;
 wire \V3/A1/A1/A1/c3 ;
 wire \V3/A1/A1/A1/M1/c1 ;
 wire \V3/A1/A1/A1/M1/c2 ;
 wire \V3/A1/A1/A1/M1/s1 ;
 wire \V3/A1/A1/A1/M2/c1 ;
 wire \V3/A1/A1/A1/M2/c2 ;
 wire \V3/A1/A1/A1/M2/s1 ;
 wire \V3/A1/A1/A1/M3/c1 ;
 wire \V3/A1/A1/A1/M3/c2 ;
 wire \V3/A1/A1/A1/M3/s1 ;
 wire \V3/A1/A1/A1/M4/c1 ;
 wire \V3/A1/A1/A1/M4/c2 ;
 wire \V3/A1/A1/A1/M4/s1 ;
 wire \V3/A1/A1/A2/c1 ;
 wire \V3/A1/A1/A2/c2 ;
 wire \V3/A1/A1/A2/c3 ;
 wire \V3/A1/A1/A2/M1/c1 ;
 wire \V3/A1/A1/A2/M1/c2 ;
 wire \V3/A1/A1/A2/M1/s1 ;
 wire \V3/A1/A1/A2/M2/c1 ;
 wire \V3/A1/A1/A2/M2/c2 ;
 wire \V3/A1/A1/A2/M2/s1 ;
 wire \V3/A1/A1/A2/M3/c1 ;
 wire \V3/A1/A1/A2/M3/c2 ;
 wire \V3/A1/A1/A2/M3/s1 ;
 wire \V3/A1/A1/A2/M4/c1 ;
 wire \V3/A1/A1/A2/M4/c2 ;
 wire \V3/A1/A1/A2/M4/s1 ;
 wire \V3/A1/A2/c1 ;
 wire \V3/A1/A2/A1/c1 ;
 wire \V3/A1/A2/A1/c2 ;
 wire \V3/A1/A2/A1/c3 ;
 wire \V3/A1/A2/A1/M1/c1 ;
 wire \V3/A1/A2/A1/M1/c2 ;
 wire \V3/A1/A2/A1/M1/s1 ;
 wire \V3/A1/A2/A1/M2/c1 ;
 wire \V3/A1/A2/A1/M2/c2 ;
 wire \V3/A1/A2/A1/M2/s1 ;
 wire \V3/A1/A2/A1/M3/c1 ;
 wire \V3/A1/A2/A1/M3/c2 ;
 wire \V3/A1/A2/A1/M3/s1 ;
 wire \V3/A1/A2/A1/M4/c1 ;
 wire \V3/A1/A2/A1/M4/c2 ;
 wire \V3/A1/A2/A1/M4/s1 ;
 wire \V3/A1/A2/A2/c1 ;
 wire \V3/A1/A2/A2/c2 ;
 wire \V3/A1/A2/A2/c3 ;
 wire \V3/A1/A2/A2/M1/c1 ;
 wire \V3/A1/A2/A2/M1/c2 ;
 wire \V3/A1/A2/A2/M1/s1 ;
 wire \V3/A1/A2/A2/M2/c1 ;
 wire \V3/A1/A2/A2/M2/c2 ;
 wire \V3/A1/A2/A2/M2/s1 ;
 wire \V3/A1/A2/A2/M3/c1 ;
 wire \V3/A1/A2/A2/M3/c2 ;
 wire \V3/A1/A2/A2/M3/s1 ;
 wire \V3/A1/A2/A2/M4/c1 ;
 wire \V3/A1/A2/A2/M4/c2 ;
 wire \V3/A1/A2/A2/M4/s1 ;
 wire \V3/A2/c1 ;
 wire \V3/A2/A1/c1 ;
 wire \V3/A2/A1/A1/c1 ;
 wire \V3/A2/A1/A1/c2 ;
 wire \V3/A2/A1/A1/c3 ;
 wire \V3/A2/A1/A1/M1/c1 ;
 wire \V3/A2/A1/A1/M1/c2 ;
 wire \V3/A2/A1/A1/M1/s1 ;
 wire \V3/A2/A1/A1/M2/c1 ;
 wire \V3/A2/A1/A1/M2/c2 ;
 wire \V3/A2/A1/A1/M2/s1 ;
 wire \V3/A2/A1/A1/M3/c1 ;
 wire \V3/A2/A1/A1/M3/c2 ;
 wire \V3/A2/A1/A1/M3/s1 ;
 wire \V3/A2/A1/A1/M4/c1 ;
 wire \V3/A2/A1/A1/M4/c2 ;
 wire \V3/A2/A1/A1/M4/s1 ;
 wire \V3/A2/A1/A2/c1 ;
 wire \V3/A2/A1/A2/c2 ;
 wire \V3/A2/A1/A2/c3 ;
 wire \V3/A2/A1/A2/M1/c1 ;
 wire \V3/A2/A1/A2/M1/c2 ;
 wire \V3/A2/A1/A2/M1/s1 ;
 wire \V3/A2/A1/A2/M2/c1 ;
 wire \V3/A2/A1/A2/M2/c2 ;
 wire \V3/A2/A1/A2/M2/s1 ;
 wire \V3/A2/A1/A2/M3/c1 ;
 wire \V3/A2/A1/A2/M3/c2 ;
 wire \V3/A2/A1/A2/M3/s1 ;
 wire \V3/A2/A1/A2/M4/c1 ;
 wire \V3/A2/A1/A2/M4/c2 ;
 wire \V3/A2/A1/A2/M4/s1 ;
 wire \V3/A2/A2/c1 ;
 wire \V3/A2/A2/A1/c1 ;
 wire \V3/A2/A2/A1/c2 ;
 wire \V3/A2/A2/A1/c3 ;
 wire \V3/A2/A2/A1/M1/c1 ;
 wire \V3/A2/A2/A1/M1/c2 ;
 wire \V3/A2/A2/A1/M1/s1 ;
 wire \V3/A2/A2/A1/M2/c1 ;
 wire \V3/A2/A2/A1/M2/c2 ;
 wire \V3/A2/A2/A1/M2/s1 ;
 wire \V3/A2/A2/A1/M3/c1 ;
 wire \V3/A2/A2/A1/M3/c2 ;
 wire \V3/A2/A2/A1/M3/s1 ;
 wire \V3/A2/A2/A1/M4/c1 ;
 wire \V3/A2/A2/A1/M4/c2 ;
 wire \V3/A2/A2/A1/M4/s1 ;
 wire \V3/A2/A2/A2/c1 ;
 wire \V3/A2/A2/A2/c2 ;
 wire \V3/A2/A2/A2/c3 ;
 wire \V3/A2/A2/A2/M1/c1 ;
 wire \V3/A2/A2/A2/M1/c2 ;
 wire \V3/A2/A2/A2/M1/s1 ;
 wire \V3/A2/A2/A2/M2/c1 ;
 wire \V3/A2/A2/A2/M2/c2 ;
 wire \V3/A2/A2/A2/M2/s1 ;
 wire \V3/A2/A2/A2/M3/c1 ;
 wire \V3/A2/A2/A2/M3/c2 ;
 wire \V3/A2/A2/A2/M3/s1 ;
 wire \V3/A2/A2/A2/M4/c1 ;
 wire \V3/A2/A2/A2/M4/c2 ;
 wire \V3/A2/A2/A2/M4/s1 ;
 wire \V3/A3/c1 ;
 wire \V3/A3/A1/c1 ;
 wire \V3/A3/A1/A1/c1 ;
 wire \V3/A3/A1/A1/c2 ;
 wire \V3/A3/A1/A1/c3 ;
 wire \V3/A3/A1/A1/M1/c1 ;
 wire \V3/A3/A1/A1/M1/c2 ;
 wire \V3/A3/A1/A1/M1/s1 ;
 wire \V3/A3/A1/A1/M2/c1 ;
 wire \V3/A3/A1/A1/M2/c2 ;
 wire \V3/A3/A1/A1/M2/s1 ;
 wire \V3/A3/A1/A1/M3/c1 ;
 wire \V3/A3/A1/A1/M3/c2 ;
 wire \V3/A3/A1/A1/M3/s1 ;
 wire \V3/A3/A1/A1/M4/c1 ;
 wire \V3/A3/A1/A1/M4/c2 ;
 wire \V3/A3/A1/A1/M4/s1 ;
 wire \V3/A3/A1/A2/c1 ;
 wire \V3/A3/A1/A2/c2 ;
 wire \V3/A3/A1/A2/c3 ;
 wire \V3/A3/A1/A2/M1/c1 ;
 wire \V3/A3/A1/A2/M1/c2 ;
 wire \V3/A3/A1/A2/M1/s1 ;
 wire \V3/A3/A1/A2/M2/c1 ;
 wire \V3/A3/A1/A2/M2/c2 ;
 wire \V3/A3/A1/A2/M2/s1 ;
 wire \V3/A3/A1/A2/M3/c1 ;
 wire \V3/A3/A1/A2/M3/c2 ;
 wire \V3/A3/A1/A2/M3/s1 ;
 wire \V3/A3/A1/A2/M4/c1 ;
 wire \V3/A3/A1/A2/M4/c2 ;
 wire \V3/A3/A1/A2/M4/s1 ;
 wire \V3/A3/A2/c1 ;
 wire \V3/A3/A2/A1/c1 ;
 wire \V3/A3/A2/A1/c2 ;
 wire \V3/A3/A2/A1/c3 ;
 wire \V3/A3/A2/A1/M1/c1 ;
 wire \V3/A3/A2/A1/M1/c2 ;
 wire \V3/A3/A2/A1/M1/s1 ;
 wire \V3/A3/A2/A1/M2/c1 ;
 wire \V3/A3/A2/A1/M2/c2 ;
 wire \V3/A3/A2/A1/M2/s1 ;
 wire \V3/A3/A2/A1/M3/c1 ;
 wire \V3/A3/A2/A1/M3/c2 ;
 wire \V3/A3/A2/A1/M3/s1 ;
 wire \V3/A3/A2/A1/M4/c1 ;
 wire \V3/A3/A2/A1/M4/c2 ;
 wire \V3/A3/A2/A1/M4/s1 ;
 wire \V3/A3/A2/A2/c1 ;
 wire \V3/A3/A2/A2/c2 ;
 wire \V3/A3/A2/A2/c3 ;
 wire \V3/A3/A2/A2/M1/c1 ;
 wire \V3/A3/A2/A2/M1/c2 ;
 wire \V3/A3/A2/A2/M1/s1 ;
 wire \V3/A3/A2/A2/M2/c1 ;
 wire \V3/A3/A2/A2/M2/c2 ;
 wire \V3/A3/A2/A2/M2/s1 ;
 wire \V3/A3/A2/A2/M3/c1 ;
 wire \V3/A3/A2/A2/M3/c2 ;
 wire \V3/A3/A2/A2/M3/s1 ;
 wire \V3/A3/A2/A2/M4/c1 ;
 wire \V3/A3/A2/A2/M4/c2 ;
 wire \V3/A3/A2/A2/M4/s1 ;
 wire \V3/V1/c1 ;
 wire \V3/V1/c2 ;
 wire \V3/V1/c3 ;
 wire \V3/V1/overflow ;
 wire \V3/V1/A1/c1 ;
 wire \V3/V1/A1/A1/c1 ;
 wire \V3/V1/A1/A1/c2 ;
 wire \V3/V1/A1/A1/c3 ;
 wire \V3/V1/A1/A1/M1/c1 ;
 wire \V3/V1/A1/A1/M1/c2 ;
 wire \V3/V1/A1/A1/M1/s1 ;
 wire \V3/V1/A1/A1/M2/c1 ;
 wire \V3/V1/A1/A1/M2/c2 ;
 wire \V3/V1/A1/A1/M2/s1 ;
 wire \V3/V1/A1/A1/M3/c1 ;
 wire \V3/V1/A1/A1/M3/c2 ;
 wire \V3/V1/A1/A1/M3/s1 ;
 wire \V3/V1/A1/A1/M4/c1 ;
 wire \V3/V1/A1/A1/M4/c2 ;
 wire \V3/V1/A1/A1/M4/s1 ;
 wire \V3/V1/A1/A2/c1 ;
 wire \V3/V1/A1/A2/c2 ;
 wire \V3/V1/A1/A2/c3 ;
 wire \V3/V1/A1/A2/M1/c1 ;
 wire \V3/V1/A1/A2/M1/c2 ;
 wire \V3/V1/A1/A2/M1/s1 ;
 wire \V3/V1/A1/A2/M2/c1 ;
 wire \V3/V1/A1/A2/M2/c2 ;
 wire \V3/V1/A1/A2/M2/s1 ;
 wire \V3/V1/A1/A2/M3/c1 ;
 wire \V3/V1/A1/A2/M3/c2 ;
 wire \V3/V1/A1/A2/M3/s1 ;
 wire \V3/V1/A1/A2/M4/c1 ;
 wire \V3/V1/A1/A2/M4/c2 ;
 wire \V3/V1/A1/A2/M4/s1 ;
 wire \V3/V1/A2/c1 ;
 wire \V3/V1/A2/A1/c1 ;
 wire \V3/V1/A2/A1/c2 ;
 wire \V3/V1/A2/A1/c3 ;
 wire \V3/V1/A2/A1/M1/c1 ;
 wire \V3/V1/A2/A1/M1/c2 ;
 wire \V3/V1/A2/A1/M1/s1 ;
 wire \V3/V1/A2/A1/M2/c1 ;
 wire \V3/V1/A2/A1/M2/c2 ;
 wire \V3/V1/A2/A1/M2/s1 ;
 wire \V3/V1/A2/A1/M3/c1 ;
 wire \V3/V1/A2/A1/M3/c2 ;
 wire \V3/V1/A2/A1/M3/s1 ;
 wire \V3/V1/A2/A1/M4/c1 ;
 wire \V3/V1/A2/A1/M4/c2 ;
 wire \V3/V1/A2/A1/M4/s1 ;
 wire \V3/V1/A2/A2/c1 ;
 wire \V3/V1/A2/A2/c2 ;
 wire \V3/V1/A2/A2/c3 ;
 wire \V3/V1/A2/A2/M1/c1 ;
 wire \V3/V1/A2/A2/M1/c2 ;
 wire \V3/V1/A2/A2/M1/s1 ;
 wire \V3/V1/A2/A2/M2/c1 ;
 wire \V3/V1/A2/A2/M2/c2 ;
 wire \V3/V1/A2/A2/M2/s1 ;
 wire \V3/V1/A2/A2/M3/c1 ;
 wire \V3/V1/A2/A2/M3/c2 ;
 wire \V3/V1/A2/A2/M3/s1 ;
 wire \V3/V1/A2/A2/M4/c1 ;
 wire \V3/V1/A2/A2/M4/c2 ;
 wire \V3/V1/A2/A2/M4/s1 ;
 wire \V3/V1/A3/c1 ;
 wire \V3/V1/A3/A1/c1 ;
 wire \V3/V1/A3/A1/c2 ;
 wire \V3/V1/A3/A1/c3 ;
 wire \V3/V1/A3/A1/M1/c1 ;
 wire \V3/V1/A3/A1/M1/c2 ;
 wire \V3/V1/A3/A1/M1/s1 ;
 wire \V3/V1/A3/A1/M2/c1 ;
 wire \V3/V1/A3/A1/M2/c2 ;
 wire \V3/V1/A3/A1/M2/s1 ;
 wire \V3/V1/A3/A1/M3/c1 ;
 wire \V3/V1/A3/A1/M3/c2 ;
 wire \V3/V1/A3/A1/M3/s1 ;
 wire \V3/V1/A3/A1/M4/c1 ;
 wire \V3/V1/A3/A1/M4/c2 ;
 wire \V3/V1/A3/A1/M4/s1 ;
 wire \V3/V1/A3/A2/c1 ;
 wire \V3/V1/A3/A2/c2 ;
 wire \V3/V1/A3/A2/c3 ;
 wire \V3/V1/A3/A2/M1/c1 ;
 wire \V3/V1/A3/A2/M1/c2 ;
 wire \V3/V1/A3/A2/M1/s1 ;
 wire \V3/V1/A3/A2/M2/c1 ;
 wire \V3/V1/A3/A2/M2/c2 ;
 wire \V3/V1/A3/A2/M2/s1 ;
 wire \V3/V1/A3/A2/M3/c1 ;
 wire \V3/V1/A3/A2/M3/c2 ;
 wire \V3/V1/A3/A2/M3/s1 ;
 wire \V3/V1/A3/A2/M4/c1 ;
 wire \V3/V1/A3/A2/M4/c2 ;
 wire \V3/V1/A3/A2/M4/s1 ;
 wire \V3/V1/V1/c1 ;
 wire \V3/V1/V1/c2 ;
 wire \V3/V1/V1/c3 ;
 wire \V3/V1/V1/overflow ;
 wire \V3/V1/V1/A1/c1 ;
 wire \V3/V1/V1/A1/c2 ;
 wire \V3/V1/V1/A1/c3 ;
 wire \V3/V1/V1/A1/M1/c1 ;
 wire \V3/V1/V1/A1/M1/c2 ;
 wire \V3/V1/V1/A1/M1/s1 ;
 wire \V3/V1/V1/A1/M2/c1 ;
 wire \V3/V1/V1/A1/M2/c2 ;
 wire \V3/V1/V1/A1/M2/s1 ;
 wire \V3/V1/V1/A1/M3/c1 ;
 wire \V3/V1/V1/A1/M3/c2 ;
 wire \V3/V1/V1/A1/M3/s1 ;
 wire \V3/V1/V1/A1/M4/c1 ;
 wire \V3/V1/V1/A1/M4/c2 ;
 wire \V3/V1/V1/A1/M4/s1 ;
 wire \V3/V1/V1/A2/c1 ;
 wire \V3/V1/V1/A2/c2 ;
 wire \V3/V1/V1/A2/c3 ;
 wire \V3/V1/V1/A2/M1/c1 ;
 wire \V3/V1/V1/A2/M1/c2 ;
 wire \V3/V1/V1/A2/M1/s1 ;
 wire \V3/V1/V1/A2/M2/c1 ;
 wire \V3/V1/V1/A2/M2/c2 ;
 wire \V3/V1/V1/A2/M2/s1 ;
 wire \V3/V1/V1/A2/M3/c1 ;
 wire \V3/V1/V1/A2/M3/c2 ;
 wire \V3/V1/V1/A2/M3/s1 ;
 wire \V3/V1/V1/A2/M4/c1 ;
 wire \V3/V1/V1/A2/M4/c2 ;
 wire \V3/V1/V1/A2/M4/s1 ;
 wire \V3/V1/V1/A3/c1 ;
 wire \V3/V1/V1/A3/c2 ;
 wire \V3/V1/V1/A3/c3 ;
 wire \V3/V1/V1/A3/M1/c1 ;
 wire \V3/V1/V1/A3/M1/c2 ;
 wire \V3/V1/V1/A3/M1/s1 ;
 wire \V3/V1/V1/A3/M2/c1 ;
 wire \V3/V1/V1/A3/M2/c2 ;
 wire \V3/V1/V1/A3/M2/s1 ;
 wire \V3/V1/V1/A3/M3/c1 ;
 wire \V3/V1/V1/A3/M3/c2 ;
 wire \V3/V1/V1/A3/M3/s1 ;
 wire \V3/V1/V1/A3/M4/c1 ;
 wire \V3/V1/V1/A3/M4/c2 ;
 wire \V3/V1/V1/A3/M4/s1 ;
 wire \V3/V1/V1/V1/w1 ;
 wire \V3/V1/V1/V1/w2 ;
 wire \V3/V1/V1/V1/w3 ;
 wire \V3/V1/V1/V1/w4 ;
 wire \V3/V1/V1/V2/w1 ;
 wire \V3/V1/V1/V2/w2 ;
 wire \V3/V1/V1/V2/w3 ;
 wire \V3/V1/V1/V2/w4 ;
 wire \V3/V1/V1/V3/w1 ;
 wire \V3/V1/V1/V3/w2 ;
 wire \V3/V1/V1/V3/w3 ;
 wire \V3/V1/V1/V3/w4 ;
 wire \V3/V1/V1/V4/w1 ;
 wire \V3/V1/V1/V4/w2 ;
 wire \V3/V1/V1/V4/w3 ;
 wire \V3/V1/V1/V4/w4 ;
 wire \V3/V1/V2/c1 ;
 wire \V3/V1/V2/c2 ;
 wire \V3/V1/V2/c3 ;
 wire \V3/V1/V2/overflow ;
 wire \V3/V1/V2/A1/c1 ;
 wire \V3/V1/V2/A1/c2 ;
 wire \V3/V1/V2/A1/c3 ;
 wire \V3/V1/V2/A1/M1/c1 ;
 wire \V3/V1/V2/A1/M1/c2 ;
 wire \V3/V1/V2/A1/M1/s1 ;
 wire \V3/V1/V2/A1/M2/c1 ;
 wire \V3/V1/V2/A1/M2/c2 ;
 wire \V3/V1/V2/A1/M2/s1 ;
 wire \V3/V1/V2/A1/M3/c1 ;
 wire \V3/V1/V2/A1/M3/c2 ;
 wire \V3/V1/V2/A1/M3/s1 ;
 wire \V3/V1/V2/A1/M4/c1 ;
 wire \V3/V1/V2/A1/M4/c2 ;
 wire \V3/V1/V2/A1/M4/s1 ;
 wire \V3/V1/V2/A2/c1 ;
 wire \V3/V1/V2/A2/c2 ;
 wire \V3/V1/V2/A2/c3 ;
 wire \V3/V1/V2/A2/M1/c1 ;
 wire \V3/V1/V2/A2/M1/c2 ;
 wire \V3/V1/V2/A2/M1/s1 ;
 wire \V3/V1/V2/A2/M2/c1 ;
 wire \V3/V1/V2/A2/M2/c2 ;
 wire \V3/V1/V2/A2/M2/s1 ;
 wire \V3/V1/V2/A2/M3/c1 ;
 wire \V3/V1/V2/A2/M3/c2 ;
 wire \V3/V1/V2/A2/M3/s1 ;
 wire \V3/V1/V2/A2/M4/c1 ;
 wire \V3/V1/V2/A2/M4/c2 ;
 wire \V3/V1/V2/A2/M4/s1 ;
 wire \V3/V1/V2/A3/c1 ;
 wire \V3/V1/V2/A3/c2 ;
 wire \V3/V1/V2/A3/c3 ;
 wire \V3/V1/V2/A3/M1/c1 ;
 wire \V3/V1/V2/A3/M1/c2 ;
 wire \V3/V1/V2/A3/M1/s1 ;
 wire \V3/V1/V2/A3/M2/c1 ;
 wire \V3/V1/V2/A3/M2/c2 ;
 wire \V3/V1/V2/A3/M2/s1 ;
 wire \V3/V1/V2/A3/M3/c1 ;
 wire \V3/V1/V2/A3/M3/c2 ;
 wire \V3/V1/V2/A3/M3/s1 ;
 wire \V3/V1/V2/A3/M4/c1 ;
 wire \V3/V1/V2/A3/M4/c2 ;
 wire \V3/V1/V2/A3/M4/s1 ;
 wire \V3/V1/V2/V1/w1 ;
 wire \V3/V1/V2/V1/w2 ;
 wire \V3/V1/V2/V1/w3 ;
 wire \V3/V1/V2/V1/w4 ;
 wire \V3/V1/V2/V2/w1 ;
 wire \V3/V1/V2/V2/w2 ;
 wire \V3/V1/V2/V2/w3 ;
 wire \V3/V1/V2/V2/w4 ;
 wire \V3/V1/V2/V3/w1 ;
 wire \V3/V1/V2/V3/w2 ;
 wire \V3/V1/V2/V3/w3 ;
 wire \V3/V1/V2/V3/w4 ;
 wire \V3/V1/V2/V4/w1 ;
 wire \V3/V1/V2/V4/w2 ;
 wire \V3/V1/V2/V4/w3 ;
 wire \V3/V1/V2/V4/w4 ;
 wire \V3/V1/V3/c1 ;
 wire \V3/V1/V3/c2 ;
 wire \V3/V1/V3/c3 ;
 wire \V3/V1/V3/overflow ;
 wire \V3/V1/V3/A1/c1 ;
 wire \V3/V1/V3/A1/c2 ;
 wire \V3/V1/V3/A1/c3 ;
 wire \V3/V1/V3/A1/M1/c1 ;
 wire \V3/V1/V3/A1/M1/c2 ;
 wire \V3/V1/V3/A1/M1/s1 ;
 wire \V3/V1/V3/A1/M2/c1 ;
 wire \V3/V1/V3/A1/M2/c2 ;
 wire \V3/V1/V3/A1/M2/s1 ;
 wire \V3/V1/V3/A1/M3/c1 ;
 wire \V3/V1/V3/A1/M3/c2 ;
 wire \V3/V1/V3/A1/M3/s1 ;
 wire \V3/V1/V3/A1/M4/c1 ;
 wire \V3/V1/V3/A1/M4/c2 ;
 wire \V3/V1/V3/A1/M4/s1 ;
 wire \V3/V1/V3/A2/c1 ;
 wire \V3/V1/V3/A2/c2 ;
 wire \V3/V1/V3/A2/c3 ;
 wire \V3/V1/V3/A2/M1/c1 ;
 wire \V3/V1/V3/A2/M1/c2 ;
 wire \V3/V1/V3/A2/M1/s1 ;
 wire \V3/V1/V3/A2/M2/c1 ;
 wire \V3/V1/V3/A2/M2/c2 ;
 wire \V3/V1/V3/A2/M2/s1 ;
 wire \V3/V1/V3/A2/M3/c1 ;
 wire \V3/V1/V3/A2/M3/c2 ;
 wire \V3/V1/V3/A2/M3/s1 ;
 wire \V3/V1/V3/A2/M4/c1 ;
 wire \V3/V1/V3/A2/M4/c2 ;
 wire \V3/V1/V3/A2/M4/s1 ;
 wire \V3/V1/V3/A3/c1 ;
 wire \V3/V1/V3/A3/c2 ;
 wire \V3/V1/V3/A3/c3 ;
 wire \V3/V1/V3/A3/M1/c1 ;
 wire \V3/V1/V3/A3/M1/c2 ;
 wire \V3/V1/V3/A3/M1/s1 ;
 wire \V3/V1/V3/A3/M2/c1 ;
 wire \V3/V1/V3/A3/M2/c2 ;
 wire \V3/V1/V3/A3/M2/s1 ;
 wire \V3/V1/V3/A3/M3/c1 ;
 wire \V3/V1/V3/A3/M3/c2 ;
 wire \V3/V1/V3/A3/M3/s1 ;
 wire \V3/V1/V3/A3/M4/c1 ;
 wire \V3/V1/V3/A3/M4/c2 ;
 wire \V3/V1/V3/A3/M4/s1 ;
 wire \V3/V1/V3/V1/w1 ;
 wire \V3/V1/V3/V1/w2 ;
 wire \V3/V1/V3/V1/w3 ;
 wire \V3/V1/V3/V1/w4 ;
 wire \V3/V1/V3/V2/w1 ;
 wire \V3/V1/V3/V2/w2 ;
 wire \V3/V1/V3/V2/w3 ;
 wire \V3/V1/V3/V2/w4 ;
 wire \V3/V1/V3/V3/w1 ;
 wire \V3/V1/V3/V3/w2 ;
 wire \V3/V1/V3/V3/w3 ;
 wire \V3/V1/V3/V3/w4 ;
 wire \V3/V1/V3/V4/w1 ;
 wire \V3/V1/V3/V4/w2 ;
 wire \V3/V1/V3/V4/w3 ;
 wire \V3/V1/V3/V4/w4 ;
 wire \V3/V1/V4/c1 ;
 wire \V3/V1/V4/c2 ;
 wire \V3/V1/V4/c3 ;
 wire \V3/V1/V4/overflow ;
 wire \V3/V1/V4/A1/c1 ;
 wire \V3/V1/V4/A1/c2 ;
 wire \V3/V1/V4/A1/c3 ;
 wire \V3/V1/V4/A1/M1/c1 ;
 wire \V3/V1/V4/A1/M1/c2 ;
 wire \V3/V1/V4/A1/M1/s1 ;
 wire \V3/V1/V4/A1/M2/c1 ;
 wire \V3/V1/V4/A1/M2/c2 ;
 wire \V3/V1/V4/A1/M2/s1 ;
 wire \V3/V1/V4/A1/M3/c1 ;
 wire \V3/V1/V4/A1/M3/c2 ;
 wire \V3/V1/V4/A1/M3/s1 ;
 wire \V3/V1/V4/A1/M4/c1 ;
 wire \V3/V1/V4/A1/M4/c2 ;
 wire \V3/V1/V4/A1/M4/s1 ;
 wire \V3/V1/V4/A2/c1 ;
 wire \V3/V1/V4/A2/c2 ;
 wire \V3/V1/V4/A2/c3 ;
 wire \V3/V1/V4/A2/M1/c1 ;
 wire \V3/V1/V4/A2/M1/c2 ;
 wire \V3/V1/V4/A2/M1/s1 ;
 wire \V3/V1/V4/A2/M2/c1 ;
 wire \V3/V1/V4/A2/M2/c2 ;
 wire \V3/V1/V4/A2/M2/s1 ;
 wire \V3/V1/V4/A2/M3/c1 ;
 wire \V3/V1/V4/A2/M3/c2 ;
 wire \V3/V1/V4/A2/M3/s1 ;
 wire \V3/V1/V4/A2/M4/c1 ;
 wire \V3/V1/V4/A2/M4/c2 ;
 wire \V3/V1/V4/A2/M4/s1 ;
 wire \V3/V1/V4/A3/c1 ;
 wire \V3/V1/V4/A3/c2 ;
 wire \V3/V1/V4/A3/c3 ;
 wire \V3/V1/V4/A3/M1/c1 ;
 wire \V3/V1/V4/A3/M1/c2 ;
 wire \V3/V1/V4/A3/M1/s1 ;
 wire \V3/V1/V4/A3/M2/c1 ;
 wire \V3/V1/V4/A3/M2/c2 ;
 wire \V3/V1/V4/A3/M2/s1 ;
 wire \V3/V1/V4/A3/M3/c1 ;
 wire \V3/V1/V4/A3/M3/c2 ;
 wire \V3/V1/V4/A3/M3/s1 ;
 wire \V3/V1/V4/A3/M4/c1 ;
 wire \V3/V1/V4/A3/M4/c2 ;
 wire \V3/V1/V4/A3/M4/s1 ;
 wire \V3/V1/V4/V1/w1 ;
 wire \V3/V1/V4/V1/w2 ;
 wire \V3/V1/V4/V1/w3 ;
 wire \V3/V1/V4/V1/w4 ;
 wire \V3/V1/V4/V2/w1 ;
 wire \V3/V1/V4/V2/w2 ;
 wire \V3/V1/V4/V2/w3 ;
 wire \V3/V1/V4/V2/w4 ;
 wire \V3/V1/V4/V3/w1 ;
 wire \V3/V1/V4/V3/w2 ;
 wire \V3/V1/V4/V3/w3 ;
 wire \V3/V1/V4/V3/w4 ;
 wire \V3/V1/V4/V4/w1 ;
 wire \V3/V1/V4/V4/w2 ;
 wire \V3/V1/V4/V4/w3 ;
 wire \V3/V1/V4/V4/w4 ;
 wire \V3/V2/c1 ;
 wire \V3/V2/c2 ;
 wire \V3/V2/c3 ;
 wire \V3/V2/overflow ;
 wire \V3/V2/A1/c1 ;
 wire \V3/V2/A1/A1/c1 ;
 wire \V3/V2/A1/A1/c2 ;
 wire \V3/V2/A1/A1/c3 ;
 wire \V3/V2/A1/A1/M1/c1 ;
 wire \V3/V2/A1/A1/M1/c2 ;
 wire \V3/V2/A1/A1/M1/s1 ;
 wire \V3/V2/A1/A1/M2/c1 ;
 wire \V3/V2/A1/A1/M2/c2 ;
 wire \V3/V2/A1/A1/M2/s1 ;
 wire \V3/V2/A1/A1/M3/c1 ;
 wire \V3/V2/A1/A1/M3/c2 ;
 wire \V3/V2/A1/A1/M3/s1 ;
 wire \V3/V2/A1/A1/M4/c1 ;
 wire \V3/V2/A1/A1/M4/c2 ;
 wire \V3/V2/A1/A1/M4/s1 ;
 wire \V3/V2/A1/A2/c1 ;
 wire \V3/V2/A1/A2/c2 ;
 wire \V3/V2/A1/A2/c3 ;
 wire \V3/V2/A1/A2/M1/c1 ;
 wire \V3/V2/A1/A2/M1/c2 ;
 wire \V3/V2/A1/A2/M1/s1 ;
 wire \V3/V2/A1/A2/M2/c1 ;
 wire \V3/V2/A1/A2/M2/c2 ;
 wire \V3/V2/A1/A2/M2/s1 ;
 wire \V3/V2/A1/A2/M3/c1 ;
 wire \V3/V2/A1/A2/M3/c2 ;
 wire \V3/V2/A1/A2/M3/s1 ;
 wire \V3/V2/A1/A2/M4/c1 ;
 wire \V3/V2/A1/A2/M4/c2 ;
 wire \V3/V2/A1/A2/M4/s1 ;
 wire \V3/V2/A2/c1 ;
 wire \V3/V2/A2/A1/c1 ;
 wire \V3/V2/A2/A1/c2 ;
 wire \V3/V2/A2/A1/c3 ;
 wire \V3/V2/A2/A1/M1/c1 ;
 wire \V3/V2/A2/A1/M1/c2 ;
 wire \V3/V2/A2/A1/M1/s1 ;
 wire \V3/V2/A2/A1/M2/c1 ;
 wire \V3/V2/A2/A1/M2/c2 ;
 wire \V3/V2/A2/A1/M2/s1 ;
 wire \V3/V2/A2/A1/M3/c1 ;
 wire \V3/V2/A2/A1/M3/c2 ;
 wire \V3/V2/A2/A1/M3/s1 ;
 wire \V3/V2/A2/A1/M4/c1 ;
 wire \V3/V2/A2/A1/M4/c2 ;
 wire \V3/V2/A2/A1/M4/s1 ;
 wire \V3/V2/A2/A2/c1 ;
 wire \V3/V2/A2/A2/c2 ;
 wire \V3/V2/A2/A2/c3 ;
 wire \V3/V2/A2/A2/M1/c1 ;
 wire \V3/V2/A2/A2/M1/c2 ;
 wire \V3/V2/A2/A2/M1/s1 ;
 wire \V3/V2/A2/A2/M2/c1 ;
 wire \V3/V2/A2/A2/M2/c2 ;
 wire \V3/V2/A2/A2/M2/s1 ;
 wire \V3/V2/A2/A2/M3/c1 ;
 wire \V3/V2/A2/A2/M3/c2 ;
 wire \V3/V2/A2/A2/M3/s1 ;
 wire \V3/V2/A2/A2/M4/c1 ;
 wire \V3/V2/A2/A2/M4/c2 ;
 wire \V3/V2/A2/A2/M4/s1 ;
 wire \V3/V2/A3/c1 ;
 wire \V3/V2/A3/A1/c1 ;
 wire \V3/V2/A3/A1/c2 ;
 wire \V3/V2/A3/A1/c3 ;
 wire \V3/V2/A3/A1/M1/c1 ;
 wire \V3/V2/A3/A1/M1/c2 ;
 wire \V3/V2/A3/A1/M1/s1 ;
 wire \V3/V2/A3/A1/M2/c1 ;
 wire \V3/V2/A3/A1/M2/c2 ;
 wire \V3/V2/A3/A1/M2/s1 ;
 wire \V3/V2/A3/A1/M3/c1 ;
 wire \V3/V2/A3/A1/M3/c2 ;
 wire \V3/V2/A3/A1/M3/s1 ;
 wire \V3/V2/A3/A1/M4/c1 ;
 wire \V3/V2/A3/A1/M4/c2 ;
 wire \V3/V2/A3/A1/M4/s1 ;
 wire \V3/V2/A3/A2/c1 ;
 wire \V3/V2/A3/A2/c2 ;
 wire \V3/V2/A3/A2/c3 ;
 wire \V3/V2/A3/A2/M1/c1 ;
 wire \V3/V2/A3/A2/M1/c2 ;
 wire \V3/V2/A3/A2/M1/s1 ;
 wire \V3/V2/A3/A2/M2/c1 ;
 wire \V3/V2/A3/A2/M2/c2 ;
 wire \V3/V2/A3/A2/M2/s1 ;
 wire \V3/V2/A3/A2/M3/c1 ;
 wire \V3/V2/A3/A2/M3/c2 ;
 wire \V3/V2/A3/A2/M3/s1 ;
 wire \V3/V2/A3/A2/M4/c1 ;
 wire \V3/V2/A3/A2/M4/c2 ;
 wire \V3/V2/A3/A2/M4/s1 ;
 wire \V3/V2/V1/c1 ;
 wire \V3/V2/V1/c2 ;
 wire \V3/V2/V1/c3 ;
 wire \V3/V2/V1/overflow ;
 wire \V3/V2/V1/A1/c1 ;
 wire \V3/V2/V1/A1/c2 ;
 wire \V3/V2/V1/A1/c3 ;
 wire \V3/V2/V1/A1/M1/c1 ;
 wire \V3/V2/V1/A1/M1/c2 ;
 wire \V3/V2/V1/A1/M1/s1 ;
 wire \V3/V2/V1/A1/M2/c1 ;
 wire \V3/V2/V1/A1/M2/c2 ;
 wire \V3/V2/V1/A1/M2/s1 ;
 wire \V3/V2/V1/A1/M3/c1 ;
 wire \V3/V2/V1/A1/M3/c2 ;
 wire \V3/V2/V1/A1/M3/s1 ;
 wire \V3/V2/V1/A1/M4/c1 ;
 wire \V3/V2/V1/A1/M4/c2 ;
 wire \V3/V2/V1/A1/M4/s1 ;
 wire \V3/V2/V1/A2/c1 ;
 wire \V3/V2/V1/A2/c2 ;
 wire \V3/V2/V1/A2/c3 ;
 wire \V3/V2/V1/A2/M1/c1 ;
 wire \V3/V2/V1/A2/M1/c2 ;
 wire \V3/V2/V1/A2/M1/s1 ;
 wire \V3/V2/V1/A2/M2/c1 ;
 wire \V3/V2/V1/A2/M2/c2 ;
 wire \V3/V2/V1/A2/M2/s1 ;
 wire \V3/V2/V1/A2/M3/c1 ;
 wire \V3/V2/V1/A2/M3/c2 ;
 wire \V3/V2/V1/A2/M3/s1 ;
 wire \V3/V2/V1/A2/M4/c1 ;
 wire \V3/V2/V1/A2/M4/c2 ;
 wire \V3/V2/V1/A2/M4/s1 ;
 wire \V3/V2/V1/A3/c1 ;
 wire \V3/V2/V1/A3/c2 ;
 wire \V3/V2/V1/A3/c3 ;
 wire \V3/V2/V1/A3/M1/c1 ;
 wire \V3/V2/V1/A3/M1/c2 ;
 wire \V3/V2/V1/A3/M1/s1 ;
 wire \V3/V2/V1/A3/M2/c1 ;
 wire \V3/V2/V1/A3/M2/c2 ;
 wire \V3/V2/V1/A3/M2/s1 ;
 wire \V3/V2/V1/A3/M3/c1 ;
 wire \V3/V2/V1/A3/M3/c2 ;
 wire \V3/V2/V1/A3/M3/s1 ;
 wire \V3/V2/V1/A3/M4/c1 ;
 wire \V3/V2/V1/A3/M4/c2 ;
 wire \V3/V2/V1/A3/M4/s1 ;
 wire \V3/V2/V1/V1/w1 ;
 wire \V3/V2/V1/V1/w2 ;
 wire \V3/V2/V1/V1/w3 ;
 wire \V3/V2/V1/V1/w4 ;
 wire \V3/V2/V1/V2/w1 ;
 wire \V3/V2/V1/V2/w2 ;
 wire \V3/V2/V1/V2/w3 ;
 wire \V3/V2/V1/V2/w4 ;
 wire \V3/V2/V1/V3/w1 ;
 wire \V3/V2/V1/V3/w2 ;
 wire \V3/V2/V1/V3/w3 ;
 wire \V3/V2/V1/V3/w4 ;
 wire \V3/V2/V1/V4/w1 ;
 wire \V3/V2/V1/V4/w2 ;
 wire \V3/V2/V1/V4/w3 ;
 wire \V3/V2/V1/V4/w4 ;
 wire \V3/V2/V2/c1 ;
 wire \V3/V2/V2/c2 ;
 wire \V3/V2/V2/c3 ;
 wire \V3/V2/V2/overflow ;
 wire \V3/V2/V2/A1/c1 ;
 wire \V3/V2/V2/A1/c2 ;
 wire \V3/V2/V2/A1/c3 ;
 wire \V3/V2/V2/A1/M1/c1 ;
 wire \V3/V2/V2/A1/M1/c2 ;
 wire \V3/V2/V2/A1/M1/s1 ;
 wire \V3/V2/V2/A1/M2/c1 ;
 wire \V3/V2/V2/A1/M2/c2 ;
 wire \V3/V2/V2/A1/M2/s1 ;
 wire \V3/V2/V2/A1/M3/c1 ;
 wire \V3/V2/V2/A1/M3/c2 ;
 wire \V3/V2/V2/A1/M3/s1 ;
 wire \V3/V2/V2/A1/M4/c1 ;
 wire \V3/V2/V2/A1/M4/c2 ;
 wire \V3/V2/V2/A1/M4/s1 ;
 wire \V3/V2/V2/A2/c1 ;
 wire \V3/V2/V2/A2/c2 ;
 wire \V3/V2/V2/A2/c3 ;
 wire \V3/V2/V2/A2/M1/c1 ;
 wire \V3/V2/V2/A2/M1/c2 ;
 wire \V3/V2/V2/A2/M1/s1 ;
 wire \V3/V2/V2/A2/M2/c1 ;
 wire \V3/V2/V2/A2/M2/c2 ;
 wire \V3/V2/V2/A2/M2/s1 ;
 wire \V3/V2/V2/A2/M3/c1 ;
 wire \V3/V2/V2/A2/M3/c2 ;
 wire \V3/V2/V2/A2/M3/s1 ;
 wire \V3/V2/V2/A2/M4/c1 ;
 wire \V3/V2/V2/A2/M4/c2 ;
 wire \V3/V2/V2/A2/M4/s1 ;
 wire \V3/V2/V2/A3/c1 ;
 wire \V3/V2/V2/A3/c2 ;
 wire \V3/V2/V2/A3/c3 ;
 wire \V3/V2/V2/A3/M1/c1 ;
 wire \V3/V2/V2/A3/M1/c2 ;
 wire \V3/V2/V2/A3/M1/s1 ;
 wire \V3/V2/V2/A3/M2/c1 ;
 wire \V3/V2/V2/A3/M2/c2 ;
 wire \V3/V2/V2/A3/M2/s1 ;
 wire \V3/V2/V2/A3/M3/c1 ;
 wire \V3/V2/V2/A3/M3/c2 ;
 wire \V3/V2/V2/A3/M3/s1 ;
 wire \V3/V2/V2/A3/M4/c1 ;
 wire \V3/V2/V2/A3/M4/c2 ;
 wire \V3/V2/V2/A3/M4/s1 ;
 wire \V3/V2/V2/V1/w1 ;
 wire \V3/V2/V2/V1/w2 ;
 wire \V3/V2/V2/V1/w3 ;
 wire \V3/V2/V2/V1/w4 ;
 wire \V3/V2/V2/V2/w1 ;
 wire \V3/V2/V2/V2/w2 ;
 wire \V3/V2/V2/V2/w3 ;
 wire \V3/V2/V2/V2/w4 ;
 wire \V3/V2/V2/V3/w1 ;
 wire \V3/V2/V2/V3/w2 ;
 wire \V3/V2/V2/V3/w3 ;
 wire \V3/V2/V2/V3/w4 ;
 wire \V3/V2/V2/V4/w1 ;
 wire \V3/V2/V2/V4/w2 ;
 wire \V3/V2/V2/V4/w3 ;
 wire \V3/V2/V2/V4/w4 ;
 wire \V3/V2/V3/c1 ;
 wire \V3/V2/V3/c2 ;
 wire \V3/V2/V3/c3 ;
 wire \V3/V2/V3/overflow ;
 wire \V3/V2/V3/A1/c1 ;
 wire \V3/V2/V3/A1/c2 ;
 wire \V3/V2/V3/A1/c3 ;
 wire \V3/V2/V3/A1/M1/c1 ;
 wire \V3/V2/V3/A1/M1/c2 ;
 wire \V3/V2/V3/A1/M1/s1 ;
 wire \V3/V2/V3/A1/M2/c1 ;
 wire \V3/V2/V3/A1/M2/c2 ;
 wire \V3/V2/V3/A1/M2/s1 ;
 wire \V3/V2/V3/A1/M3/c1 ;
 wire \V3/V2/V3/A1/M3/c2 ;
 wire \V3/V2/V3/A1/M3/s1 ;
 wire \V3/V2/V3/A1/M4/c1 ;
 wire \V3/V2/V3/A1/M4/c2 ;
 wire \V3/V2/V3/A1/M4/s1 ;
 wire \V3/V2/V3/A2/c1 ;
 wire \V3/V2/V3/A2/c2 ;
 wire \V3/V2/V3/A2/c3 ;
 wire \V3/V2/V3/A2/M1/c1 ;
 wire \V3/V2/V3/A2/M1/c2 ;
 wire \V3/V2/V3/A2/M1/s1 ;
 wire \V3/V2/V3/A2/M2/c1 ;
 wire \V3/V2/V3/A2/M2/c2 ;
 wire \V3/V2/V3/A2/M2/s1 ;
 wire \V3/V2/V3/A2/M3/c1 ;
 wire \V3/V2/V3/A2/M3/c2 ;
 wire \V3/V2/V3/A2/M3/s1 ;
 wire \V3/V2/V3/A2/M4/c1 ;
 wire \V3/V2/V3/A2/M4/c2 ;
 wire \V3/V2/V3/A2/M4/s1 ;
 wire \V3/V2/V3/A3/c1 ;
 wire \V3/V2/V3/A3/c2 ;
 wire \V3/V2/V3/A3/c3 ;
 wire \V3/V2/V3/A3/M1/c1 ;
 wire \V3/V2/V3/A3/M1/c2 ;
 wire \V3/V2/V3/A3/M1/s1 ;
 wire \V3/V2/V3/A3/M2/c1 ;
 wire \V3/V2/V3/A3/M2/c2 ;
 wire \V3/V2/V3/A3/M2/s1 ;
 wire \V3/V2/V3/A3/M3/c1 ;
 wire \V3/V2/V3/A3/M3/c2 ;
 wire \V3/V2/V3/A3/M3/s1 ;
 wire \V3/V2/V3/A3/M4/c1 ;
 wire \V3/V2/V3/A3/M4/c2 ;
 wire \V3/V2/V3/A3/M4/s1 ;
 wire \V3/V2/V3/V1/w1 ;
 wire \V3/V2/V3/V1/w2 ;
 wire \V3/V2/V3/V1/w3 ;
 wire \V3/V2/V3/V1/w4 ;
 wire \V3/V2/V3/V2/w1 ;
 wire \V3/V2/V3/V2/w2 ;
 wire \V3/V2/V3/V2/w3 ;
 wire \V3/V2/V3/V2/w4 ;
 wire \V3/V2/V3/V3/w1 ;
 wire \V3/V2/V3/V3/w2 ;
 wire \V3/V2/V3/V3/w3 ;
 wire \V3/V2/V3/V3/w4 ;
 wire \V3/V2/V3/V4/w1 ;
 wire \V3/V2/V3/V4/w2 ;
 wire \V3/V2/V3/V4/w3 ;
 wire \V3/V2/V3/V4/w4 ;
 wire \V3/V2/V4/c1 ;
 wire \V3/V2/V4/c2 ;
 wire \V3/V2/V4/c3 ;
 wire \V3/V2/V4/overflow ;
 wire \V3/V2/V4/A1/c1 ;
 wire \V3/V2/V4/A1/c2 ;
 wire \V3/V2/V4/A1/c3 ;
 wire \V3/V2/V4/A1/M1/c1 ;
 wire \V3/V2/V4/A1/M1/c2 ;
 wire \V3/V2/V4/A1/M1/s1 ;
 wire \V3/V2/V4/A1/M2/c1 ;
 wire \V3/V2/V4/A1/M2/c2 ;
 wire \V3/V2/V4/A1/M2/s1 ;
 wire \V3/V2/V4/A1/M3/c1 ;
 wire \V3/V2/V4/A1/M3/c2 ;
 wire \V3/V2/V4/A1/M3/s1 ;
 wire \V3/V2/V4/A1/M4/c1 ;
 wire \V3/V2/V4/A1/M4/c2 ;
 wire \V3/V2/V4/A1/M4/s1 ;
 wire \V3/V2/V4/A2/c1 ;
 wire \V3/V2/V4/A2/c2 ;
 wire \V3/V2/V4/A2/c3 ;
 wire \V3/V2/V4/A2/M1/c1 ;
 wire \V3/V2/V4/A2/M1/c2 ;
 wire \V3/V2/V4/A2/M1/s1 ;
 wire \V3/V2/V4/A2/M2/c1 ;
 wire \V3/V2/V4/A2/M2/c2 ;
 wire \V3/V2/V4/A2/M2/s1 ;
 wire \V3/V2/V4/A2/M3/c1 ;
 wire \V3/V2/V4/A2/M3/c2 ;
 wire \V3/V2/V4/A2/M3/s1 ;
 wire \V3/V2/V4/A2/M4/c1 ;
 wire \V3/V2/V4/A2/M4/c2 ;
 wire \V3/V2/V4/A2/M4/s1 ;
 wire \V3/V2/V4/A3/c1 ;
 wire \V3/V2/V4/A3/c2 ;
 wire \V3/V2/V4/A3/c3 ;
 wire \V3/V2/V4/A3/M1/c1 ;
 wire \V3/V2/V4/A3/M1/c2 ;
 wire \V3/V2/V4/A3/M1/s1 ;
 wire \V3/V2/V4/A3/M2/c1 ;
 wire \V3/V2/V4/A3/M2/c2 ;
 wire \V3/V2/V4/A3/M2/s1 ;
 wire \V3/V2/V4/A3/M3/c1 ;
 wire \V3/V2/V4/A3/M3/c2 ;
 wire \V3/V2/V4/A3/M3/s1 ;
 wire \V3/V2/V4/A3/M4/c1 ;
 wire \V3/V2/V4/A3/M4/c2 ;
 wire \V3/V2/V4/A3/M4/s1 ;
 wire \V3/V2/V4/V1/w1 ;
 wire \V3/V2/V4/V1/w2 ;
 wire \V3/V2/V4/V1/w3 ;
 wire \V3/V2/V4/V1/w4 ;
 wire \V3/V2/V4/V2/w1 ;
 wire \V3/V2/V4/V2/w2 ;
 wire \V3/V2/V4/V2/w3 ;
 wire \V3/V2/V4/V2/w4 ;
 wire \V3/V2/V4/V3/w1 ;
 wire \V3/V2/V4/V3/w2 ;
 wire \V3/V2/V4/V3/w3 ;
 wire \V3/V2/V4/V3/w4 ;
 wire \V3/V2/V4/V4/w1 ;
 wire \V3/V2/V4/V4/w2 ;
 wire \V3/V2/V4/V4/w3 ;
 wire \V3/V2/V4/V4/w4 ;
 wire \V3/V3/c1 ;
 wire \V3/V3/c2 ;
 wire \V3/V3/c3 ;
 wire \V3/V3/overflow ;
 wire \V3/V3/A1/c1 ;
 wire \V3/V3/A1/A1/c1 ;
 wire \V3/V3/A1/A1/c2 ;
 wire \V3/V3/A1/A1/c3 ;
 wire \V3/V3/A1/A1/M1/c1 ;
 wire \V3/V3/A1/A1/M1/c2 ;
 wire \V3/V3/A1/A1/M1/s1 ;
 wire \V3/V3/A1/A1/M2/c1 ;
 wire \V3/V3/A1/A1/M2/c2 ;
 wire \V3/V3/A1/A1/M2/s1 ;
 wire \V3/V3/A1/A1/M3/c1 ;
 wire \V3/V3/A1/A1/M3/c2 ;
 wire \V3/V3/A1/A1/M3/s1 ;
 wire \V3/V3/A1/A1/M4/c1 ;
 wire \V3/V3/A1/A1/M4/c2 ;
 wire \V3/V3/A1/A1/M4/s1 ;
 wire \V3/V3/A1/A2/c1 ;
 wire \V3/V3/A1/A2/c2 ;
 wire \V3/V3/A1/A2/c3 ;
 wire \V3/V3/A1/A2/M1/c1 ;
 wire \V3/V3/A1/A2/M1/c2 ;
 wire \V3/V3/A1/A2/M1/s1 ;
 wire \V3/V3/A1/A2/M2/c1 ;
 wire \V3/V3/A1/A2/M2/c2 ;
 wire \V3/V3/A1/A2/M2/s1 ;
 wire \V3/V3/A1/A2/M3/c1 ;
 wire \V3/V3/A1/A2/M3/c2 ;
 wire \V3/V3/A1/A2/M3/s1 ;
 wire \V3/V3/A1/A2/M4/c1 ;
 wire \V3/V3/A1/A2/M4/c2 ;
 wire \V3/V3/A1/A2/M4/s1 ;
 wire \V3/V3/A2/c1 ;
 wire \V3/V3/A2/A1/c1 ;
 wire \V3/V3/A2/A1/c2 ;
 wire \V3/V3/A2/A1/c3 ;
 wire \V3/V3/A2/A1/M1/c1 ;
 wire \V3/V3/A2/A1/M1/c2 ;
 wire \V3/V3/A2/A1/M1/s1 ;
 wire \V3/V3/A2/A1/M2/c1 ;
 wire \V3/V3/A2/A1/M2/c2 ;
 wire \V3/V3/A2/A1/M2/s1 ;
 wire \V3/V3/A2/A1/M3/c1 ;
 wire \V3/V3/A2/A1/M3/c2 ;
 wire \V3/V3/A2/A1/M3/s1 ;
 wire \V3/V3/A2/A1/M4/c1 ;
 wire \V3/V3/A2/A1/M4/c2 ;
 wire \V3/V3/A2/A1/M4/s1 ;
 wire \V3/V3/A2/A2/c1 ;
 wire \V3/V3/A2/A2/c2 ;
 wire \V3/V3/A2/A2/c3 ;
 wire \V3/V3/A2/A2/M1/c1 ;
 wire \V3/V3/A2/A2/M1/c2 ;
 wire \V3/V3/A2/A2/M1/s1 ;
 wire \V3/V3/A2/A2/M2/c1 ;
 wire \V3/V3/A2/A2/M2/c2 ;
 wire \V3/V3/A2/A2/M2/s1 ;
 wire \V3/V3/A2/A2/M3/c1 ;
 wire \V3/V3/A2/A2/M3/c2 ;
 wire \V3/V3/A2/A2/M3/s1 ;
 wire \V3/V3/A2/A2/M4/c1 ;
 wire \V3/V3/A2/A2/M4/c2 ;
 wire \V3/V3/A2/A2/M4/s1 ;
 wire \V3/V3/A3/c1 ;
 wire \V3/V3/A3/A1/c1 ;
 wire \V3/V3/A3/A1/c2 ;
 wire \V3/V3/A3/A1/c3 ;
 wire \V3/V3/A3/A1/M1/c1 ;
 wire \V3/V3/A3/A1/M1/c2 ;
 wire \V3/V3/A3/A1/M1/s1 ;
 wire \V3/V3/A3/A1/M2/c1 ;
 wire \V3/V3/A3/A1/M2/c2 ;
 wire \V3/V3/A3/A1/M2/s1 ;
 wire \V3/V3/A3/A1/M3/c1 ;
 wire \V3/V3/A3/A1/M3/c2 ;
 wire \V3/V3/A3/A1/M3/s1 ;
 wire \V3/V3/A3/A1/M4/c1 ;
 wire \V3/V3/A3/A1/M4/c2 ;
 wire \V3/V3/A3/A1/M4/s1 ;
 wire \V3/V3/A3/A2/c1 ;
 wire \V3/V3/A3/A2/c2 ;
 wire \V3/V3/A3/A2/c3 ;
 wire \V3/V3/A3/A2/M1/c1 ;
 wire \V3/V3/A3/A2/M1/c2 ;
 wire \V3/V3/A3/A2/M1/s1 ;
 wire \V3/V3/A3/A2/M2/c1 ;
 wire \V3/V3/A3/A2/M2/c2 ;
 wire \V3/V3/A3/A2/M2/s1 ;
 wire \V3/V3/A3/A2/M3/c1 ;
 wire \V3/V3/A3/A2/M3/c2 ;
 wire \V3/V3/A3/A2/M3/s1 ;
 wire \V3/V3/A3/A2/M4/c1 ;
 wire \V3/V3/A3/A2/M4/c2 ;
 wire \V3/V3/A3/A2/M4/s1 ;
 wire \V3/V3/V1/c1 ;
 wire \V3/V3/V1/c2 ;
 wire \V3/V3/V1/c3 ;
 wire \V3/V3/V1/overflow ;
 wire \V3/V3/V1/A1/c1 ;
 wire \V3/V3/V1/A1/c2 ;
 wire \V3/V3/V1/A1/c3 ;
 wire \V3/V3/V1/A1/M1/c1 ;
 wire \V3/V3/V1/A1/M1/c2 ;
 wire \V3/V3/V1/A1/M1/s1 ;
 wire \V3/V3/V1/A1/M2/c1 ;
 wire \V3/V3/V1/A1/M2/c2 ;
 wire \V3/V3/V1/A1/M2/s1 ;
 wire \V3/V3/V1/A1/M3/c1 ;
 wire \V3/V3/V1/A1/M3/c2 ;
 wire \V3/V3/V1/A1/M3/s1 ;
 wire \V3/V3/V1/A1/M4/c1 ;
 wire \V3/V3/V1/A1/M4/c2 ;
 wire \V3/V3/V1/A1/M4/s1 ;
 wire \V3/V3/V1/A2/c1 ;
 wire \V3/V3/V1/A2/c2 ;
 wire \V3/V3/V1/A2/c3 ;
 wire \V3/V3/V1/A2/M1/c1 ;
 wire \V3/V3/V1/A2/M1/c2 ;
 wire \V3/V3/V1/A2/M1/s1 ;
 wire \V3/V3/V1/A2/M2/c1 ;
 wire \V3/V3/V1/A2/M2/c2 ;
 wire \V3/V3/V1/A2/M2/s1 ;
 wire \V3/V3/V1/A2/M3/c1 ;
 wire \V3/V3/V1/A2/M3/c2 ;
 wire \V3/V3/V1/A2/M3/s1 ;
 wire \V3/V3/V1/A2/M4/c1 ;
 wire \V3/V3/V1/A2/M4/c2 ;
 wire \V3/V3/V1/A2/M4/s1 ;
 wire \V3/V3/V1/A3/c1 ;
 wire \V3/V3/V1/A3/c2 ;
 wire \V3/V3/V1/A3/c3 ;
 wire \V3/V3/V1/A3/M1/c1 ;
 wire \V3/V3/V1/A3/M1/c2 ;
 wire \V3/V3/V1/A3/M1/s1 ;
 wire \V3/V3/V1/A3/M2/c1 ;
 wire \V3/V3/V1/A3/M2/c2 ;
 wire \V3/V3/V1/A3/M2/s1 ;
 wire \V3/V3/V1/A3/M3/c1 ;
 wire \V3/V3/V1/A3/M3/c2 ;
 wire \V3/V3/V1/A3/M3/s1 ;
 wire \V3/V3/V1/A3/M4/c1 ;
 wire \V3/V3/V1/A3/M4/c2 ;
 wire \V3/V3/V1/A3/M4/s1 ;
 wire \V3/V3/V1/V1/w1 ;
 wire \V3/V3/V1/V1/w2 ;
 wire \V3/V3/V1/V1/w3 ;
 wire \V3/V3/V1/V1/w4 ;
 wire \V3/V3/V1/V2/w1 ;
 wire \V3/V3/V1/V2/w2 ;
 wire \V3/V3/V1/V2/w3 ;
 wire \V3/V3/V1/V2/w4 ;
 wire \V3/V3/V1/V3/w1 ;
 wire \V3/V3/V1/V3/w2 ;
 wire \V3/V3/V1/V3/w3 ;
 wire \V3/V3/V1/V3/w4 ;
 wire \V3/V3/V1/V4/w1 ;
 wire \V3/V3/V1/V4/w2 ;
 wire \V3/V3/V1/V4/w3 ;
 wire \V3/V3/V1/V4/w4 ;
 wire \V3/V3/V2/c1 ;
 wire \V3/V3/V2/c2 ;
 wire \V3/V3/V2/c3 ;
 wire \V3/V3/V2/overflow ;
 wire \V3/V3/V2/A1/c1 ;
 wire \V3/V3/V2/A1/c2 ;
 wire \V3/V3/V2/A1/c3 ;
 wire \V3/V3/V2/A1/M1/c1 ;
 wire \V3/V3/V2/A1/M1/c2 ;
 wire \V3/V3/V2/A1/M1/s1 ;
 wire \V3/V3/V2/A1/M2/c1 ;
 wire \V3/V3/V2/A1/M2/c2 ;
 wire \V3/V3/V2/A1/M2/s1 ;
 wire \V3/V3/V2/A1/M3/c1 ;
 wire \V3/V3/V2/A1/M3/c2 ;
 wire \V3/V3/V2/A1/M3/s1 ;
 wire \V3/V3/V2/A1/M4/c1 ;
 wire \V3/V3/V2/A1/M4/c2 ;
 wire \V3/V3/V2/A1/M4/s1 ;
 wire \V3/V3/V2/A2/c1 ;
 wire \V3/V3/V2/A2/c2 ;
 wire \V3/V3/V2/A2/c3 ;
 wire \V3/V3/V2/A2/M1/c1 ;
 wire \V3/V3/V2/A2/M1/c2 ;
 wire \V3/V3/V2/A2/M1/s1 ;
 wire \V3/V3/V2/A2/M2/c1 ;
 wire \V3/V3/V2/A2/M2/c2 ;
 wire \V3/V3/V2/A2/M2/s1 ;
 wire \V3/V3/V2/A2/M3/c1 ;
 wire \V3/V3/V2/A2/M3/c2 ;
 wire \V3/V3/V2/A2/M3/s1 ;
 wire \V3/V3/V2/A2/M4/c1 ;
 wire \V3/V3/V2/A2/M4/c2 ;
 wire \V3/V3/V2/A2/M4/s1 ;
 wire \V3/V3/V2/A3/c1 ;
 wire \V3/V3/V2/A3/c2 ;
 wire \V3/V3/V2/A3/c3 ;
 wire \V3/V3/V2/A3/M1/c1 ;
 wire \V3/V3/V2/A3/M1/c2 ;
 wire \V3/V3/V2/A3/M1/s1 ;
 wire \V3/V3/V2/A3/M2/c1 ;
 wire \V3/V3/V2/A3/M2/c2 ;
 wire \V3/V3/V2/A3/M2/s1 ;
 wire \V3/V3/V2/A3/M3/c1 ;
 wire \V3/V3/V2/A3/M3/c2 ;
 wire \V3/V3/V2/A3/M3/s1 ;
 wire \V3/V3/V2/A3/M4/c1 ;
 wire \V3/V3/V2/A3/M4/c2 ;
 wire \V3/V3/V2/A3/M4/s1 ;
 wire \V3/V3/V2/V1/w1 ;
 wire \V3/V3/V2/V1/w2 ;
 wire \V3/V3/V2/V1/w3 ;
 wire \V3/V3/V2/V1/w4 ;
 wire \V3/V3/V2/V2/w1 ;
 wire \V3/V3/V2/V2/w2 ;
 wire \V3/V3/V2/V2/w3 ;
 wire \V3/V3/V2/V2/w4 ;
 wire \V3/V3/V2/V3/w1 ;
 wire \V3/V3/V2/V3/w2 ;
 wire \V3/V3/V2/V3/w3 ;
 wire \V3/V3/V2/V3/w4 ;
 wire \V3/V3/V2/V4/w1 ;
 wire \V3/V3/V2/V4/w2 ;
 wire \V3/V3/V2/V4/w3 ;
 wire \V3/V3/V2/V4/w4 ;
 wire \V3/V3/V3/c1 ;
 wire \V3/V3/V3/c2 ;
 wire \V3/V3/V3/c3 ;
 wire \V3/V3/V3/overflow ;
 wire \V3/V3/V3/A1/c1 ;
 wire \V3/V3/V3/A1/c2 ;
 wire \V3/V3/V3/A1/c3 ;
 wire \V3/V3/V3/A1/M1/c1 ;
 wire \V3/V3/V3/A1/M1/c2 ;
 wire \V3/V3/V3/A1/M1/s1 ;
 wire \V3/V3/V3/A1/M2/c1 ;
 wire \V3/V3/V3/A1/M2/c2 ;
 wire \V3/V3/V3/A1/M2/s1 ;
 wire \V3/V3/V3/A1/M3/c1 ;
 wire \V3/V3/V3/A1/M3/c2 ;
 wire \V3/V3/V3/A1/M3/s1 ;
 wire \V3/V3/V3/A1/M4/c1 ;
 wire \V3/V3/V3/A1/M4/c2 ;
 wire \V3/V3/V3/A1/M4/s1 ;
 wire \V3/V3/V3/A2/c1 ;
 wire \V3/V3/V3/A2/c2 ;
 wire \V3/V3/V3/A2/c3 ;
 wire \V3/V3/V3/A2/M1/c1 ;
 wire \V3/V3/V3/A2/M1/c2 ;
 wire \V3/V3/V3/A2/M1/s1 ;
 wire \V3/V3/V3/A2/M2/c1 ;
 wire \V3/V3/V3/A2/M2/c2 ;
 wire \V3/V3/V3/A2/M2/s1 ;
 wire \V3/V3/V3/A2/M3/c1 ;
 wire \V3/V3/V3/A2/M3/c2 ;
 wire \V3/V3/V3/A2/M3/s1 ;
 wire \V3/V3/V3/A2/M4/c1 ;
 wire \V3/V3/V3/A2/M4/c2 ;
 wire \V3/V3/V3/A2/M4/s1 ;
 wire \V3/V3/V3/A3/c1 ;
 wire \V3/V3/V3/A3/c2 ;
 wire \V3/V3/V3/A3/c3 ;
 wire \V3/V3/V3/A3/M1/c1 ;
 wire \V3/V3/V3/A3/M1/c2 ;
 wire \V3/V3/V3/A3/M1/s1 ;
 wire \V3/V3/V3/A3/M2/c1 ;
 wire \V3/V3/V3/A3/M2/c2 ;
 wire \V3/V3/V3/A3/M2/s1 ;
 wire \V3/V3/V3/A3/M3/c1 ;
 wire \V3/V3/V3/A3/M3/c2 ;
 wire \V3/V3/V3/A3/M3/s1 ;
 wire \V3/V3/V3/A3/M4/c1 ;
 wire \V3/V3/V3/A3/M4/c2 ;
 wire \V3/V3/V3/A3/M4/s1 ;
 wire \V3/V3/V3/V1/w1 ;
 wire \V3/V3/V3/V1/w2 ;
 wire \V3/V3/V3/V1/w3 ;
 wire \V3/V3/V3/V1/w4 ;
 wire \V3/V3/V3/V2/w1 ;
 wire \V3/V3/V3/V2/w2 ;
 wire \V3/V3/V3/V2/w3 ;
 wire \V3/V3/V3/V2/w4 ;
 wire \V3/V3/V3/V3/w1 ;
 wire \V3/V3/V3/V3/w2 ;
 wire \V3/V3/V3/V3/w3 ;
 wire \V3/V3/V3/V3/w4 ;
 wire \V3/V3/V3/V4/w1 ;
 wire \V3/V3/V3/V4/w2 ;
 wire \V3/V3/V3/V4/w3 ;
 wire \V3/V3/V3/V4/w4 ;
 wire \V3/V3/V4/c1 ;
 wire \V3/V3/V4/c2 ;
 wire \V3/V3/V4/c3 ;
 wire \V3/V3/V4/overflow ;
 wire \V3/V3/V4/A1/c1 ;
 wire \V3/V3/V4/A1/c2 ;
 wire \V3/V3/V4/A1/c3 ;
 wire \V3/V3/V4/A1/M1/c1 ;
 wire \V3/V3/V4/A1/M1/c2 ;
 wire \V3/V3/V4/A1/M1/s1 ;
 wire \V3/V3/V4/A1/M2/c1 ;
 wire \V3/V3/V4/A1/M2/c2 ;
 wire \V3/V3/V4/A1/M2/s1 ;
 wire \V3/V3/V4/A1/M3/c1 ;
 wire \V3/V3/V4/A1/M3/c2 ;
 wire \V3/V3/V4/A1/M3/s1 ;
 wire \V3/V3/V4/A1/M4/c1 ;
 wire \V3/V3/V4/A1/M4/c2 ;
 wire \V3/V3/V4/A1/M4/s1 ;
 wire \V3/V3/V4/A2/c1 ;
 wire \V3/V3/V4/A2/c2 ;
 wire \V3/V3/V4/A2/c3 ;
 wire \V3/V3/V4/A2/M1/c1 ;
 wire \V3/V3/V4/A2/M1/c2 ;
 wire \V3/V3/V4/A2/M1/s1 ;
 wire \V3/V3/V4/A2/M2/c1 ;
 wire \V3/V3/V4/A2/M2/c2 ;
 wire \V3/V3/V4/A2/M2/s1 ;
 wire \V3/V3/V4/A2/M3/c1 ;
 wire \V3/V3/V4/A2/M3/c2 ;
 wire \V3/V3/V4/A2/M3/s1 ;
 wire \V3/V3/V4/A2/M4/c1 ;
 wire \V3/V3/V4/A2/M4/c2 ;
 wire \V3/V3/V4/A2/M4/s1 ;
 wire \V3/V3/V4/A3/c1 ;
 wire \V3/V3/V4/A3/c2 ;
 wire \V3/V3/V4/A3/c3 ;
 wire \V3/V3/V4/A3/M1/c1 ;
 wire \V3/V3/V4/A3/M1/c2 ;
 wire \V3/V3/V4/A3/M1/s1 ;
 wire \V3/V3/V4/A3/M2/c1 ;
 wire \V3/V3/V4/A3/M2/c2 ;
 wire \V3/V3/V4/A3/M2/s1 ;
 wire \V3/V3/V4/A3/M3/c1 ;
 wire \V3/V3/V4/A3/M3/c2 ;
 wire \V3/V3/V4/A3/M3/s1 ;
 wire \V3/V3/V4/A3/M4/c1 ;
 wire \V3/V3/V4/A3/M4/c2 ;
 wire \V3/V3/V4/A3/M4/s1 ;
 wire \V3/V3/V4/V1/w1 ;
 wire \V3/V3/V4/V1/w2 ;
 wire \V3/V3/V4/V1/w3 ;
 wire \V3/V3/V4/V1/w4 ;
 wire \V3/V3/V4/V2/w1 ;
 wire \V3/V3/V4/V2/w2 ;
 wire \V3/V3/V4/V2/w3 ;
 wire \V3/V3/V4/V2/w4 ;
 wire \V3/V3/V4/V3/w1 ;
 wire \V3/V3/V4/V3/w2 ;
 wire \V3/V3/V4/V3/w3 ;
 wire \V3/V3/V4/V3/w4 ;
 wire \V3/V3/V4/V4/w1 ;
 wire \V3/V3/V4/V4/w2 ;
 wire \V3/V3/V4/V4/w3 ;
 wire \V3/V3/V4/V4/w4 ;
 wire \V3/V4/c1 ;
 wire \V3/V4/c2 ;
 wire \V3/V4/c3 ;
 wire \V3/V4/overflow ;
 wire \V3/V4/A1/c1 ;
 wire \V3/V4/A1/A1/c1 ;
 wire \V3/V4/A1/A1/c2 ;
 wire \V3/V4/A1/A1/c3 ;
 wire \V3/V4/A1/A1/M1/c1 ;
 wire \V3/V4/A1/A1/M1/c2 ;
 wire \V3/V4/A1/A1/M1/s1 ;
 wire \V3/V4/A1/A1/M2/c1 ;
 wire \V3/V4/A1/A1/M2/c2 ;
 wire \V3/V4/A1/A1/M2/s1 ;
 wire \V3/V4/A1/A1/M3/c1 ;
 wire \V3/V4/A1/A1/M3/c2 ;
 wire \V3/V4/A1/A1/M3/s1 ;
 wire \V3/V4/A1/A1/M4/c1 ;
 wire \V3/V4/A1/A1/M4/c2 ;
 wire \V3/V4/A1/A1/M4/s1 ;
 wire \V3/V4/A1/A2/c1 ;
 wire \V3/V4/A1/A2/c2 ;
 wire \V3/V4/A1/A2/c3 ;
 wire \V3/V4/A1/A2/M1/c1 ;
 wire \V3/V4/A1/A2/M1/c2 ;
 wire \V3/V4/A1/A2/M1/s1 ;
 wire \V3/V4/A1/A2/M2/c1 ;
 wire \V3/V4/A1/A2/M2/c2 ;
 wire \V3/V4/A1/A2/M2/s1 ;
 wire \V3/V4/A1/A2/M3/c1 ;
 wire \V3/V4/A1/A2/M3/c2 ;
 wire \V3/V4/A1/A2/M3/s1 ;
 wire \V3/V4/A1/A2/M4/c1 ;
 wire \V3/V4/A1/A2/M4/c2 ;
 wire \V3/V4/A1/A2/M4/s1 ;
 wire \V3/V4/A2/c1 ;
 wire \V3/V4/A2/A1/c1 ;
 wire \V3/V4/A2/A1/c2 ;
 wire \V3/V4/A2/A1/c3 ;
 wire \V3/V4/A2/A1/M1/c1 ;
 wire \V3/V4/A2/A1/M1/c2 ;
 wire \V3/V4/A2/A1/M1/s1 ;
 wire \V3/V4/A2/A1/M2/c1 ;
 wire \V3/V4/A2/A1/M2/c2 ;
 wire \V3/V4/A2/A1/M2/s1 ;
 wire \V3/V4/A2/A1/M3/c1 ;
 wire \V3/V4/A2/A1/M3/c2 ;
 wire \V3/V4/A2/A1/M3/s1 ;
 wire \V3/V4/A2/A1/M4/c1 ;
 wire \V3/V4/A2/A1/M4/c2 ;
 wire \V3/V4/A2/A1/M4/s1 ;
 wire \V3/V4/A2/A2/c1 ;
 wire \V3/V4/A2/A2/c2 ;
 wire \V3/V4/A2/A2/c3 ;
 wire \V3/V4/A2/A2/M1/c1 ;
 wire \V3/V4/A2/A2/M1/c2 ;
 wire \V3/V4/A2/A2/M1/s1 ;
 wire \V3/V4/A2/A2/M2/c1 ;
 wire \V3/V4/A2/A2/M2/c2 ;
 wire \V3/V4/A2/A2/M2/s1 ;
 wire \V3/V4/A2/A2/M3/c1 ;
 wire \V3/V4/A2/A2/M3/c2 ;
 wire \V3/V4/A2/A2/M3/s1 ;
 wire \V3/V4/A2/A2/M4/c1 ;
 wire \V3/V4/A2/A2/M4/c2 ;
 wire \V3/V4/A2/A2/M4/s1 ;
 wire \V3/V4/A3/c1 ;
 wire \V3/V4/A3/A1/c1 ;
 wire \V3/V4/A3/A1/c2 ;
 wire \V3/V4/A3/A1/c3 ;
 wire \V3/V4/A3/A1/M1/c1 ;
 wire \V3/V4/A3/A1/M1/c2 ;
 wire \V3/V4/A3/A1/M1/s1 ;
 wire \V3/V4/A3/A1/M2/c1 ;
 wire \V3/V4/A3/A1/M2/c2 ;
 wire \V3/V4/A3/A1/M2/s1 ;
 wire \V3/V4/A3/A1/M3/c1 ;
 wire \V3/V4/A3/A1/M3/c2 ;
 wire \V3/V4/A3/A1/M3/s1 ;
 wire \V3/V4/A3/A1/M4/c1 ;
 wire \V3/V4/A3/A1/M4/c2 ;
 wire \V3/V4/A3/A1/M4/s1 ;
 wire \V3/V4/A3/A2/c1 ;
 wire \V3/V4/A3/A2/c2 ;
 wire \V3/V4/A3/A2/c3 ;
 wire \V3/V4/A3/A2/M1/c1 ;
 wire \V3/V4/A3/A2/M1/c2 ;
 wire \V3/V4/A3/A2/M1/s1 ;
 wire \V3/V4/A3/A2/M2/c1 ;
 wire \V3/V4/A3/A2/M2/c2 ;
 wire \V3/V4/A3/A2/M2/s1 ;
 wire \V3/V4/A3/A2/M3/c1 ;
 wire \V3/V4/A3/A2/M3/c2 ;
 wire \V3/V4/A3/A2/M3/s1 ;
 wire \V3/V4/A3/A2/M4/c1 ;
 wire \V3/V4/A3/A2/M4/c2 ;
 wire \V3/V4/A3/A2/M4/s1 ;
 wire \V3/V4/V1/c1 ;
 wire \V3/V4/V1/c2 ;
 wire \V3/V4/V1/c3 ;
 wire \V3/V4/V1/overflow ;
 wire \V3/V4/V1/A1/c1 ;
 wire \V3/V4/V1/A1/c2 ;
 wire \V3/V4/V1/A1/c3 ;
 wire \V3/V4/V1/A1/M1/c1 ;
 wire \V3/V4/V1/A1/M1/c2 ;
 wire \V3/V4/V1/A1/M1/s1 ;
 wire \V3/V4/V1/A1/M2/c1 ;
 wire \V3/V4/V1/A1/M2/c2 ;
 wire \V3/V4/V1/A1/M2/s1 ;
 wire \V3/V4/V1/A1/M3/c1 ;
 wire \V3/V4/V1/A1/M3/c2 ;
 wire \V3/V4/V1/A1/M3/s1 ;
 wire \V3/V4/V1/A1/M4/c1 ;
 wire \V3/V4/V1/A1/M4/c2 ;
 wire \V3/V4/V1/A1/M4/s1 ;
 wire \V3/V4/V1/A2/c1 ;
 wire \V3/V4/V1/A2/c2 ;
 wire \V3/V4/V1/A2/c3 ;
 wire \V3/V4/V1/A2/M1/c1 ;
 wire \V3/V4/V1/A2/M1/c2 ;
 wire \V3/V4/V1/A2/M1/s1 ;
 wire \V3/V4/V1/A2/M2/c1 ;
 wire \V3/V4/V1/A2/M2/c2 ;
 wire \V3/V4/V1/A2/M2/s1 ;
 wire \V3/V4/V1/A2/M3/c1 ;
 wire \V3/V4/V1/A2/M3/c2 ;
 wire \V3/V4/V1/A2/M3/s1 ;
 wire \V3/V4/V1/A2/M4/c1 ;
 wire \V3/V4/V1/A2/M4/c2 ;
 wire \V3/V4/V1/A2/M4/s1 ;
 wire \V3/V4/V1/A3/c1 ;
 wire \V3/V4/V1/A3/c2 ;
 wire \V3/V4/V1/A3/c3 ;
 wire \V3/V4/V1/A3/M1/c1 ;
 wire \V3/V4/V1/A3/M1/c2 ;
 wire \V3/V4/V1/A3/M1/s1 ;
 wire \V3/V4/V1/A3/M2/c1 ;
 wire \V3/V4/V1/A3/M2/c2 ;
 wire \V3/V4/V1/A3/M2/s1 ;
 wire \V3/V4/V1/A3/M3/c1 ;
 wire \V3/V4/V1/A3/M3/c2 ;
 wire \V3/V4/V1/A3/M3/s1 ;
 wire \V3/V4/V1/A3/M4/c1 ;
 wire \V3/V4/V1/A3/M4/c2 ;
 wire \V3/V4/V1/A3/M4/s1 ;
 wire \V3/V4/V1/V1/w1 ;
 wire \V3/V4/V1/V1/w2 ;
 wire \V3/V4/V1/V1/w3 ;
 wire \V3/V4/V1/V1/w4 ;
 wire \V3/V4/V1/V2/w1 ;
 wire \V3/V4/V1/V2/w2 ;
 wire \V3/V4/V1/V2/w3 ;
 wire \V3/V4/V1/V2/w4 ;
 wire \V3/V4/V1/V3/w1 ;
 wire \V3/V4/V1/V3/w2 ;
 wire \V3/V4/V1/V3/w3 ;
 wire \V3/V4/V1/V3/w4 ;
 wire \V3/V4/V1/V4/w1 ;
 wire \V3/V4/V1/V4/w2 ;
 wire \V3/V4/V1/V4/w3 ;
 wire \V3/V4/V1/V4/w4 ;
 wire \V3/V4/V2/c1 ;
 wire \V3/V4/V2/c2 ;
 wire \V3/V4/V2/c3 ;
 wire \V3/V4/V2/overflow ;
 wire \V3/V4/V2/A1/c1 ;
 wire \V3/V4/V2/A1/c2 ;
 wire \V3/V4/V2/A1/c3 ;
 wire \V3/V4/V2/A1/M1/c1 ;
 wire \V3/V4/V2/A1/M1/c2 ;
 wire \V3/V4/V2/A1/M1/s1 ;
 wire \V3/V4/V2/A1/M2/c1 ;
 wire \V3/V4/V2/A1/M2/c2 ;
 wire \V3/V4/V2/A1/M2/s1 ;
 wire \V3/V4/V2/A1/M3/c1 ;
 wire \V3/V4/V2/A1/M3/c2 ;
 wire \V3/V4/V2/A1/M3/s1 ;
 wire \V3/V4/V2/A1/M4/c1 ;
 wire \V3/V4/V2/A1/M4/c2 ;
 wire \V3/V4/V2/A1/M4/s1 ;
 wire \V3/V4/V2/A2/c1 ;
 wire \V3/V4/V2/A2/c2 ;
 wire \V3/V4/V2/A2/c3 ;
 wire \V3/V4/V2/A2/M1/c1 ;
 wire \V3/V4/V2/A2/M1/c2 ;
 wire \V3/V4/V2/A2/M1/s1 ;
 wire \V3/V4/V2/A2/M2/c1 ;
 wire \V3/V4/V2/A2/M2/c2 ;
 wire \V3/V4/V2/A2/M2/s1 ;
 wire \V3/V4/V2/A2/M3/c1 ;
 wire \V3/V4/V2/A2/M3/c2 ;
 wire \V3/V4/V2/A2/M3/s1 ;
 wire \V3/V4/V2/A2/M4/c1 ;
 wire \V3/V4/V2/A2/M4/c2 ;
 wire \V3/V4/V2/A2/M4/s1 ;
 wire \V3/V4/V2/A3/c1 ;
 wire \V3/V4/V2/A3/c2 ;
 wire \V3/V4/V2/A3/c3 ;
 wire \V3/V4/V2/A3/M1/c1 ;
 wire \V3/V4/V2/A3/M1/c2 ;
 wire \V3/V4/V2/A3/M1/s1 ;
 wire \V3/V4/V2/A3/M2/c1 ;
 wire \V3/V4/V2/A3/M2/c2 ;
 wire \V3/V4/V2/A3/M2/s1 ;
 wire \V3/V4/V2/A3/M3/c1 ;
 wire \V3/V4/V2/A3/M3/c2 ;
 wire \V3/V4/V2/A3/M3/s1 ;
 wire \V3/V4/V2/A3/M4/c1 ;
 wire \V3/V4/V2/A3/M4/c2 ;
 wire \V3/V4/V2/A3/M4/s1 ;
 wire \V3/V4/V2/V1/w1 ;
 wire \V3/V4/V2/V1/w2 ;
 wire \V3/V4/V2/V1/w3 ;
 wire \V3/V4/V2/V1/w4 ;
 wire \V3/V4/V2/V2/w1 ;
 wire \V3/V4/V2/V2/w2 ;
 wire \V3/V4/V2/V2/w3 ;
 wire \V3/V4/V2/V2/w4 ;
 wire \V3/V4/V2/V3/w1 ;
 wire \V3/V4/V2/V3/w2 ;
 wire \V3/V4/V2/V3/w3 ;
 wire \V3/V4/V2/V3/w4 ;
 wire \V3/V4/V2/V4/w1 ;
 wire \V3/V4/V2/V4/w2 ;
 wire \V3/V4/V2/V4/w3 ;
 wire \V3/V4/V2/V4/w4 ;
 wire \V3/V4/V3/c1 ;
 wire \V3/V4/V3/c2 ;
 wire \V3/V4/V3/c3 ;
 wire \V3/V4/V3/overflow ;
 wire \V3/V4/V3/A1/c1 ;
 wire \V3/V4/V3/A1/c2 ;
 wire \V3/V4/V3/A1/c3 ;
 wire \V3/V4/V3/A1/M1/c1 ;
 wire \V3/V4/V3/A1/M1/c2 ;
 wire \V3/V4/V3/A1/M1/s1 ;
 wire \V3/V4/V3/A1/M2/c1 ;
 wire \V3/V4/V3/A1/M2/c2 ;
 wire \V3/V4/V3/A1/M2/s1 ;
 wire \V3/V4/V3/A1/M3/c1 ;
 wire \V3/V4/V3/A1/M3/c2 ;
 wire \V3/V4/V3/A1/M3/s1 ;
 wire \V3/V4/V3/A1/M4/c1 ;
 wire \V3/V4/V3/A1/M4/c2 ;
 wire \V3/V4/V3/A1/M4/s1 ;
 wire \V3/V4/V3/A2/c1 ;
 wire \V3/V4/V3/A2/c2 ;
 wire \V3/V4/V3/A2/c3 ;
 wire \V3/V4/V3/A2/M1/c1 ;
 wire \V3/V4/V3/A2/M1/c2 ;
 wire \V3/V4/V3/A2/M1/s1 ;
 wire \V3/V4/V3/A2/M2/c1 ;
 wire \V3/V4/V3/A2/M2/c2 ;
 wire \V3/V4/V3/A2/M2/s1 ;
 wire \V3/V4/V3/A2/M3/c1 ;
 wire \V3/V4/V3/A2/M3/c2 ;
 wire \V3/V4/V3/A2/M3/s1 ;
 wire \V3/V4/V3/A2/M4/c1 ;
 wire \V3/V4/V3/A2/M4/c2 ;
 wire \V3/V4/V3/A2/M4/s1 ;
 wire \V3/V4/V3/A3/c1 ;
 wire \V3/V4/V3/A3/c2 ;
 wire \V3/V4/V3/A3/c3 ;
 wire \V3/V4/V3/A3/M1/c1 ;
 wire \V3/V4/V3/A3/M1/c2 ;
 wire \V3/V4/V3/A3/M1/s1 ;
 wire \V3/V4/V3/A3/M2/c1 ;
 wire \V3/V4/V3/A3/M2/c2 ;
 wire \V3/V4/V3/A3/M2/s1 ;
 wire \V3/V4/V3/A3/M3/c1 ;
 wire \V3/V4/V3/A3/M3/c2 ;
 wire \V3/V4/V3/A3/M3/s1 ;
 wire \V3/V4/V3/A3/M4/c1 ;
 wire \V3/V4/V3/A3/M4/c2 ;
 wire \V3/V4/V3/A3/M4/s1 ;
 wire \V3/V4/V3/V1/w1 ;
 wire \V3/V4/V3/V1/w2 ;
 wire \V3/V4/V3/V1/w3 ;
 wire \V3/V4/V3/V1/w4 ;
 wire \V3/V4/V3/V2/w1 ;
 wire \V3/V4/V3/V2/w2 ;
 wire \V3/V4/V3/V2/w3 ;
 wire \V3/V4/V3/V2/w4 ;
 wire \V3/V4/V3/V3/w1 ;
 wire \V3/V4/V3/V3/w2 ;
 wire \V3/V4/V3/V3/w3 ;
 wire \V3/V4/V3/V3/w4 ;
 wire \V3/V4/V3/V4/w1 ;
 wire \V3/V4/V3/V4/w2 ;
 wire \V3/V4/V3/V4/w3 ;
 wire \V3/V4/V3/V4/w4 ;
 wire \V3/V4/V4/c1 ;
 wire \V3/V4/V4/c2 ;
 wire \V3/V4/V4/c3 ;
 wire \V3/V4/V4/overflow ;
 wire \V3/V4/V4/A1/c1 ;
 wire \V3/V4/V4/A1/c2 ;
 wire \V3/V4/V4/A1/c3 ;
 wire \V3/V4/V4/A1/M1/c1 ;
 wire \V3/V4/V4/A1/M1/c2 ;
 wire \V3/V4/V4/A1/M1/s1 ;
 wire \V3/V4/V4/A1/M2/c1 ;
 wire \V3/V4/V4/A1/M2/c2 ;
 wire \V3/V4/V4/A1/M2/s1 ;
 wire \V3/V4/V4/A1/M3/c1 ;
 wire \V3/V4/V4/A1/M3/c2 ;
 wire \V3/V4/V4/A1/M3/s1 ;
 wire \V3/V4/V4/A1/M4/c1 ;
 wire \V3/V4/V4/A1/M4/c2 ;
 wire \V3/V4/V4/A1/M4/s1 ;
 wire \V3/V4/V4/A2/c1 ;
 wire \V3/V4/V4/A2/c2 ;
 wire \V3/V4/V4/A2/c3 ;
 wire \V3/V4/V4/A2/M1/c1 ;
 wire \V3/V4/V4/A2/M1/c2 ;
 wire \V3/V4/V4/A2/M1/s1 ;
 wire \V3/V4/V4/A2/M2/c1 ;
 wire \V3/V4/V4/A2/M2/c2 ;
 wire \V3/V4/V4/A2/M2/s1 ;
 wire \V3/V4/V4/A2/M3/c1 ;
 wire \V3/V4/V4/A2/M3/c2 ;
 wire \V3/V4/V4/A2/M3/s1 ;
 wire \V3/V4/V4/A2/M4/c1 ;
 wire \V3/V4/V4/A2/M4/c2 ;
 wire \V3/V4/V4/A2/M4/s1 ;
 wire \V3/V4/V4/A3/c1 ;
 wire \V3/V4/V4/A3/c2 ;
 wire \V3/V4/V4/A3/c3 ;
 wire \V3/V4/V4/A3/M1/c1 ;
 wire \V3/V4/V4/A3/M1/c2 ;
 wire \V3/V4/V4/A3/M1/s1 ;
 wire \V3/V4/V4/A3/M2/c1 ;
 wire \V3/V4/V4/A3/M2/c2 ;
 wire \V3/V4/V4/A3/M2/s1 ;
 wire \V3/V4/V4/A3/M3/c1 ;
 wire \V3/V4/V4/A3/M3/c2 ;
 wire \V3/V4/V4/A3/M3/s1 ;
 wire \V3/V4/V4/A3/M4/c1 ;
 wire \V3/V4/V4/A3/M4/c2 ;
 wire \V3/V4/V4/A3/M4/s1 ;
 wire \V3/V4/V4/V1/w1 ;
 wire \V3/V4/V4/V1/w2 ;
 wire \V3/V4/V4/V1/w3 ;
 wire \V3/V4/V4/V1/w4 ;
 wire \V3/V4/V4/V2/w1 ;
 wire \V3/V4/V4/V2/w2 ;
 wire \V3/V4/V4/V2/w3 ;
 wire \V3/V4/V4/V2/w4 ;
 wire \V3/V4/V4/V3/w1 ;
 wire \V3/V4/V4/V3/w2 ;
 wire \V3/V4/V4/V3/w3 ;
 wire \V3/V4/V4/V3/w4 ;
 wire \V3/V4/V4/V4/w1 ;
 wire \V3/V4/V4/V4/w2 ;
 wire \V3/V4/V4/V4/w3 ;
 wire \V3/V4/V4/V4/w4 ;
 wire \V4/c1 ;
 wire \V4/c2 ;
 wire \V4/c3 ;
 wire \V4/overflow ;
 wire \V4/A1/c1 ;
 wire \V4/A1/A1/c1 ;
 wire \V4/A1/A1/A1/c1 ;
 wire \V4/A1/A1/A1/c2 ;
 wire \V4/A1/A1/A1/c3 ;
 wire \V4/A1/A1/A1/M1/c1 ;
 wire \V4/A1/A1/A1/M1/c2 ;
 wire \V4/A1/A1/A1/M1/s1 ;
 wire \V4/A1/A1/A1/M2/c1 ;
 wire \V4/A1/A1/A1/M2/c2 ;
 wire \V4/A1/A1/A1/M2/s1 ;
 wire \V4/A1/A1/A1/M3/c1 ;
 wire \V4/A1/A1/A1/M3/c2 ;
 wire \V4/A1/A1/A1/M3/s1 ;
 wire \V4/A1/A1/A1/M4/c1 ;
 wire \V4/A1/A1/A1/M4/c2 ;
 wire \V4/A1/A1/A1/M4/s1 ;
 wire \V4/A1/A1/A2/c1 ;
 wire \V4/A1/A1/A2/c2 ;
 wire \V4/A1/A1/A2/c3 ;
 wire \V4/A1/A1/A2/M1/c1 ;
 wire \V4/A1/A1/A2/M1/c2 ;
 wire \V4/A1/A1/A2/M1/s1 ;
 wire \V4/A1/A1/A2/M2/c1 ;
 wire \V4/A1/A1/A2/M2/c2 ;
 wire \V4/A1/A1/A2/M2/s1 ;
 wire \V4/A1/A1/A2/M3/c1 ;
 wire \V4/A1/A1/A2/M3/c2 ;
 wire \V4/A1/A1/A2/M3/s1 ;
 wire \V4/A1/A1/A2/M4/c1 ;
 wire \V4/A1/A1/A2/M4/c2 ;
 wire \V4/A1/A1/A2/M4/s1 ;
 wire \V4/A1/A2/c1 ;
 wire \V4/A1/A2/A1/c1 ;
 wire \V4/A1/A2/A1/c2 ;
 wire \V4/A1/A2/A1/c3 ;
 wire \V4/A1/A2/A1/M1/c1 ;
 wire \V4/A1/A2/A1/M1/c2 ;
 wire \V4/A1/A2/A1/M1/s1 ;
 wire \V4/A1/A2/A1/M2/c1 ;
 wire \V4/A1/A2/A1/M2/c2 ;
 wire \V4/A1/A2/A1/M2/s1 ;
 wire \V4/A1/A2/A1/M3/c1 ;
 wire \V4/A1/A2/A1/M3/c2 ;
 wire \V4/A1/A2/A1/M3/s1 ;
 wire \V4/A1/A2/A1/M4/c1 ;
 wire \V4/A1/A2/A1/M4/c2 ;
 wire \V4/A1/A2/A1/M4/s1 ;
 wire \V4/A1/A2/A2/c1 ;
 wire \V4/A1/A2/A2/c2 ;
 wire \V4/A1/A2/A2/c3 ;
 wire \V4/A1/A2/A2/M1/c1 ;
 wire \V4/A1/A2/A2/M1/c2 ;
 wire \V4/A1/A2/A2/M1/s1 ;
 wire \V4/A1/A2/A2/M2/c1 ;
 wire \V4/A1/A2/A2/M2/c2 ;
 wire \V4/A1/A2/A2/M2/s1 ;
 wire \V4/A1/A2/A2/M3/c1 ;
 wire \V4/A1/A2/A2/M3/c2 ;
 wire \V4/A1/A2/A2/M3/s1 ;
 wire \V4/A1/A2/A2/M4/c1 ;
 wire \V4/A1/A2/A2/M4/c2 ;
 wire \V4/A1/A2/A2/M4/s1 ;
 wire \V4/A2/c1 ;
 wire \V4/A2/A1/c1 ;
 wire \V4/A2/A1/A1/c1 ;
 wire \V4/A2/A1/A1/c2 ;
 wire \V4/A2/A1/A1/c3 ;
 wire \V4/A2/A1/A1/M1/c1 ;
 wire \V4/A2/A1/A1/M1/c2 ;
 wire \V4/A2/A1/A1/M1/s1 ;
 wire \V4/A2/A1/A1/M2/c1 ;
 wire \V4/A2/A1/A1/M2/c2 ;
 wire \V4/A2/A1/A1/M2/s1 ;
 wire \V4/A2/A1/A1/M3/c1 ;
 wire \V4/A2/A1/A1/M3/c2 ;
 wire \V4/A2/A1/A1/M3/s1 ;
 wire \V4/A2/A1/A1/M4/c1 ;
 wire \V4/A2/A1/A1/M4/c2 ;
 wire \V4/A2/A1/A1/M4/s1 ;
 wire \V4/A2/A1/A2/c1 ;
 wire \V4/A2/A1/A2/c2 ;
 wire \V4/A2/A1/A2/c3 ;
 wire \V4/A2/A1/A2/M1/c1 ;
 wire \V4/A2/A1/A2/M1/c2 ;
 wire \V4/A2/A1/A2/M1/s1 ;
 wire \V4/A2/A1/A2/M2/c1 ;
 wire \V4/A2/A1/A2/M2/c2 ;
 wire \V4/A2/A1/A2/M2/s1 ;
 wire \V4/A2/A1/A2/M3/c1 ;
 wire \V4/A2/A1/A2/M3/c2 ;
 wire \V4/A2/A1/A2/M3/s1 ;
 wire \V4/A2/A1/A2/M4/c1 ;
 wire \V4/A2/A1/A2/M4/c2 ;
 wire \V4/A2/A1/A2/M4/s1 ;
 wire \V4/A2/A2/c1 ;
 wire \V4/A2/A2/A1/c1 ;
 wire \V4/A2/A2/A1/c2 ;
 wire \V4/A2/A2/A1/c3 ;
 wire \V4/A2/A2/A1/M1/c1 ;
 wire \V4/A2/A2/A1/M1/c2 ;
 wire \V4/A2/A2/A1/M1/s1 ;
 wire \V4/A2/A2/A1/M2/c1 ;
 wire \V4/A2/A2/A1/M2/c2 ;
 wire \V4/A2/A2/A1/M2/s1 ;
 wire \V4/A2/A2/A1/M3/c1 ;
 wire \V4/A2/A2/A1/M3/c2 ;
 wire \V4/A2/A2/A1/M3/s1 ;
 wire \V4/A2/A2/A1/M4/c1 ;
 wire \V4/A2/A2/A1/M4/c2 ;
 wire \V4/A2/A2/A1/M4/s1 ;
 wire \V4/A2/A2/A2/c1 ;
 wire \V4/A2/A2/A2/c2 ;
 wire \V4/A2/A2/A2/c3 ;
 wire \V4/A2/A2/A2/M1/c1 ;
 wire \V4/A2/A2/A2/M1/c2 ;
 wire \V4/A2/A2/A2/M1/s1 ;
 wire \V4/A2/A2/A2/M2/c1 ;
 wire \V4/A2/A2/A2/M2/c2 ;
 wire \V4/A2/A2/A2/M2/s1 ;
 wire \V4/A2/A2/A2/M3/c1 ;
 wire \V4/A2/A2/A2/M3/c2 ;
 wire \V4/A2/A2/A2/M3/s1 ;
 wire \V4/A2/A2/A2/M4/c1 ;
 wire \V4/A2/A2/A2/M4/c2 ;
 wire \V4/A2/A2/A2/M4/s1 ;
 wire \V4/A3/c1 ;
 wire \V4/A3/A1/c1 ;
 wire \V4/A3/A1/A1/c1 ;
 wire \V4/A3/A1/A1/c2 ;
 wire \V4/A3/A1/A1/c3 ;
 wire \V4/A3/A1/A1/M1/c1 ;
 wire \V4/A3/A1/A1/M1/c2 ;
 wire \V4/A3/A1/A1/M1/s1 ;
 wire \V4/A3/A1/A1/M2/c1 ;
 wire \V4/A3/A1/A1/M2/c2 ;
 wire \V4/A3/A1/A1/M2/s1 ;
 wire \V4/A3/A1/A1/M3/c1 ;
 wire \V4/A3/A1/A1/M3/c2 ;
 wire \V4/A3/A1/A1/M3/s1 ;
 wire \V4/A3/A1/A1/M4/c1 ;
 wire \V4/A3/A1/A1/M4/c2 ;
 wire \V4/A3/A1/A1/M4/s1 ;
 wire \V4/A3/A1/A2/c1 ;
 wire \V4/A3/A1/A2/c2 ;
 wire \V4/A3/A1/A2/c3 ;
 wire \V4/A3/A1/A2/M1/c1 ;
 wire \V4/A3/A1/A2/M1/c2 ;
 wire \V4/A3/A1/A2/M1/s1 ;
 wire \V4/A3/A1/A2/M2/c1 ;
 wire \V4/A3/A1/A2/M2/c2 ;
 wire \V4/A3/A1/A2/M2/s1 ;
 wire \V4/A3/A1/A2/M3/c1 ;
 wire \V4/A3/A1/A2/M3/c2 ;
 wire \V4/A3/A1/A2/M3/s1 ;
 wire \V4/A3/A1/A2/M4/c1 ;
 wire \V4/A3/A1/A2/M4/c2 ;
 wire \V4/A3/A1/A2/M4/s1 ;
 wire \V4/A3/A2/c1 ;
 wire \V4/A3/A2/A1/c1 ;
 wire \V4/A3/A2/A1/c2 ;
 wire \V4/A3/A2/A1/c3 ;
 wire \V4/A3/A2/A1/M1/c1 ;
 wire \V4/A3/A2/A1/M1/c2 ;
 wire \V4/A3/A2/A1/M1/s1 ;
 wire \V4/A3/A2/A1/M2/c1 ;
 wire \V4/A3/A2/A1/M2/c2 ;
 wire \V4/A3/A2/A1/M2/s1 ;
 wire \V4/A3/A2/A1/M3/c1 ;
 wire \V4/A3/A2/A1/M3/c2 ;
 wire \V4/A3/A2/A1/M3/s1 ;
 wire \V4/A3/A2/A1/M4/c1 ;
 wire \V4/A3/A2/A1/M4/c2 ;
 wire \V4/A3/A2/A1/M4/s1 ;
 wire \V4/A3/A2/A2/c1 ;
 wire \V4/A3/A2/A2/c2 ;
 wire \V4/A3/A2/A2/c3 ;
 wire \V4/A3/A2/A2/M1/c1 ;
 wire \V4/A3/A2/A2/M1/c2 ;
 wire \V4/A3/A2/A2/M1/s1 ;
 wire \V4/A3/A2/A2/M2/c1 ;
 wire \V4/A3/A2/A2/M2/c2 ;
 wire \V4/A3/A2/A2/M2/s1 ;
 wire \V4/A3/A2/A2/M3/c1 ;
 wire \V4/A3/A2/A2/M3/c2 ;
 wire \V4/A3/A2/A2/M3/s1 ;
 wire \V4/A3/A2/A2/M4/c1 ;
 wire \V4/A3/A2/A2/M4/c2 ;
 wire \V4/A3/A2/A2/M4/s1 ;
 wire \V4/V1/c1 ;
 wire \V4/V1/c2 ;
 wire \V4/V1/c3 ;
 wire \V4/V1/overflow ;
 wire \V4/V1/A1/c1 ;
 wire \V4/V1/A1/A1/c1 ;
 wire \V4/V1/A1/A1/c2 ;
 wire \V4/V1/A1/A1/c3 ;
 wire \V4/V1/A1/A1/M1/c1 ;
 wire \V4/V1/A1/A1/M1/c2 ;
 wire \V4/V1/A1/A1/M1/s1 ;
 wire \V4/V1/A1/A1/M2/c1 ;
 wire \V4/V1/A1/A1/M2/c2 ;
 wire \V4/V1/A1/A1/M2/s1 ;
 wire \V4/V1/A1/A1/M3/c1 ;
 wire \V4/V1/A1/A1/M3/c2 ;
 wire \V4/V1/A1/A1/M3/s1 ;
 wire \V4/V1/A1/A1/M4/c1 ;
 wire \V4/V1/A1/A1/M4/c2 ;
 wire \V4/V1/A1/A1/M4/s1 ;
 wire \V4/V1/A1/A2/c1 ;
 wire \V4/V1/A1/A2/c2 ;
 wire \V4/V1/A1/A2/c3 ;
 wire \V4/V1/A1/A2/M1/c1 ;
 wire \V4/V1/A1/A2/M1/c2 ;
 wire \V4/V1/A1/A2/M1/s1 ;
 wire \V4/V1/A1/A2/M2/c1 ;
 wire \V4/V1/A1/A2/M2/c2 ;
 wire \V4/V1/A1/A2/M2/s1 ;
 wire \V4/V1/A1/A2/M3/c1 ;
 wire \V4/V1/A1/A2/M3/c2 ;
 wire \V4/V1/A1/A2/M3/s1 ;
 wire \V4/V1/A1/A2/M4/c1 ;
 wire \V4/V1/A1/A2/M4/c2 ;
 wire \V4/V1/A1/A2/M4/s1 ;
 wire \V4/V1/A2/c1 ;
 wire \V4/V1/A2/A1/c1 ;
 wire \V4/V1/A2/A1/c2 ;
 wire \V4/V1/A2/A1/c3 ;
 wire \V4/V1/A2/A1/M1/c1 ;
 wire \V4/V1/A2/A1/M1/c2 ;
 wire \V4/V1/A2/A1/M1/s1 ;
 wire \V4/V1/A2/A1/M2/c1 ;
 wire \V4/V1/A2/A1/M2/c2 ;
 wire \V4/V1/A2/A1/M2/s1 ;
 wire \V4/V1/A2/A1/M3/c1 ;
 wire \V4/V1/A2/A1/M3/c2 ;
 wire \V4/V1/A2/A1/M3/s1 ;
 wire \V4/V1/A2/A1/M4/c1 ;
 wire \V4/V1/A2/A1/M4/c2 ;
 wire \V4/V1/A2/A1/M4/s1 ;
 wire \V4/V1/A2/A2/c1 ;
 wire \V4/V1/A2/A2/c2 ;
 wire \V4/V1/A2/A2/c3 ;
 wire \V4/V1/A2/A2/M1/c1 ;
 wire \V4/V1/A2/A2/M1/c2 ;
 wire \V4/V1/A2/A2/M1/s1 ;
 wire \V4/V1/A2/A2/M2/c1 ;
 wire \V4/V1/A2/A2/M2/c2 ;
 wire \V4/V1/A2/A2/M2/s1 ;
 wire \V4/V1/A2/A2/M3/c1 ;
 wire \V4/V1/A2/A2/M3/c2 ;
 wire \V4/V1/A2/A2/M3/s1 ;
 wire \V4/V1/A2/A2/M4/c1 ;
 wire \V4/V1/A2/A2/M4/c2 ;
 wire \V4/V1/A2/A2/M4/s1 ;
 wire \V4/V1/A3/c1 ;
 wire \V4/V1/A3/A1/c1 ;
 wire \V4/V1/A3/A1/c2 ;
 wire \V4/V1/A3/A1/c3 ;
 wire \V4/V1/A3/A1/M1/c1 ;
 wire \V4/V1/A3/A1/M1/c2 ;
 wire \V4/V1/A3/A1/M1/s1 ;
 wire \V4/V1/A3/A1/M2/c1 ;
 wire \V4/V1/A3/A1/M2/c2 ;
 wire \V4/V1/A3/A1/M2/s1 ;
 wire \V4/V1/A3/A1/M3/c1 ;
 wire \V4/V1/A3/A1/M3/c2 ;
 wire \V4/V1/A3/A1/M3/s1 ;
 wire \V4/V1/A3/A1/M4/c1 ;
 wire \V4/V1/A3/A1/M4/c2 ;
 wire \V4/V1/A3/A1/M4/s1 ;
 wire \V4/V1/A3/A2/c1 ;
 wire \V4/V1/A3/A2/c2 ;
 wire \V4/V1/A3/A2/c3 ;
 wire \V4/V1/A3/A2/M1/c1 ;
 wire \V4/V1/A3/A2/M1/c2 ;
 wire \V4/V1/A3/A2/M1/s1 ;
 wire \V4/V1/A3/A2/M2/c1 ;
 wire \V4/V1/A3/A2/M2/c2 ;
 wire \V4/V1/A3/A2/M2/s1 ;
 wire \V4/V1/A3/A2/M3/c1 ;
 wire \V4/V1/A3/A2/M3/c2 ;
 wire \V4/V1/A3/A2/M3/s1 ;
 wire \V4/V1/A3/A2/M4/c1 ;
 wire \V4/V1/A3/A2/M4/c2 ;
 wire \V4/V1/A3/A2/M4/s1 ;
 wire \V4/V1/V1/c1 ;
 wire \V4/V1/V1/c2 ;
 wire \V4/V1/V1/c3 ;
 wire \V4/V1/V1/overflow ;
 wire \V4/V1/V1/A1/c1 ;
 wire \V4/V1/V1/A1/c2 ;
 wire \V4/V1/V1/A1/c3 ;
 wire \V4/V1/V1/A1/M1/c1 ;
 wire \V4/V1/V1/A1/M1/c2 ;
 wire \V4/V1/V1/A1/M1/s1 ;
 wire \V4/V1/V1/A1/M2/c1 ;
 wire \V4/V1/V1/A1/M2/c2 ;
 wire \V4/V1/V1/A1/M2/s1 ;
 wire \V4/V1/V1/A1/M3/c1 ;
 wire \V4/V1/V1/A1/M3/c2 ;
 wire \V4/V1/V1/A1/M3/s1 ;
 wire \V4/V1/V1/A1/M4/c1 ;
 wire \V4/V1/V1/A1/M4/c2 ;
 wire \V4/V1/V1/A1/M4/s1 ;
 wire \V4/V1/V1/A2/c1 ;
 wire \V4/V1/V1/A2/c2 ;
 wire \V4/V1/V1/A2/c3 ;
 wire \V4/V1/V1/A2/M1/c1 ;
 wire \V4/V1/V1/A2/M1/c2 ;
 wire \V4/V1/V1/A2/M1/s1 ;
 wire \V4/V1/V1/A2/M2/c1 ;
 wire \V4/V1/V1/A2/M2/c2 ;
 wire \V4/V1/V1/A2/M2/s1 ;
 wire \V4/V1/V1/A2/M3/c1 ;
 wire \V4/V1/V1/A2/M3/c2 ;
 wire \V4/V1/V1/A2/M3/s1 ;
 wire \V4/V1/V1/A2/M4/c1 ;
 wire \V4/V1/V1/A2/M4/c2 ;
 wire \V4/V1/V1/A2/M4/s1 ;
 wire \V4/V1/V1/A3/c1 ;
 wire \V4/V1/V1/A3/c2 ;
 wire \V4/V1/V1/A3/c3 ;
 wire \V4/V1/V1/A3/M1/c1 ;
 wire \V4/V1/V1/A3/M1/c2 ;
 wire \V4/V1/V1/A3/M1/s1 ;
 wire \V4/V1/V1/A3/M2/c1 ;
 wire \V4/V1/V1/A3/M2/c2 ;
 wire \V4/V1/V1/A3/M2/s1 ;
 wire \V4/V1/V1/A3/M3/c1 ;
 wire \V4/V1/V1/A3/M3/c2 ;
 wire \V4/V1/V1/A3/M3/s1 ;
 wire \V4/V1/V1/A3/M4/c1 ;
 wire \V4/V1/V1/A3/M4/c2 ;
 wire \V4/V1/V1/A3/M4/s1 ;
 wire \V4/V1/V1/V1/w1 ;
 wire \V4/V1/V1/V1/w2 ;
 wire \V4/V1/V1/V1/w3 ;
 wire \V4/V1/V1/V1/w4 ;
 wire \V4/V1/V1/V2/w1 ;
 wire \V4/V1/V1/V2/w2 ;
 wire \V4/V1/V1/V2/w3 ;
 wire \V4/V1/V1/V2/w4 ;
 wire \V4/V1/V1/V3/w1 ;
 wire \V4/V1/V1/V3/w2 ;
 wire \V4/V1/V1/V3/w3 ;
 wire \V4/V1/V1/V3/w4 ;
 wire \V4/V1/V1/V4/w1 ;
 wire \V4/V1/V1/V4/w2 ;
 wire \V4/V1/V1/V4/w3 ;
 wire \V4/V1/V1/V4/w4 ;
 wire \V4/V1/V2/c1 ;
 wire \V4/V1/V2/c2 ;
 wire \V4/V1/V2/c3 ;
 wire \V4/V1/V2/overflow ;
 wire \V4/V1/V2/A1/c1 ;
 wire \V4/V1/V2/A1/c2 ;
 wire \V4/V1/V2/A1/c3 ;
 wire \V4/V1/V2/A1/M1/c1 ;
 wire \V4/V1/V2/A1/M1/c2 ;
 wire \V4/V1/V2/A1/M1/s1 ;
 wire \V4/V1/V2/A1/M2/c1 ;
 wire \V4/V1/V2/A1/M2/c2 ;
 wire \V4/V1/V2/A1/M2/s1 ;
 wire \V4/V1/V2/A1/M3/c1 ;
 wire \V4/V1/V2/A1/M3/c2 ;
 wire \V4/V1/V2/A1/M3/s1 ;
 wire \V4/V1/V2/A1/M4/c1 ;
 wire \V4/V1/V2/A1/M4/c2 ;
 wire \V4/V1/V2/A1/M4/s1 ;
 wire \V4/V1/V2/A2/c1 ;
 wire \V4/V1/V2/A2/c2 ;
 wire \V4/V1/V2/A2/c3 ;
 wire \V4/V1/V2/A2/M1/c1 ;
 wire \V4/V1/V2/A2/M1/c2 ;
 wire \V4/V1/V2/A2/M1/s1 ;
 wire \V4/V1/V2/A2/M2/c1 ;
 wire \V4/V1/V2/A2/M2/c2 ;
 wire \V4/V1/V2/A2/M2/s1 ;
 wire \V4/V1/V2/A2/M3/c1 ;
 wire \V4/V1/V2/A2/M3/c2 ;
 wire \V4/V1/V2/A2/M3/s1 ;
 wire \V4/V1/V2/A2/M4/c1 ;
 wire \V4/V1/V2/A2/M4/c2 ;
 wire \V4/V1/V2/A2/M4/s1 ;
 wire \V4/V1/V2/A3/c1 ;
 wire \V4/V1/V2/A3/c2 ;
 wire \V4/V1/V2/A3/c3 ;
 wire \V4/V1/V2/A3/M1/c1 ;
 wire \V4/V1/V2/A3/M1/c2 ;
 wire \V4/V1/V2/A3/M1/s1 ;
 wire \V4/V1/V2/A3/M2/c1 ;
 wire \V4/V1/V2/A3/M2/c2 ;
 wire \V4/V1/V2/A3/M2/s1 ;
 wire \V4/V1/V2/A3/M3/c1 ;
 wire \V4/V1/V2/A3/M3/c2 ;
 wire \V4/V1/V2/A3/M3/s1 ;
 wire \V4/V1/V2/A3/M4/c1 ;
 wire \V4/V1/V2/A3/M4/c2 ;
 wire \V4/V1/V2/A3/M4/s1 ;
 wire \V4/V1/V2/V1/w1 ;
 wire \V4/V1/V2/V1/w2 ;
 wire \V4/V1/V2/V1/w3 ;
 wire \V4/V1/V2/V1/w4 ;
 wire \V4/V1/V2/V2/w1 ;
 wire \V4/V1/V2/V2/w2 ;
 wire \V4/V1/V2/V2/w3 ;
 wire \V4/V1/V2/V2/w4 ;
 wire \V4/V1/V2/V3/w1 ;
 wire \V4/V1/V2/V3/w2 ;
 wire \V4/V1/V2/V3/w3 ;
 wire \V4/V1/V2/V3/w4 ;
 wire \V4/V1/V2/V4/w1 ;
 wire \V4/V1/V2/V4/w2 ;
 wire \V4/V1/V2/V4/w3 ;
 wire \V4/V1/V2/V4/w4 ;
 wire \V4/V1/V3/c1 ;
 wire \V4/V1/V3/c2 ;
 wire \V4/V1/V3/c3 ;
 wire \V4/V1/V3/overflow ;
 wire \V4/V1/V3/A1/c1 ;
 wire \V4/V1/V3/A1/c2 ;
 wire \V4/V1/V3/A1/c3 ;
 wire \V4/V1/V3/A1/M1/c1 ;
 wire \V4/V1/V3/A1/M1/c2 ;
 wire \V4/V1/V3/A1/M1/s1 ;
 wire \V4/V1/V3/A1/M2/c1 ;
 wire \V4/V1/V3/A1/M2/c2 ;
 wire \V4/V1/V3/A1/M2/s1 ;
 wire \V4/V1/V3/A1/M3/c1 ;
 wire \V4/V1/V3/A1/M3/c2 ;
 wire \V4/V1/V3/A1/M3/s1 ;
 wire \V4/V1/V3/A1/M4/c1 ;
 wire \V4/V1/V3/A1/M4/c2 ;
 wire \V4/V1/V3/A1/M4/s1 ;
 wire \V4/V1/V3/A2/c1 ;
 wire \V4/V1/V3/A2/c2 ;
 wire \V4/V1/V3/A2/c3 ;
 wire \V4/V1/V3/A2/M1/c1 ;
 wire \V4/V1/V3/A2/M1/c2 ;
 wire \V4/V1/V3/A2/M1/s1 ;
 wire \V4/V1/V3/A2/M2/c1 ;
 wire \V4/V1/V3/A2/M2/c2 ;
 wire \V4/V1/V3/A2/M2/s1 ;
 wire \V4/V1/V3/A2/M3/c1 ;
 wire \V4/V1/V3/A2/M3/c2 ;
 wire \V4/V1/V3/A2/M3/s1 ;
 wire \V4/V1/V3/A2/M4/c1 ;
 wire \V4/V1/V3/A2/M4/c2 ;
 wire \V4/V1/V3/A2/M4/s1 ;
 wire \V4/V1/V3/A3/c1 ;
 wire \V4/V1/V3/A3/c2 ;
 wire \V4/V1/V3/A3/c3 ;
 wire \V4/V1/V3/A3/M1/c1 ;
 wire \V4/V1/V3/A3/M1/c2 ;
 wire \V4/V1/V3/A3/M1/s1 ;
 wire \V4/V1/V3/A3/M2/c1 ;
 wire \V4/V1/V3/A3/M2/c2 ;
 wire \V4/V1/V3/A3/M2/s1 ;
 wire \V4/V1/V3/A3/M3/c1 ;
 wire \V4/V1/V3/A3/M3/c2 ;
 wire \V4/V1/V3/A3/M3/s1 ;
 wire \V4/V1/V3/A3/M4/c1 ;
 wire \V4/V1/V3/A3/M4/c2 ;
 wire \V4/V1/V3/A3/M4/s1 ;
 wire \V4/V1/V3/V1/w1 ;
 wire \V4/V1/V3/V1/w2 ;
 wire \V4/V1/V3/V1/w3 ;
 wire \V4/V1/V3/V1/w4 ;
 wire \V4/V1/V3/V2/w1 ;
 wire \V4/V1/V3/V2/w2 ;
 wire \V4/V1/V3/V2/w3 ;
 wire \V4/V1/V3/V2/w4 ;
 wire \V4/V1/V3/V3/w1 ;
 wire \V4/V1/V3/V3/w2 ;
 wire \V4/V1/V3/V3/w3 ;
 wire \V4/V1/V3/V3/w4 ;
 wire \V4/V1/V3/V4/w1 ;
 wire \V4/V1/V3/V4/w2 ;
 wire \V4/V1/V3/V4/w3 ;
 wire \V4/V1/V3/V4/w4 ;
 wire \V4/V1/V4/c1 ;
 wire \V4/V1/V4/c2 ;
 wire \V4/V1/V4/c3 ;
 wire \V4/V1/V4/overflow ;
 wire \V4/V1/V4/A1/c1 ;
 wire \V4/V1/V4/A1/c2 ;
 wire \V4/V1/V4/A1/c3 ;
 wire \V4/V1/V4/A1/M1/c1 ;
 wire \V4/V1/V4/A1/M1/c2 ;
 wire \V4/V1/V4/A1/M1/s1 ;
 wire \V4/V1/V4/A1/M2/c1 ;
 wire \V4/V1/V4/A1/M2/c2 ;
 wire \V4/V1/V4/A1/M2/s1 ;
 wire \V4/V1/V4/A1/M3/c1 ;
 wire \V4/V1/V4/A1/M3/c2 ;
 wire \V4/V1/V4/A1/M3/s1 ;
 wire \V4/V1/V4/A1/M4/c1 ;
 wire \V4/V1/V4/A1/M4/c2 ;
 wire \V4/V1/V4/A1/M4/s1 ;
 wire \V4/V1/V4/A2/c1 ;
 wire \V4/V1/V4/A2/c2 ;
 wire \V4/V1/V4/A2/c3 ;
 wire \V4/V1/V4/A2/M1/c1 ;
 wire \V4/V1/V4/A2/M1/c2 ;
 wire \V4/V1/V4/A2/M1/s1 ;
 wire \V4/V1/V4/A2/M2/c1 ;
 wire \V4/V1/V4/A2/M2/c2 ;
 wire \V4/V1/V4/A2/M2/s1 ;
 wire \V4/V1/V4/A2/M3/c1 ;
 wire \V4/V1/V4/A2/M3/c2 ;
 wire \V4/V1/V4/A2/M3/s1 ;
 wire \V4/V1/V4/A2/M4/c1 ;
 wire \V4/V1/V4/A2/M4/c2 ;
 wire \V4/V1/V4/A2/M4/s1 ;
 wire \V4/V1/V4/A3/c1 ;
 wire \V4/V1/V4/A3/c2 ;
 wire \V4/V1/V4/A3/c3 ;
 wire \V4/V1/V4/A3/M1/c1 ;
 wire \V4/V1/V4/A3/M1/c2 ;
 wire \V4/V1/V4/A3/M1/s1 ;
 wire \V4/V1/V4/A3/M2/c1 ;
 wire \V4/V1/V4/A3/M2/c2 ;
 wire \V4/V1/V4/A3/M2/s1 ;
 wire \V4/V1/V4/A3/M3/c1 ;
 wire \V4/V1/V4/A3/M3/c2 ;
 wire \V4/V1/V4/A3/M3/s1 ;
 wire \V4/V1/V4/A3/M4/c1 ;
 wire \V4/V1/V4/A3/M4/c2 ;
 wire \V4/V1/V4/A3/M4/s1 ;
 wire \V4/V1/V4/V1/w1 ;
 wire \V4/V1/V4/V1/w2 ;
 wire \V4/V1/V4/V1/w3 ;
 wire \V4/V1/V4/V1/w4 ;
 wire \V4/V1/V4/V2/w1 ;
 wire \V4/V1/V4/V2/w2 ;
 wire \V4/V1/V4/V2/w3 ;
 wire \V4/V1/V4/V2/w4 ;
 wire \V4/V1/V4/V3/w1 ;
 wire \V4/V1/V4/V3/w2 ;
 wire \V4/V1/V4/V3/w3 ;
 wire \V4/V1/V4/V3/w4 ;
 wire \V4/V1/V4/V4/w1 ;
 wire \V4/V1/V4/V4/w2 ;
 wire \V4/V1/V4/V4/w3 ;
 wire \V4/V1/V4/V4/w4 ;
 wire \V4/V2/c1 ;
 wire \V4/V2/c2 ;
 wire \V4/V2/c3 ;
 wire \V4/V2/overflow ;
 wire \V4/V2/A1/c1 ;
 wire \V4/V2/A1/A1/c1 ;
 wire \V4/V2/A1/A1/c2 ;
 wire \V4/V2/A1/A1/c3 ;
 wire \V4/V2/A1/A1/M1/c1 ;
 wire \V4/V2/A1/A1/M1/c2 ;
 wire \V4/V2/A1/A1/M1/s1 ;
 wire \V4/V2/A1/A1/M2/c1 ;
 wire \V4/V2/A1/A1/M2/c2 ;
 wire \V4/V2/A1/A1/M2/s1 ;
 wire \V4/V2/A1/A1/M3/c1 ;
 wire \V4/V2/A1/A1/M3/c2 ;
 wire \V4/V2/A1/A1/M3/s1 ;
 wire \V4/V2/A1/A1/M4/c1 ;
 wire \V4/V2/A1/A1/M4/c2 ;
 wire \V4/V2/A1/A1/M4/s1 ;
 wire \V4/V2/A1/A2/c1 ;
 wire \V4/V2/A1/A2/c2 ;
 wire \V4/V2/A1/A2/c3 ;
 wire \V4/V2/A1/A2/M1/c1 ;
 wire \V4/V2/A1/A2/M1/c2 ;
 wire \V4/V2/A1/A2/M1/s1 ;
 wire \V4/V2/A1/A2/M2/c1 ;
 wire \V4/V2/A1/A2/M2/c2 ;
 wire \V4/V2/A1/A2/M2/s1 ;
 wire \V4/V2/A1/A2/M3/c1 ;
 wire \V4/V2/A1/A2/M3/c2 ;
 wire \V4/V2/A1/A2/M3/s1 ;
 wire \V4/V2/A1/A2/M4/c1 ;
 wire \V4/V2/A1/A2/M4/c2 ;
 wire \V4/V2/A1/A2/M4/s1 ;
 wire \V4/V2/A2/c1 ;
 wire \V4/V2/A2/A1/c1 ;
 wire \V4/V2/A2/A1/c2 ;
 wire \V4/V2/A2/A1/c3 ;
 wire \V4/V2/A2/A1/M1/c1 ;
 wire \V4/V2/A2/A1/M1/c2 ;
 wire \V4/V2/A2/A1/M1/s1 ;
 wire \V4/V2/A2/A1/M2/c1 ;
 wire \V4/V2/A2/A1/M2/c2 ;
 wire \V4/V2/A2/A1/M2/s1 ;
 wire \V4/V2/A2/A1/M3/c1 ;
 wire \V4/V2/A2/A1/M3/c2 ;
 wire \V4/V2/A2/A1/M3/s1 ;
 wire \V4/V2/A2/A1/M4/c1 ;
 wire \V4/V2/A2/A1/M4/c2 ;
 wire \V4/V2/A2/A1/M4/s1 ;
 wire \V4/V2/A2/A2/c1 ;
 wire \V4/V2/A2/A2/c2 ;
 wire \V4/V2/A2/A2/c3 ;
 wire \V4/V2/A2/A2/M1/c1 ;
 wire \V4/V2/A2/A2/M1/c2 ;
 wire \V4/V2/A2/A2/M1/s1 ;
 wire \V4/V2/A2/A2/M2/c1 ;
 wire \V4/V2/A2/A2/M2/c2 ;
 wire \V4/V2/A2/A2/M2/s1 ;
 wire \V4/V2/A2/A2/M3/c1 ;
 wire \V4/V2/A2/A2/M3/c2 ;
 wire \V4/V2/A2/A2/M3/s1 ;
 wire \V4/V2/A2/A2/M4/c1 ;
 wire \V4/V2/A2/A2/M4/c2 ;
 wire \V4/V2/A2/A2/M4/s1 ;
 wire \V4/V2/A3/c1 ;
 wire \V4/V2/A3/A1/c1 ;
 wire \V4/V2/A3/A1/c2 ;
 wire \V4/V2/A3/A1/c3 ;
 wire \V4/V2/A3/A1/M1/c1 ;
 wire \V4/V2/A3/A1/M1/c2 ;
 wire \V4/V2/A3/A1/M1/s1 ;
 wire \V4/V2/A3/A1/M2/c1 ;
 wire \V4/V2/A3/A1/M2/c2 ;
 wire \V4/V2/A3/A1/M2/s1 ;
 wire \V4/V2/A3/A1/M3/c1 ;
 wire \V4/V2/A3/A1/M3/c2 ;
 wire \V4/V2/A3/A1/M3/s1 ;
 wire \V4/V2/A3/A1/M4/c1 ;
 wire \V4/V2/A3/A1/M4/c2 ;
 wire \V4/V2/A3/A1/M4/s1 ;
 wire \V4/V2/A3/A2/c1 ;
 wire \V4/V2/A3/A2/c2 ;
 wire \V4/V2/A3/A2/c3 ;
 wire \V4/V2/A3/A2/M1/c1 ;
 wire \V4/V2/A3/A2/M1/c2 ;
 wire \V4/V2/A3/A2/M1/s1 ;
 wire \V4/V2/A3/A2/M2/c1 ;
 wire \V4/V2/A3/A2/M2/c2 ;
 wire \V4/V2/A3/A2/M2/s1 ;
 wire \V4/V2/A3/A2/M3/c1 ;
 wire \V4/V2/A3/A2/M3/c2 ;
 wire \V4/V2/A3/A2/M3/s1 ;
 wire \V4/V2/A3/A2/M4/c1 ;
 wire \V4/V2/A3/A2/M4/c2 ;
 wire \V4/V2/A3/A2/M4/s1 ;
 wire \V4/V2/V1/c1 ;
 wire \V4/V2/V1/c2 ;
 wire \V4/V2/V1/c3 ;
 wire \V4/V2/V1/overflow ;
 wire \V4/V2/V1/A1/c1 ;
 wire \V4/V2/V1/A1/c2 ;
 wire \V4/V2/V1/A1/c3 ;
 wire \V4/V2/V1/A1/M1/c1 ;
 wire \V4/V2/V1/A1/M1/c2 ;
 wire \V4/V2/V1/A1/M1/s1 ;
 wire \V4/V2/V1/A1/M2/c1 ;
 wire \V4/V2/V1/A1/M2/c2 ;
 wire \V4/V2/V1/A1/M2/s1 ;
 wire \V4/V2/V1/A1/M3/c1 ;
 wire \V4/V2/V1/A1/M3/c2 ;
 wire \V4/V2/V1/A1/M3/s1 ;
 wire \V4/V2/V1/A1/M4/c1 ;
 wire \V4/V2/V1/A1/M4/c2 ;
 wire \V4/V2/V1/A1/M4/s1 ;
 wire \V4/V2/V1/A2/c1 ;
 wire \V4/V2/V1/A2/c2 ;
 wire \V4/V2/V1/A2/c3 ;
 wire \V4/V2/V1/A2/M1/c1 ;
 wire \V4/V2/V1/A2/M1/c2 ;
 wire \V4/V2/V1/A2/M1/s1 ;
 wire \V4/V2/V1/A2/M2/c1 ;
 wire \V4/V2/V1/A2/M2/c2 ;
 wire \V4/V2/V1/A2/M2/s1 ;
 wire \V4/V2/V1/A2/M3/c1 ;
 wire \V4/V2/V1/A2/M3/c2 ;
 wire \V4/V2/V1/A2/M3/s1 ;
 wire \V4/V2/V1/A2/M4/c1 ;
 wire \V4/V2/V1/A2/M4/c2 ;
 wire \V4/V2/V1/A2/M4/s1 ;
 wire \V4/V2/V1/A3/c1 ;
 wire \V4/V2/V1/A3/c2 ;
 wire \V4/V2/V1/A3/c3 ;
 wire \V4/V2/V1/A3/M1/c1 ;
 wire \V4/V2/V1/A3/M1/c2 ;
 wire \V4/V2/V1/A3/M1/s1 ;
 wire \V4/V2/V1/A3/M2/c1 ;
 wire \V4/V2/V1/A3/M2/c2 ;
 wire \V4/V2/V1/A3/M2/s1 ;
 wire \V4/V2/V1/A3/M3/c1 ;
 wire \V4/V2/V1/A3/M3/c2 ;
 wire \V4/V2/V1/A3/M3/s1 ;
 wire \V4/V2/V1/A3/M4/c1 ;
 wire \V4/V2/V1/A3/M4/c2 ;
 wire \V4/V2/V1/A3/M4/s1 ;
 wire \V4/V2/V1/V1/w1 ;
 wire \V4/V2/V1/V1/w2 ;
 wire \V4/V2/V1/V1/w3 ;
 wire \V4/V2/V1/V1/w4 ;
 wire \V4/V2/V1/V2/w1 ;
 wire \V4/V2/V1/V2/w2 ;
 wire \V4/V2/V1/V2/w3 ;
 wire \V4/V2/V1/V2/w4 ;
 wire \V4/V2/V1/V3/w1 ;
 wire \V4/V2/V1/V3/w2 ;
 wire \V4/V2/V1/V3/w3 ;
 wire \V4/V2/V1/V3/w4 ;
 wire \V4/V2/V1/V4/w1 ;
 wire \V4/V2/V1/V4/w2 ;
 wire \V4/V2/V1/V4/w3 ;
 wire \V4/V2/V1/V4/w4 ;
 wire \V4/V2/V2/c1 ;
 wire \V4/V2/V2/c2 ;
 wire \V4/V2/V2/c3 ;
 wire \V4/V2/V2/overflow ;
 wire \V4/V2/V2/A1/c1 ;
 wire \V4/V2/V2/A1/c2 ;
 wire \V4/V2/V2/A1/c3 ;
 wire \V4/V2/V2/A1/M1/c1 ;
 wire \V4/V2/V2/A1/M1/c2 ;
 wire \V4/V2/V2/A1/M1/s1 ;
 wire \V4/V2/V2/A1/M2/c1 ;
 wire \V4/V2/V2/A1/M2/c2 ;
 wire \V4/V2/V2/A1/M2/s1 ;
 wire \V4/V2/V2/A1/M3/c1 ;
 wire \V4/V2/V2/A1/M3/c2 ;
 wire \V4/V2/V2/A1/M3/s1 ;
 wire \V4/V2/V2/A1/M4/c1 ;
 wire \V4/V2/V2/A1/M4/c2 ;
 wire \V4/V2/V2/A1/M4/s1 ;
 wire \V4/V2/V2/A2/c1 ;
 wire \V4/V2/V2/A2/c2 ;
 wire \V4/V2/V2/A2/c3 ;
 wire \V4/V2/V2/A2/M1/c1 ;
 wire \V4/V2/V2/A2/M1/c2 ;
 wire \V4/V2/V2/A2/M1/s1 ;
 wire \V4/V2/V2/A2/M2/c1 ;
 wire \V4/V2/V2/A2/M2/c2 ;
 wire \V4/V2/V2/A2/M2/s1 ;
 wire \V4/V2/V2/A2/M3/c1 ;
 wire \V4/V2/V2/A2/M3/c2 ;
 wire \V4/V2/V2/A2/M3/s1 ;
 wire \V4/V2/V2/A2/M4/c1 ;
 wire \V4/V2/V2/A2/M4/c2 ;
 wire \V4/V2/V2/A2/M4/s1 ;
 wire \V4/V2/V2/A3/c1 ;
 wire \V4/V2/V2/A3/c2 ;
 wire \V4/V2/V2/A3/c3 ;
 wire \V4/V2/V2/A3/M1/c1 ;
 wire \V4/V2/V2/A3/M1/c2 ;
 wire \V4/V2/V2/A3/M1/s1 ;
 wire \V4/V2/V2/A3/M2/c1 ;
 wire \V4/V2/V2/A3/M2/c2 ;
 wire \V4/V2/V2/A3/M2/s1 ;
 wire \V4/V2/V2/A3/M3/c1 ;
 wire \V4/V2/V2/A3/M3/c2 ;
 wire \V4/V2/V2/A3/M3/s1 ;
 wire \V4/V2/V2/A3/M4/c1 ;
 wire \V4/V2/V2/A3/M4/c2 ;
 wire \V4/V2/V2/A3/M4/s1 ;
 wire \V4/V2/V2/V1/w1 ;
 wire \V4/V2/V2/V1/w2 ;
 wire \V4/V2/V2/V1/w3 ;
 wire \V4/V2/V2/V1/w4 ;
 wire \V4/V2/V2/V2/w1 ;
 wire \V4/V2/V2/V2/w2 ;
 wire \V4/V2/V2/V2/w3 ;
 wire \V4/V2/V2/V2/w4 ;
 wire \V4/V2/V2/V3/w1 ;
 wire \V4/V2/V2/V3/w2 ;
 wire \V4/V2/V2/V3/w3 ;
 wire \V4/V2/V2/V3/w4 ;
 wire \V4/V2/V2/V4/w1 ;
 wire \V4/V2/V2/V4/w2 ;
 wire \V4/V2/V2/V4/w3 ;
 wire \V4/V2/V2/V4/w4 ;
 wire \V4/V2/V3/c1 ;
 wire \V4/V2/V3/c2 ;
 wire \V4/V2/V3/c3 ;
 wire \V4/V2/V3/overflow ;
 wire \V4/V2/V3/A1/c1 ;
 wire \V4/V2/V3/A1/c2 ;
 wire \V4/V2/V3/A1/c3 ;
 wire \V4/V2/V3/A1/M1/c1 ;
 wire \V4/V2/V3/A1/M1/c2 ;
 wire \V4/V2/V3/A1/M1/s1 ;
 wire \V4/V2/V3/A1/M2/c1 ;
 wire \V4/V2/V3/A1/M2/c2 ;
 wire \V4/V2/V3/A1/M2/s1 ;
 wire \V4/V2/V3/A1/M3/c1 ;
 wire \V4/V2/V3/A1/M3/c2 ;
 wire \V4/V2/V3/A1/M3/s1 ;
 wire \V4/V2/V3/A1/M4/c1 ;
 wire \V4/V2/V3/A1/M4/c2 ;
 wire \V4/V2/V3/A1/M4/s1 ;
 wire \V4/V2/V3/A2/c1 ;
 wire \V4/V2/V3/A2/c2 ;
 wire \V4/V2/V3/A2/c3 ;
 wire \V4/V2/V3/A2/M1/c1 ;
 wire \V4/V2/V3/A2/M1/c2 ;
 wire \V4/V2/V3/A2/M1/s1 ;
 wire \V4/V2/V3/A2/M2/c1 ;
 wire \V4/V2/V3/A2/M2/c2 ;
 wire \V4/V2/V3/A2/M2/s1 ;
 wire \V4/V2/V3/A2/M3/c1 ;
 wire \V4/V2/V3/A2/M3/c2 ;
 wire \V4/V2/V3/A2/M3/s1 ;
 wire \V4/V2/V3/A2/M4/c1 ;
 wire \V4/V2/V3/A2/M4/c2 ;
 wire \V4/V2/V3/A2/M4/s1 ;
 wire \V4/V2/V3/A3/c1 ;
 wire \V4/V2/V3/A3/c2 ;
 wire \V4/V2/V3/A3/c3 ;
 wire \V4/V2/V3/A3/M1/c1 ;
 wire \V4/V2/V3/A3/M1/c2 ;
 wire \V4/V2/V3/A3/M1/s1 ;
 wire \V4/V2/V3/A3/M2/c1 ;
 wire \V4/V2/V3/A3/M2/c2 ;
 wire \V4/V2/V3/A3/M2/s1 ;
 wire \V4/V2/V3/A3/M3/c1 ;
 wire \V4/V2/V3/A3/M3/c2 ;
 wire \V4/V2/V3/A3/M3/s1 ;
 wire \V4/V2/V3/A3/M4/c1 ;
 wire \V4/V2/V3/A3/M4/c2 ;
 wire \V4/V2/V3/A3/M4/s1 ;
 wire \V4/V2/V3/V1/w1 ;
 wire \V4/V2/V3/V1/w2 ;
 wire \V4/V2/V3/V1/w3 ;
 wire \V4/V2/V3/V1/w4 ;
 wire \V4/V2/V3/V2/w1 ;
 wire \V4/V2/V3/V2/w2 ;
 wire \V4/V2/V3/V2/w3 ;
 wire \V4/V2/V3/V2/w4 ;
 wire \V4/V2/V3/V3/w1 ;
 wire \V4/V2/V3/V3/w2 ;
 wire \V4/V2/V3/V3/w3 ;
 wire \V4/V2/V3/V3/w4 ;
 wire \V4/V2/V3/V4/w1 ;
 wire \V4/V2/V3/V4/w2 ;
 wire \V4/V2/V3/V4/w3 ;
 wire \V4/V2/V3/V4/w4 ;
 wire \V4/V2/V4/c1 ;
 wire \V4/V2/V4/c2 ;
 wire \V4/V2/V4/c3 ;
 wire \V4/V2/V4/overflow ;
 wire \V4/V2/V4/A1/c1 ;
 wire \V4/V2/V4/A1/c2 ;
 wire \V4/V2/V4/A1/c3 ;
 wire \V4/V2/V4/A1/M1/c1 ;
 wire \V4/V2/V4/A1/M1/c2 ;
 wire \V4/V2/V4/A1/M1/s1 ;
 wire \V4/V2/V4/A1/M2/c1 ;
 wire \V4/V2/V4/A1/M2/c2 ;
 wire \V4/V2/V4/A1/M2/s1 ;
 wire \V4/V2/V4/A1/M3/c1 ;
 wire \V4/V2/V4/A1/M3/c2 ;
 wire \V4/V2/V4/A1/M3/s1 ;
 wire \V4/V2/V4/A1/M4/c1 ;
 wire \V4/V2/V4/A1/M4/c2 ;
 wire \V4/V2/V4/A1/M4/s1 ;
 wire \V4/V2/V4/A2/c1 ;
 wire \V4/V2/V4/A2/c2 ;
 wire \V4/V2/V4/A2/c3 ;
 wire \V4/V2/V4/A2/M1/c1 ;
 wire \V4/V2/V4/A2/M1/c2 ;
 wire \V4/V2/V4/A2/M1/s1 ;
 wire \V4/V2/V4/A2/M2/c1 ;
 wire \V4/V2/V4/A2/M2/c2 ;
 wire \V4/V2/V4/A2/M2/s1 ;
 wire \V4/V2/V4/A2/M3/c1 ;
 wire \V4/V2/V4/A2/M3/c2 ;
 wire \V4/V2/V4/A2/M3/s1 ;
 wire \V4/V2/V4/A2/M4/c1 ;
 wire \V4/V2/V4/A2/M4/c2 ;
 wire \V4/V2/V4/A2/M4/s1 ;
 wire \V4/V2/V4/A3/c1 ;
 wire \V4/V2/V4/A3/c2 ;
 wire \V4/V2/V4/A3/c3 ;
 wire \V4/V2/V4/A3/M1/c1 ;
 wire \V4/V2/V4/A3/M1/c2 ;
 wire \V4/V2/V4/A3/M1/s1 ;
 wire \V4/V2/V4/A3/M2/c1 ;
 wire \V4/V2/V4/A3/M2/c2 ;
 wire \V4/V2/V4/A3/M2/s1 ;
 wire \V4/V2/V4/A3/M3/c1 ;
 wire \V4/V2/V4/A3/M3/c2 ;
 wire \V4/V2/V4/A3/M3/s1 ;
 wire \V4/V2/V4/A3/M4/c1 ;
 wire \V4/V2/V4/A3/M4/c2 ;
 wire \V4/V2/V4/A3/M4/s1 ;
 wire \V4/V2/V4/V1/w1 ;
 wire \V4/V2/V4/V1/w2 ;
 wire \V4/V2/V4/V1/w3 ;
 wire \V4/V2/V4/V1/w4 ;
 wire \V4/V2/V4/V2/w1 ;
 wire \V4/V2/V4/V2/w2 ;
 wire \V4/V2/V4/V2/w3 ;
 wire \V4/V2/V4/V2/w4 ;
 wire \V4/V2/V4/V3/w1 ;
 wire \V4/V2/V4/V3/w2 ;
 wire \V4/V2/V4/V3/w3 ;
 wire \V4/V2/V4/V3/w4 ;
 wire \V4/V2/V4/V4/w1 ;
 wire \V4/V2/V4/V4/w2 ;
 wire \V4/V2/V4/V4/w3 ;
 wire \V4/V2/V4/V4/w4 ;
 wire \V4/V3/c1 ;
 wire \V4/V3/c2 ;
 wire \V4/V3/c3 ;
 wire \V4/V3/overflow ;
 wire \V4/V3/A1/c1 ;
 wire \V4/V3/A1/A1/c1 ;
 wire \V4/V3/A1/A1/c2 ;
 wire \V4/V3/A1/A1/c3 ;
 wire \V4/V3/A1/A1/M1/c1 ;
 wire \V4/V3/A1/A1/M1/c2 ;
 wire \V4/V3/A1/A1/M1/s1 ;
 wire \V4/V3/A1/A1/M2/c1 ;
 wire \V4/V3/A1/A1/M2/c2 ;
 wire \V4/V3/A1/A1/M2/s1 ;
 wire \V4/V3/A1/A1/M3/c1 ;
 wire \V4/V3/A1/A1/M3/c2 ;
 wire \V4/V3/A1/A1/M3/s1 ;
 wire \V4/V3/A1/A1/M4/c1 ;
 wire \V4/V3/A1/A1/M4/c2 ;
 wire \V4/V3/A1/A1/M4/s1 ;
 wire \V4/V3/A1/A2/c1 ;
 wire \V4/V3/A1/A2/c2 ;
 wire \V4/V3/A1/A2/c3 ;
 wire \V4/V3/A1/A2/M1/c1 ;
 wire \V4/V3/A1/A2/M1/c2 ;
 wire \V4/V3/A1/A2/M1/s1 ;
 wire \V4/V3/A1/A2/M2/c1 ;
 wire \V4/V3/A1/A2/M2/c2 ;
 wire \V4/V3/A1/A2/M2/s1 ;
 wire \V4/V3/A1/A2/M3/c1 ;
 wire \V4/V3/A1/A2/M3/c2 ;
 wire \V4/V3/A1/A2/M3/s1 ;
 wire \V4/V3/A1/A2/M4/c1 ;
 wire \V4/V3/A1/A2/M4/c2 ;
 wire \V4/V3/A1/A2/M4/s1 ;
 wire \V4/V3/A2/c1 ;
 wire \V4/V3/A2/A1/c1 ;
 wire \V4/V3/A2/A1/c2 ;
 wire \V4/V3/A2/A1/c3 ;
 wire \V4/V3/A2/A1/M1/c1 ;
 wire \V4/V3/A2/A1/M1/c2 ;
 wire \V4/V3/A2/A1/M1/s1 ;
 wire \V4/V3/A2/A1/M2/c1 ;
 wire \V4/V3/A2/A1/M2/c2 ;
 wire \V4/V3/A2/A1/M2/s1 ;
 wire \V4/V3/A2/A1/M3/c1 ;
 wire \V4/V3/A2/A1/M3/c2 ;
 wire \V4/V3/A2/A1/M3/s1 ;
 wire \V4/V3/A2/A1/M4/c1 ;
 wire \V4/V3/A2/A1/M4/c2 ;
 wire \V4/V3/A2/A1/M4/s1 ;
 wire \V4/V3/A2/A2/c1 ;
 wire \V4/V3/A2/A2/c2 ;
 wire \V4/V3/A2/A2/c3 ;
 wire \V4/V3/A2/A2/M1/c1 ;
 wire \V4/V3/A2/A2/M1/c2 ;
 wire \V4/V3/A2/A2/M1/s1 ;
 wire \V4/V3/A2/A2/M2/c1 ;
 wire \V4/V3/A2/A2/M2/c2 ;
 wire \V4/V3/A2/A2/M2/s1 ;
 wire \V4/V3/A2/A2/M3/c1 ;
 wire \V4/V3/A2/A2/M3/c2 ;
 wire \V4/V3/A2/A2/M3/s1 ;
 wire \V4/V3/A2/A2/M4/c1 ;
 wire \V4/V3/A2/A2/M4/c2 ;
 wire \V4/V3/A2/A2/M4/s1 ;
 wire \V4/V3/A3/c1 ;
 wire \V4/V3/A3/A1/c1 ;
 wire \V4/V3/A3/A1/c2 ;
 wire \V4/V3/A3/A1/c3 ;
 wire \V4/V3/A3/A1/M1/c1 ;
 wire \V4/V3/A3/A1/M1/c2 ;
 wire \V4/V3/A3/A1/M1/s1 ;
 wire \V4/V3/A3/A1/M2/c1 ;
 wire \V4/V3/A3/A1/M2/c2 ;
 wire \V4/V3/A3/A1/M2/s1 ;
 wire \V4/V3/A3/A1/M3/c1 ;
 wire \V4/V3/A3/A1/M3/c2 ;
 wire \V4/V3/A3/A1/M3/s1 ;
 wire \V4/V3/A3/A1/M4/c1 ;
 wire \V4/V3/A3/A1/M4/c2 ;
 wire \V4/V3/A3/A1/M4/s1 ;
 wire \V4/V3/A3/A2/c1 ;
 wire \V4/V3/A3/A2/c2 ;
 wire \V4/V3/A3/A2/c3 ;
 wire \V4/V3/A3/A2/M1/c1 ;
 wire \V4/V3/A3/A2/M1/c2 ;
 wire \V4/V3/A3/A2/M1/s1 ;
 wire \V4/V3/A3/A2/M2/c1 ;
 wire \V4/V3/A3/A2/M2/c2 ;
 wire \V4/V3/A3/A2/M2/s1 ;
 wire \V4/V3/A3/A2/M3/c1 ;
 wire \V4/V3/A3/A2/M3/c2 ;
 wire \V4/V3/A3/A2/M3/s1 ;
 wire \V4/V3/A3/A2/M4/c1 ;
 wire \V4/V3/A3/A2/M4/c2 ;
 wire \V4/V3/A3/A2/M4/s1 ;
 wire \V4/V3/V1/c1 ;
 wire \V4/V3/V1/c2 ;
 wire \V4/V3/V1/c3 ;
 wire \V4/V3/V1/overflow ;
 wire \V4/V3/V1/A1/c1 ;
 wire \V4/V3/V1/A1/c2 ;
 wire \V4/V3/V1/A1/c3 ;
 wire \V4/V3/V1/A1/M1/c1 ;
 wire \V4/V3/V1/A1/M1/c2 ;
 wire \V4/V3/V1/A1/M1/s1 ;
 wire \V4/V3/V1/A1/M2/c1 ;
 wire \V4/V3/V1/A1/M2/c2 ;
 wire \V4/V3/V1/A1/M2/s1 ;
 wire \V4/V3/V1/A1/M3/c1 ;
 wire \V4/V3/V1/A1/M3/c2 ;
 wire \V4/V3/V1/A1/M3/s1 ;
 wire \V4/V3/V1/A1/M4/c1 ;
 wire \V4/V3/V1/A1/M4/c2 ;
 wire \V4/V3/V1/A1/M4/s1 ;
 wire \V4/V3/V1/A2/c1 ;
 wire \V4/V3/V1/A2/c2 ;
 wire \V4/V3/V1/A2/c3 ;
 wire \V4/V3/V1/A2/M1/c1 ;
 wire \V4/V3/V1/A2/M1/c2 ;
 wire \V4/V3/V1/A2/M1/s1 ;
 wire \V4/V3/V1/A2/M2/c1 ;
 wire \V4/V3/V1/A2/M2/c2 ;
 wire \V4/V3/V1/A2/M2/s1 ;
 wire \V4/V3/V1/A2/M3/c1 ;
 wire \V4/V3/V1/A2/M3/c2 ;
 wire \V4/V3/V1/A2/M3/s1 ;
 wire \V4/V3/V1/A2/M4/c1 ;
 wire \V4/V3/V1/A2/M4/c2 ;
 wire \V4/V3/V1/A2/M4/s1 ;
 wire \V4/V3/V1/A3/c1 ;
 wire \V4/V3/V1/A3/c2 ;
 wire \V4/V3/V1/A3/c3 ;
 wire \V4/V3/V1/A3/M1/c1 ;
 wire \V4/V3/V1/A3/M1/c2 ;
 wire \V4/V3/V1/A3/M1/s1 ;
 wire \V4/V3/V1/A3/M2/c1 ;
 wire \V4/V3/V1/A3/M2/c2 ;
 wire \V4/V3/V1/A3/M2/s1 ;
 wire \V4/V3/V1/A3/M3/c1 ;
 wire \V4/V3/V1/A3/M3/c2 ;
 wire \V4/V3/V1/A3/M3/s1 ;
 wire \V4/V3/V1/A3/M4/c1 ;
 wire \V4/V3/V1/A3/M4/c2 ;
 wire \V4/V3/V1/A3/M4/s1 ;
 wire \V4/V3/V1/V1/w1 ;
 wire \V4/V3/V1/V1/w2 ;
 wire \V4/V3/V1/V1/w3 ;
 wire \V4/V3/V1/V1/w4 ;
 wire \V4/V3/V1/V2/w1 ;
 wire \V4/V3/V1/V2/w2 ;
 wire \V4/V3/V1/V2/w3 ;
 wire \V4/V3/V1/V2/w4 ;
 wire \V4/V3/V1/V3/w1 ;
 wire \V4/V3/V1/V3/w2 ;
 wire \V4/V3/V1/V3/w3 ;
 wire \V4/V3/V1/V3/w4 ;
 wire \V4/V3/V1/V4/w1 ;
 wire \V4/V3/V1/V4/w2 ;
 wire \V4/V3/V1/V4/w3 ;
 wire \V4/V3/V1/V4/w4 ;
 wire \V4/V3/V2/c1 ;
 wire \V4/V3/V2/c2 ;
 wire \V4/V3/V2/c3 ;
 wire \V4/V3/V2/overflow ;
 wire \V4/V3/V2/A1/c1 ;
 wire \V4/V3/V2/A1/c2 ;
 wire \V4/V3/V2/A1/c3 ;
 wire \V4/V3/V2/A1/M1/c1 ;
 wire \V4/V3/V2/A1/M1/c2 ;
 wire \V4/V3/V2/A1/M1/s1 ;
 wire \V4/V3/V2/A1/M2/c1 ;
 wire \V4/V3/V2/A1/M2/c2 ;
 wire \V4/V3/V2/A1/M2/s1 ;
 wire \V4/V3/V2/A1/M3/c1 ;
 wire \V4/V3/V2/A1/M3/c2 ;
 wire \V4/V3/V2/A1/M3/s1 ;
 wire \V4/V3/V2/A1/M4/c1 ;
 wire \V4/V3/V2/A1/M4/c2 ;
 wire \V4/V3/V2/A1/M4/s1 ;
 wire \V4/V3/V2/A2/c1 ;
 wire \V4/V3/V2/A2/c2 ;
 wire \V4/V3/V2/A2/c3 ;
 wire \V4/V3/V2/A2/M1/c1 ;
 wire \V4/V3/V2/A2/M1/c2 ;
 wire \V4/V3/V2/A2/M1/s1 ;
 wire \V4/V3/V2/A2/M2/c1 ;
 wire \V4/V3/V2/A2/M2/c2 ;
 wire \V4/V3/V2/A2/M2/s1 ;
 wire \V4/V3/V2/A2/M3/c1 ;
 wire \V4/V3/V2/A2/M3/c2 ;
 wire \V4/V3/V2/A2/M3/s1 ;
 wire \V4/V3/V2/A2/M4/c1 ;
 wire \V4/V3/V2/A2/M4/c2 ;
 wire \V4/V3/V2/A2/M4/s1 ;
 wire \V4/V3/V2/A3/c1 ;
 wire \V4/V3/V2/A3/c2 ;
 wire \V4/V3/V2/A3/c3 ;
 wire \V4/V3/V2/A3/M1/c1 ;
 wire \V4/V3/V2/A3/M1/c2 ;
 wire \V4/V3/V2/A3/M1/s1 ;
 wire \V4/V3/V2/A3/M2/c1 ;
 wire \V4/V3/V2/A3/M2/c2 ;
 wire \V4/V3/V2/A3/M2/s1 ;
 wire \V4/V3/V2/A3/M3/c1 ;
 wire \V4/V3/V2/A3/M3/c2 ;
 wire \V4/V3/V2/A3/M3/s1 ;
 wire \V4/V3/V2/A3/M4/c1 ;
 wire \V4/V3/V2/A3/M4/c2 ;
 wire \V4/V3/V2/A3/M4/s1 ;
 wire \V4/V3/V2/V1/w1 ;
 wire \V4/V3/V2/V1/w2 ;
 wire \V4/V3/V2/V1/w3 ;
 wire \V4/V3/V2/V1/w4 ;
 wire \V4/V3/V2/V2/w1 ;
 wire \V4/V3/V2/V2/w2 ;
 wire \V4/V3/V2/V2/w3 ;
 wire \V4/V3/V2/V2/w4 ;
 wire \V4/V3/V2/V3/w1 ;
 wire \V4/V3/V2/V3/w2 ;
 wire \V4/V3/V2/V3/w3 ;
 wire \V4/V3/V2/V3/w4 ;
 wire \V4/V3/V2/V4/w1 ;
 wire \V4/V3/V2/V4/w2 ;
 wire \V4/V3/V2/V4/w3 ;
 wire \V4/V3/V2/V4/w4 ;
 wire \V4/V3/V3/c1 ;
 wire \V4/V3/V3/c2 ;
 wire \V4/V3/V3/c3 ;
 wire \V4/V3/V3/overflow ;
 wire \V4/V3/V3/A1/c1 ;
 wire \V4/V3/V3/A1/c2 ;
 wire \V4/V3/V3/A1/c3 ;
 wire \V4/V3/V3/A1/M1/c1 ;
 wire \V4/V3/V3/A1/M1/c2 ;
 wire \V4/V3/V3/A1/M1/s1 ;
 wire \V4/V3/V3/A1/M2/c1 ;
 wire \V4/V3/V3/A1/M2/c2 ;
 wire \V4/V3/V3/A1/M2/s1 ;
 wire \V4/V3/V3/A1/M3/c1 ;
 wire \V4/V3/V3/A1/M3/c2 ;
 wire \V4/V3/V3/A1/M3/s1 ;
 wire \V4/V3/V3/A1/M4/c1 ;
 wire \V4/V3/V3/A1/M4/c2 ;
 wire \V4/V3/V3/A1/M4/s1 ;
 wire \V4/V3/V3/A2/c1 ;
 wire \V4/V3/V3/A2/c2 ;
 wire \V4/V3/V3/A2/c3 ;
 wire \V4/V3/V3/A2/M1/c1 ;
 wire \V4/V3/V3/A2/M1/c2 ;
 wire \V4/V3/V3/A2/M1/s1 ;
 wire \V4/V3/V3/A2/M2/c1 ;
 wire \V4/V3/V3/A2/M2/c2 ;
 wire \V4/V3/V3/A2/M2/s1 ;
 wire \V4/V3/V3/A2/M3/c1 ;
 wire \V4/V3/V3/A2/M3/c2 ;
 wire \V4/V3/V3/A2/M3/s1 ;
 wire \V4/V3/V3/A2/M4/c1 ;
 wire \V4/V3/V3/A2/M4/c2 ;
 wire \V4/V3/V3/A2/M4/s1 ;
 wire \V4/V3/V3/A3/c1 ;
 wire \V4/V3/V3/A3/c2 ;
 wire \V4/V3/V3/A3/c3 ;
 wire \V4/V3/V3/A3/M1/c1 ;
 wire \V4/V3/V3/A3/M1/c2 ;
 wire \V4/V3/V3/A3/M1/s1 ;
 wire \V4/V3/V3/A3/M2/c1 ;
 wire \V4/V3/V3/A3/M2/c2 ;
 wire \V4/V3/V3/A3/M2/s1 ;
 wire \V4/V3/V3/A3/M3/c1 ;
 wire \V4/V3/V3/A3/M3/c2 ;
 wire \V4/V3/V3/A3/M3/s1 ;
 wire \V4/V3/V3/A3/M4/c1 ;
 wire \V4/V3/V3/A3/M4/c2 ;
 wire \V4/V3/V3/A3/M4/s1 ;
 wire \V4/V3/V3/V1/w1 ;
 wire \V4/V3/V3/V1/w2 ;
 wire \V4/V3/V3/V1/w3 ;
 wire \V4/V3/V3/V1/w4 ;
 wire \V4/V3/V3/V2/w1 ;
 wire \V4/V3/V3/V2/w2 ;
 wire \V4/V3/V3/V2/w3 ;
 wire \V4/V3/V3/V2/w4 ;
 wire \V4/V3/V3/V3/w1 ;
 wire \V4/V3/V3/V3/w2 ;
 wire \V4/V3/V3/V3/w3 ;
 wire \V4/V3/V3/V3/w4 ;
 wire \V4/V3/V3/V4/w1 ;
 wire \V4/V3/V3/V4/w2 ;
 wire \V4/V3/V3/V4/w3 ;
 wire \V4/V3/V3/V4/w4 ;
 wire \V4/V3/V4/c1 ;
 wire \V4/V3/V4/c2 ;
 wire \V4/V3/V4/c3 ;
 wire \V4/V3/V4/overflow ;
 wire \V4/V3/V4/A1/c1 ;
 wire \V4/V3/V4/A1/c2 ;
 wire \V4/V3/V4/A1/c3 ;
 wire \V4/V3/V4/A1/M1/c1 ;
 wire \V4/V3/V4/A1/M1/c2 ;
 wire \V4/V3/V4/A1/M1/s1 ;
 wire \V4/V3/V4/A1/M2/c1 ;
 wire \V4/V3/V4/A1/M2/c2 ;
 wire \V4/V3/V4/A1/M2/s1 ;
 wire \V4/V3/V4/A1/M3/c1 ;
 wire \V4/V3/V4/A1/M3/c2 ;
 wire \V4/V3/V4/A1/M3/s1 ;
 wire \V4/V3/V4/A1/M4/c1 ;
 wire \V4/V3/V4/A1/M4/c2 ;
 wire \V4/V3/V4/A1/M4/s1 ;
 wire \V4/V3/V4/A2/c1 ;
 wire \V4/V3/V4/A2/c2 ;
 wire \V4/V3/V4/A2/c3 ;
 wire \V4/V3/V4/A2/M1/c1 ;
 wire \V4/V3/V4/A2/M1/c2 ;
 wire \V4/V3/V4/A2/M1/s1 ;
 wire \V4/V3/V4/A2/M2/c1 ;
 wire \V4/V3/V4/A2/M2/c2 ;
 wire \V4/V3/V4/A2/M2/s1 ;
 wire \V4/V3/V4/A2/M3/c1 ;
 wire \V4/V3/V4/A2/M3/c2 ;
 wire \V4/V3/V4/A2/M3/s1 ;
 wire \V4/V3/V4/A2/M4/c1 ;
 wire \V4/V3/V4/A2/M4/c2 ;
 wire \V4/V3/V4/A2/M4/s1 ;
 wire \V4/V3/V4/A3/c1 ;
 wire \V4/V3/V4/A3/c2 ;
 wire \V4/V3/V4/A3/c3 ;
 wire \V4/V3/V4/A3/M1/c1 ;
 wire \V4/V3/V4/A3/M1/c2 ;
 wire \V4/V3/V4/A3/M1/s1 ;
 wire \V4/V3/V4/A3/M2/c1 ;
 wire \V4/V3/V4/A3/M2/c2 ;
 wire \V4/V3/V4/A3/M2/s1 ;
 wire \V4/V3/V4/A3/M3/c1 ;
 wire \V4/V3/V4/A3/M3/c2 ;
 wire \V4/V3/V4/A3/M3/s1 ;
 wire \V4/V3/V4/A3/M4/c1 ;
 wire \V4/V3/V4/A3/M4/c2 ;
 wire \V4/V3/V4/A3/M4/s1 ;
 wire \V4/V3/V4/V1/w1 ;
 wire \V4/V3/V4/V1/w2 ;
 wire \V4/V3/V4/V1/w3 ;
 wire \V4/V3/V4/V1/w4 ;
 wire \V4/V3/V4/V2/w1 ;
 wire \V4/V3/V4/V2/w2 ;
 wire \V4/V3/V4/V2/w3 ;
 wire \V4/V3/V4/V2/w4 ;
 wire \V4/V3/V4/V3/w1 ;
 wire \V4/V3/V4/V3/w2 ;
 wire \V4/V3/V4/V3/w3 ;
 wire \V4/V3/V4/V3/w4 ;
 wire \V4/V3/V4/V4/w1 ;
 wire \V4/V3/V4/V4/w2 ;
 wire \V4/V3/V4/V4/w3 ;
 wire \V4/V3/V4/V4/w4 ;
 wire \V4/V4/c1 ;
 wire \V4/V4/c2 ;
 wire \V4/V4/c3 ;
 wire \V4/V4/overflow ;
 wire \V4/V4/A1/c1 ;
 wire \V4/V4/A1/A1/c1 ;
 wire \V4/V4/A1/A1/c2 ;
 wire \V4/V4/A1/A1/c3 ;
 wire \V4/V4/A1/A1/M1/c1 ;
 wire \V4/V4/A1/A1/M1/c2 ;
 wire \V4/V4/A1/A1/M1/s1 ;
 wire \V4/V4/A1/A1/M2/c1 ;
 wire \V4/V4/A1/A1/M2/c2 ;
 wire \V4/V4/A1/A1/M2/s1 ;
 wire \V4/V4/A1/A1/M3/c1 ;
 wire \V4/V4/A1/A1/M3/c2 ;
 wire \V4/V4/A1/A1/M3/s1 ;
 wire \V4/V4/A1/A1/M4/c1 ;
 wire \V4/V4/A1/A1/M4/c2 ;
 wire \V4/V4/A1/A1/M4/s1 ;
 wire \V4/V4/A1/A2/c1 ;
 wire \V4/V4/A1/A2/c2 ;
 wire \V4/V4/A1/A2/c3 ;
 wire \V4/V4/A1/A2/M1/c1 ;
 wire \V4/V4/A1/A2/M1/c2 ;
 wire \V4/V4/A1/A2/M1/s1 ;
 wire \V4/V4/A1/A2/M2/c1 ;
 wire \V4/V4/A1/A2/M2/c2 ;
 wire \V4/V4/A1/A2/M2/s1 ;
 wire \V4/V4/A1/A2/M3/c1 ;
 wire \V4/V4/A1/A2/M3/c2 ;
 wire \V4/V4/A1/A2/M3/s1 ;
 wire \V4/V4/A1/A2/M4/c1 ;
 wire \V4/V4/A1/A2/M4/c2 ;
 wire \V4/V4/A1/A2/M4/s1 ;
 wire \V4/V4/A2/c1 ;
 wire \V4/V4/A2/A1/c1 ;
 wire \V4/V4/A2/A1/c2 ;
 wire \V4/V4/A2/A1/c3 ;
 wire \V4/V4/A2/A1/M1/c1 ;
 wire \V4/V4/A2/A1/M1/c2 ;
 wire \V4/V4/A2/A1/M1/s1 ;
 wire \V4/V4/A2/A1/M2/c1 ;
 wire \V4/V4/A2/A1/M2/c2 ;
 wire \V4/V4/A2/A1/M2/s1 ;
 wire \V4/V4/A2/A1/M3/c1 ;
 wire \V4/V4/A2/A1/M3/c2 ;
 wire \V4/V4/A2/A1/M3/s1 ;
 wire \V4/V4/A2/A1/M4/c1 ;
 wire \V4/V4/A2/A1/M4/c2 ;
 wire \V4/V4/A2/A1/M4/s1 ;
 wire \V4/V4/A2/A2/c1 ;
 wire \V4/V4/A2/A2/c2 ;
 wire \V4/V4/A2/A2/c3 ;
 wire \V4/V4/A2/A2/M1/c1 ;
 wire \V4/V4/A2/A2/M1/c2 ;
 wire \V4/V4/A2/A2/M1/s1 ;
 wire \V4/V4/A2/A2/M2/c1 ;
 wire \V4/V4/A2/A2/M2/c2 ;
 wire \V4/V4/A2/A2/M2/s1 ;
 wire \V4/V4/A2/A2/M3/c1 ;
 wire \V4/V4/A2/A2/M3/c2 ;
 wire \V4/V4/A2/A2/M3/s1 ;
 wire \V4/V4/A2/A2/M4/c1 ;
 wire \V4/V4/A2/A2/M4/c2 ;
 wire \V4/V4/A2/A2/M4/s1 ;
 wire \V4/V4/A3/c1 ;
 wire \V4/V4/A3/A1/c1 ;
 wire \V4/V4/A3/A1/c2 ;
 wire \V4/V4/A3/A1/c3 ;
 wire \V4/V4/A3/A1/M1/c1 ;
 wire \V4/V4/A3/A1/M1/c2 ;
 wire \V4/V4/A3/A1/M1/s1 ;
 wire \V4/V4/A3/A1/M2/c1 ;
 wire \V4/V4/A3/A1/M2/c2 ;
 wire \V4/V4/A3/A1/M2/s1 ;
 wire \V4/V4/A3/A1/M3/c1 ;
 wire \V4/V4/A3/A1/M3/c2 ;
 wire \V4/V4/A3/A1/M3/s1 ;
 wire \V4/V4/A3/A1/M4/c1 ;
 wire \V4/V4/A3/A1/M4/c2 ;
 wire \V4/V4/A3/A1/M4/s1 ;
 wire \V4/V4/A3/A2/c1 ;
 wire \V4/V4/A3/A2/c2 ;
 wire \V4/V4/A3/A2/c3 ;
 wire \V4/V4/A3/A2/M1/c1 ;
 wire \V4/V4/A3/A2/M1/c2 ;
 wire \V4/V4/A3/A2/M1/s1 ;
 wire \V4/V4/A3/A2/M2/c1 ;
 wire \V4/V4/A3/A2/M2/c2 ;
 wire \V4/V4/A3/A2/M2/s1 ;
 wire \V4/V4/A3/A2/M3/c1 ;
 wire \V4/V4/A3/A2/M3/c2 ;
 wire \V4/V4/A3/A2/M3/s1 ;
 wire \V4/V4/A3/A2/M4/c1 ;
 wire \V4/V4/A3/A2/M4/c2 ;
 wire \V4/V4/A3/A2/M4/s1 ;
 wire \V4/V4/V1/c1 ;
 wire \V4/V4/V1/c2 ;
 wire \V4/V4/V1/c3 ;
 wire \V4/V4/V1/overflow ;
 wire \V4/V4/V1/A1/c1 ;
 wire \V4/V4/V1/A1/c2 ;
 wire \V4/V4/V1/A1/c3 ;
 wire \V4/V4/V1/A1/M1/c1 ;
 wire \V4/V4/V1/A1/M1/c2 ;
 wire \V4/V4/V1/A1/M1/s1 ;
 wire \V4/V4/V1/A1/M2/c1 ;
 wire \V4/V4/V1/A1/M2/c2 ;
 wire \V4/V4/V1/A1/M2/s1 ;
 wire \V4/V4/V1/A1/M3/c1 ;
 wire \V4/V4/V1/A1/M3/c2 ;
 wire \V4/V4/V1/A1/M3/s1 ;
 wire \V4/V4/V1/A1/M4/c1 ;
 wire \V4/V4/V1/A1/M4/c2 ;
 wire \V4/V4/V1/A1/M4/s1 ;
 wire \V4/V4/V1/A2/c1 ;
 wire \V4/V4/V1/A2/c2 ;
 wire \V4/V4/V1/A2/c3 ;
 wire \V4/V4/V1/A2/M1/c1 ;
 wire \V4/V4/V1/A2/M1/c2 ;
 wire \V4/V4/V1/A2/M1/s1 ;
 wire \V4/V4/V1/A2/M2/c1 ;
 wire \V4/V4/V1/A2/M2/c2 ;
 wire \V4/V4/V1/A2/M2/s1 ;
 wire \V4/V4/V1/A2/M3/c1 ;
 wire \V4/V4/V1/A2/M3/c2 ;
 wire \V4/V4/V1/A2/M3/s1 ;
 wire \V4/V4/V1/A2/M4/c1 ;
 wire \V4/V4/V1/A2/M4/c2 ;
 wire \V4/V4/V1/A2/M4/s1 ;
 wire \V4/V4/V1/A3/c1 ;
 wire \V4/V4/V1/A3/c2 ;
 wire \V4/V4/V1/A3/c3 ;
 wire \V4/V4/V1/A3/M1/c1 ;
 wire \V4/V4/V1/A3/M1/c2 ;
 wire \V4/V4/V1/A3/M1/s1 ;
 wire \V4/V4/V1/A3/M2/c1 ;
 wire \V4/V4/V1/A3/M2/c2 ;
 wire \V4/V4/V1/A3/M2/s1 ;
 wire \V4/V4/V1/A3/M3/c1 ;
 wire \V4/V4/V1/A3/M3/c2 ;
 wire \V4/V4/V1/A3/M3/s1 ;
 wire \V4/V4/V1/A3/M4/c1 ;
 wire \V4/V4/V1/A3/M4/c2 ;
 wire \V4/V4/V1/A3/M4/s1 ;
 wire \V4/V4/V1/V1/w1 ;
 wire \V4/V4/V1/V1/w2 ;
 wire \V4/V4/V1/V1/w3 ;
 wire \V4/V4/V1/V1/w4 ;
 wire \V4/V4/V1/V2/w1 ;
 wire \V4/V4/V1/V2/w2 ;
 wire \V4/V4/V1/V2/w3 ;
 wire \V4/V4/V1/V2/w4 ;
 wire \V4/V4/V1/V3/w1 ;
 wire \V4/V4/V1/V3/w2 ;
 wire \V4/V4/V1/V3/w3 ;
 wire \V4/V4/V1/V3/w4 ;
 wire \V4/V4/V1/V4/w1 ;
 wire \V4/V4/V1/V4/w2 ;
 wire \V4/V4/V1/V4/w3 ;
 wire \V4/V4/V1/V4/w4 ;
 wire \V4/V4/V2/c1 ;
 wire \V4/V4/V2/c2 ;
 wire \V4/V4/V2/c3 ;
 wire \V4/V4/V2/overflow ;
 wire \V4/V4/V2/A1/c1 ;
 wire \V4/V4/V2/A1/c2 ;
 wire \V4/V4/V2/A1/c3 ;
 wire \V4/V4/V2/A1/M1/c1 ;
 wire \V4/V4/V2/A1/M1/c2 ;
 wire \V4/V4/V2/A1/M1/s1 ;
 wire \V4/V4/V2/A1/M2/c1 ;
 wire \V4/V4/V2/A1/M2/c2 ;
 wire \V4/V4/V2/A1/M2/s1 ;
 wire \V4/V4/V2/A1/M3/c1 ;
 wire \V4/V4/V2/A1/M3/c2 ;
 wire \V4/V4/V2/A1/M3/s1 ;
 wire \V4/V4/V2/A1/M4/c1 ;
 wire \V4/V4/V2/A1/M4/c2 ;
 wire \V4/V4/V2/A1/M4/s1 ;
 wire \V4/V4/V2/A2/c1 ;
 wire \V4/V4/V2/A2/c2 ;
 wire \V4/V4/V2/A2/c3 ;
 wire \V4/V4/V2/A2/M1/c1 ;
 wire \V4/V4/V2/A2/M1/c2 ;
 wire \V4/V4/V2/A2/M1/s1 ;
 wire \V4/V4/V2/A2/M2/c1 ;
 wire \V4/V4/V2/A2/M2/c2 ;
 wire \V4/V4/V2/A2/M2/s1 ;
 wire \V4/V4/V2/A2/M3/c1 ;
 wire \V4/V4/V2/A2/M3/c2 ;
 wire \V4/V4/V2/A2/M3/s1 ;
 wire \V4/V4/V2/A2/M4/c1 ;
 wire \V4/V4/V2/A2/M4/c2 ;
 wire \V4/V4/V2/A2/M4/s1 ;
 wire \V4/V4/V2/A3/c1 ;
 wire \V4/V4/V2/A3/c2 ;
 wire \V4/V4/V2/A3/c3 ;
 wire \V4/V4/V2/A3/M1/c1 ;
 wire \V4/V4/V2/A3/M1/c2 ;
 wire \V4/V4/V2/A3/M1/s1 ;
 wire \V4/V4/V2/A3/M2/c1 ;
 wire \V4/V4/V2/A3/M2/c2 ;
 wire \V4/V4/V2/A3/M2/s1 ;
 wire \V4/V4/V2/A3/M3/c1 ;
 wire \V4/V4/V2/A3/M3/c2 ;
 wire \V4/V4/V2/A3/M3/s1 ;
 wire \V4/V4/V2/A3/M4/c1 ;
 wire \V4/V4/V2/A3/M4/c2 ;
 wire \V4/V4/V2/A3/M4/s1 ;
 wire \V4/V4/V2/V1/w1 ;
 wire \V4/V4/V2/V1/w2 ;
 wire \V4/V4/V2/V1/w3 ;
 wire \V4/V4/V2/V1/w4 ;
 wire \V4/V4/V2/V2/w1 ;
 wire \V4/V4/V2/V2/w2 ;
 wire \V4/V4/V2/V2/w3 ;
 wire \V4/V4/V2/V2/w4 ;
 wire \V4/V4/V2/V3/w1 ;
 wire \V4/V4/V2/V3/w2 ;
 wire \V4/V4/V2/V3/w3 ;
 wire \V4/V4/V2/V3/w4 ;
 wire \V4/V4/V2/V4/w1 ;
 wire \V4/V4/V2/V4/w2 ;
 wire \V4/V4/V2/V4/w3 ;
 wire \V4/V4/V2/V4/w4 ;
 wire \V4/V4/V3/c1 ;
 wire \V4/V4/V3/c2 ;
 wire \V4/V4/V3/c3 ;
 wire \V4/V4/V3/overflow ;
 wire \V4/V4/V3/A1/c1 ;
 wire \V4/V4/V3/A1/c2 ;
 wire \V4/V4/V3/A1/c3 ;
 wire \V4/V4/V3/A1/M1/c1 ;
 wire \V4/V4/V3/A1/M1/c2 ;
 wire \V4/V4/V3/A1/M1/s1 ;
 wire \V4/V4/V3/A1/M2/c1 ;
 wire \V4/V4/V3/A1/M2/c2 ;
 wire \V4/V4/V3/A1/M2/s1 ;
 wire \V4/V4/V3/A1/M3/c1 ;
 wire \V4/V4/V3/A1/M3/c2 ;
 wire \V4/V4/V3/A1/M3/s1 ;
 wire \V4/V4/V3/A1/M4/c1 ;
 wire \V4/V4/V3/A1/M4/c2 ;
 wire \V4/V4/V3/A1/M4/s1 ;
 wire \V4/V4/V3/A2/c1 ;
 wire \V4/V4/V3/A2/c2 ;
 wire \V4/V4/V3/A2/c3 ;
 wire \V4/V4/V3/A2/M1/c1 ;
 wire \V4/V4/V3/A2/M1/c2 ;
 wire \V4/V4/V3/A2/M1/s1 ;
 wire \V4/V4/V3/A2/M2/c1 ;
 wire \V4/V4/V3/A2/M2/c2 ;
 wire \V4/V4/V3/A2/M2/s1 ;
 wire \V4/V4/V3/A2/M3/c1 ;
 wire \V4/V4/V3/A2/M3/c2 ;
 wire \V4/V4/V3/A2/M3/s1 ;
 wire \V4/V4/V3/A2/M4/c1 ;
 wire \V4/V4/V3/A2/M4/c2 ;
 wire \V4/V4/V3/A2/M4/s1 ;
 wire \V4/V4/V3/A3/c1 ;
 wire \V4/V4/V3/A3/c2 ;
 wire \V4/V4/V3/A3/c3 ;
 wire \V4/V4/V3/A3/M1/c1 ;
 wire \V4/V4/V3/A3/M1/c2 ;
 wire \V4/V4/V3/A3/M1/s1 ;
 wire \V4/V4/V3/A3/M2/c1 ;
 wire \V4/V4/V3/A3/M2/c2 ;
 wire \V4/V4/V3/A3/M2/s1 ;
 wire \V4/V4/V3/A3/M3/c1 ;
 wire \V4/V4/V3/A3/M3/c2 ;
 wire \V4/V4/V3/A3/M3/s1 ;
 wire \V4/V4/V3/A3/M4/c1 ;
 wire \V4/V4/V3/A3/M4/c2 ;
 wire \V4/V4/V3/A3/M4/s1 ;
 wire \V4/V4/V3/V1/w1 ;
 wire \V4/V4/V3/V1/w2 ;
 wire \V4/V4/V3/V1/w3 ;
 wire \V4/V4/V3/V1/w4 ;
 wire \V4/V4/V3/V2/w1 ;
 wire \V4/V4/V3/V2/w2 ;
 wire \V4/V4/V3/V2/w3 ;
 wire \V4/V4/V3/V2/w4 ;
 wire \V4/V4/V3/V3/w1 ;
 wire \V4/V4/V3/V3/w2 ;
 wire \V4/V4/V3/V3/w3 ;
 wire \V4/V4/V3/V3/w4 ;
 wire \V4/V4/V3/V4/w1 ;
 wire \V4/V4/V3/V4/w2 ;
 wire \V4/V4/V3/V4/w3 ;
 wire \V4/V4/V3/V4/w4 ;
 wire \V4/V4/V4/c1 ;
 wire \V4/V4/V4/c2 ;
 wire \V4/V4/V4/c3 ;
 wire \V4/V4/V4/overflow ;
 wire \V4/V4/V4/A1/c1 ;
 wire \V4/V4/V4/A1/c2 ;
 wire \V4/V4/V4/A1/c3 ;
 wire \V4/V4/V4/A1/M1/c1 ;
 wire \V4/V4/V4/A1/M1/c2 ;
 wire \V4/V4/V4/A1/M1/s1 ;
 wire \V4/V4/V4/A1/M2/c1 ;
 wire \V4/V4/V4/A1/M2/c2 ;
 wire \V4/V4/V4/A1/M2/s1 ;
 wire \V4/V4/V4/A1/M3/c1 ;
 wire \V4/V4/V4/A1/M3/c2 ;
 wire \V4/V4/V4/A1/M3/s1 ;
 wire \V4/V4/V4/A1/M4/c1 ;
 wire \V4/V4/V4/A1/M4/c2 ;
 wire \V4/V4/V4/A1/M4/s1 ;
 wire \V4/V4/V4/A2/c1 ;
 wire \V4/V4/V4/A2/c2 ;
 wire \V4/V4/V4/A2/c3 ;
 wire \V4/V4/V4/A2/M1/c1 ;
 wire \V4/V4/V4/A2/M1/c2 ;
 wire \V4/V4/V4/A2/M1/s1 ;
 wire \V4/V4/V4/A2/M2/c1 ;
 wire \V4/V4/V4/A2/M2/c2 ;
 wire \V4/V4/V4/A2/M2/s1 ;
 wire \V4/V4/V4/A2/M3/c1 ;
 wire \V4/V4/V4/A2/M3/c2 ;
 wire \V4/V4/V4/A2/M3/s1 ;
 wire \V4/V4/V4/A2/M4/c1 ;
 wire \V4/V4/V4/A2/M4/c2 ;
 wire \V4/V4/V4/A2/M4/s1 ;
 wire \V4/V4/V4/A3/c1 ;
 wire \V4/V4/V4/A3/c2 ;
 wire \V4/V4/V4/A3/c3 ;
 wire \V4/V4/V4/A3/M1/c1 ;
 wire \V4/V4/V4/A3/M1/c2 ;
 wire \V4/V4/V4/A3/M1/s1 ;
 wire \V4/V4/V4/A3/M2/c1 ;
 wire \V4/V4/V4/A3/M2/c2 ;
 wire \V4/V4/V4/A3/M2/s1 ;
 wire \V4/V4/V4/A3/M3/c1 ;
 wire \V4/V4/V4/A3/M3/c2 ;
 wire \V4/V4/V4/A3/M3/s1 ;
 wire \V4/V4/V4/A3/M4/c1 ;
 wire \V4/V4/V4/A3/M4/c2 ;
 wire \V4/V4/V4/A3/M4/s1 ;
 wire \V4/V4/V4/V1/w1 ;
 wire \V4/V4/V4/V1/w2 ;
 wire \V4/V4/V4/V1/w3 ;
 wire \V4/V4/V4/V1/w4 ;
 wire \V4/V4/V4/V2/w1 ;
 wire \V4/V4/V4/V2/w2 ;
 wire \V4/V4/V4/V2/w3 ;
 wire \V4/V4/V4/V2/w4 ;
 wire \V4/V4/V4/V3/w1 ;
 wire \V4/V4/V4/V3/w2 ;
 wire \V4/V4/V4/V3/w3 ;
 wire \V4/V4/V4/V3/w4 ;
 wire \V4/V4/V4/V4/w1 ;
 wire \V4/V4/V4/V4/w2 ;
 wire \V4/V4/V4/V4/w3 ;
 wire \V4/V4/V4/V4/w4 ;
 wire [3:0] \V1/V1/V1/s1 ;
 wire [3:0] \V1/V1/V1/s2 ;
 wire [3:0] \V1/V1/V1/v1 ;
 wire [3:0] \V1/V1/V1/v2 ;
 wire [3:0] \V1/V1/V1/v3 ;
 wire [3:0] \V1/V1/V1/v4 ;
 wire [3:0] \V1/V1/V2/s1 ;
 wire [3:0] \V1/V1/V2/s2 ;
 wire [3:0] \V1/V1/V2/v1 ;
 wire [3:0] \V1/V1/V2/v2 ;
 wire [3:0] \V1/V1/V2/v3 ;
 wire [3:0] \V1/V1/V2/v4 ;
 wire [3:0] \V1/V1/V3/s1 ;
 wire [3:0] \V1/V1/V3/s2 ;
 wire [3:0] \V1/V1/V3/v1 ;
 wire [3:0] \V1/V1/V3/v2 ;
 wire [3:0] \V1/V1/V3/v3 ;
 wire [3:0] \V1/V1/V3/v4 ;
 wire [3:0] \V1/V1/V4/s1 ;
 wire [3:0] \V1/V1/V4/s2 ;
 wire [3:0] \V1/V1/V4/v1 ;
 wire [3:0] \V1/V1/V4/v2 ;
 wire [3:0] \V1/V1/V4/v3 ;
 wire [3:0] \V1/V1/V4/v4 ;
 wire [7:0] \V1/V1/s1 ;
 wire [7:0] \V1/V1/s2 ;
 wire [7:0] \V1/V1/v1 ;
 wire [7:0] \V1/V1/v2 ;
 wire [7:0] \V1/V1/v3 ;
 wire [7:0] \V1/V1/v4 ;
 wire [3:0] \V1/V2/V1/s1 ;
 wire [3:0] \V1/V2/V1/s2 ;
 wire [3:0] \V1/V2/V1/v1 ;
 wire [3:0] \V1/V2/V1/v2 ;
 wire [3:0] \V1/V2/V1/v3 ;
 wire [3:0] \V1/V2/V1/v4 ;
 wire [3:0] \V1/V2/V2/s1 ;
 wire [3:0] \V1/V2/V2/s2 ;
 wire [3:0] \V1/V2/V2/v1 ;
 wire [3:0] \V1/V2/V2/v2 ;
 wire [3:0] \V1/V2/V2/v3 ;
 wire [3:0] \V1/V2/V2/v4 ;
 wire [3:0] \V1/V2/V3/s1 ;
 wire [3:0] \V1/V2/V3/s2 ;
 wire [3:0] \V1/V2/V3/v1 ;
 wire [3:0] \V1/V2/V3/v2 ;
 wire [3:0] \V1/V2/V3/v3 ;
 wire [3:0] \V1/V2/V3/v4 ;
 wire [3:0] \V1/V2/V4/s1 ;
 wire [3:0] \V1/V2/V4/s2 ;
 wire [3:0] \V1/V2/V4/v1 ;
 wire [3:0] \V1/V2/V4/v2 ;
 wire [3:0] \V1/V2/V4/v3 ;
 wire [3:0] \V1/V2/V4/v4 ;
 wire [7:0] \V1/V2/s1 ;
 wire [7:0] \V1/V2/s2 ;
 wire [7:0] \V1/V2/v1 ;
 wire [7:0] \V1/V2/v2 ;
 wire [7:0] \V1/V2/v3 ;
 wire [7:0] \V1/V2/v4 ;
 wire [3:0] \V1/V3/V1/s1 ;
 wire [3:0] \V1/V3/V1/s2 ;
 wire [3:0] \V1/V3/V1/v1 ;
 wire [3:0] \V1/V3/V1/v2 ;
 wire [3:0] \V1/V3/V1/v3 ;
 wire [3:0] \V1/V3/V1/v4 ;
 wire [3:0] \V1/V3/V2/s1 ;
 wire [3:0] \V1/V3/V2/s2 ;
 wire [3:0] \V1/V3/V2/v1 ;
 wire [3:0] \V1/V3/V2/v2 ;
 wire [3:0] \V1/V3/V2/v3 ;
 wire [3:0] \V1/V3/V2/v4 ;
 wire [3:0] \V1/V3/V3/s1 ;
 wire [3:0] \V1/V3/V3/s2 ;
 wire [3:0] \V1/V3/V3/v1 ;
 wire [3:0] \V1/V3/V3/v2 ;
 wire [3:0] \V1/V3/V3/v3 ;
 wire [3:0] \V1/V3/V3/v4 ;
 wire [3:0] \V1/V3/V4/s1 ;
 wire [3:0] \V1/V3/V4/s2 ;
 wire [3:0] \V1/V3/V4/v1 ;
 wire [3:0] \V1/V3/V4/v2 ;
 wire [3:0] \V1/V3/V4/v3 ;
 wire [3:0] \V1/V3/V4/v4 ;
 wire [7:0] \V1/V3/s1 ;
 wire [7:0] \V1/V3/s2 ;
 wire [7:0] \V1/V3/v1 ;
 wire [7:0] \V1/V3/v2 ;
 wire [7:0] \V1/V3/v3 ;
 wire [7:0] \V1/V3/v4 ;
 wire [3:0] \V1/V4/V1/s1 ;
 wire [3:0] \V1/V4/V1/s2 ;
 wire [3:0] \V1/V4/V1/v1 ;
 wire [3:0] \V1/V4/V1/v2 ;
 wire [3:0] \V1/V4/V1/v3 ;
 wire [3:0] \V1/V4/V1/v4 ;
 wire [3:0] \V1/V4/V2/s1 ;
 wire [3:0] \V1/V4/V2/s2 ;
 wire [3:0] \V1/V4/V2/v1 ;
 wire [3:0] \V1/V4/V2/v2 ;
 wire [3:0] \V1/V4/V2/v3 ;
 wire [3:0] \V1/V4/V2/v4 ;
 wire [3:0] \V1/V4/V3/s1 ;
 wire [3:0] \V1/V4/V3/s2 ;
 wire [3:0] \V1/V4/V3/v1 ;
 wire [3:0] \V1/V4/V3/v2 ;
 wire [3:0] \V1/V4/V3/v3 ;
 wire [3:0] \V1/V4/V3/v4 ;
 wire [3:0] \V1/V4/V4/s1 ;
 wire [3:0] \V1/V4/V4/s2 ;
 wire [3:0] \V1/V4/V4/v1 ;
 wire [3:0] \V1/V4/V4/v2 ;
 wire [3:0] \V1/V4/V4/v3 ;
 wire [3:0] \V1/V4/V4/v4 ;
 wire [7:0] \V1/V4/s1 ;
 wire [7:0] \V1/V4/s2 ;
 wire [7:0] \V1/V4/v1 ;
 wire [7:0] \V1/V4/v2 ;
 wire [7:0] \V1/V4/v3 ;
 wire [7:0] \V1/V4/v4 ;
 wire [15:0] \V1/s1 ;
 wire [15:0] \V1/s2 ;
 wire [15:0] \V1/v1 ;
 wire [15:0] \V1/v2 ;
 wire [15:0] \V1/v3 ;
 wire [15:0] \V1/v4 ;
 wire [3:0] \V2/V1/V1/s1 ;
 wire [3:0] \V2/V1/V1/s2 ;
 wire [3:0] \V2/V1/V1/v1 ;
 wire [3:0] \V2/V1/V1/v2 ;
 wire [3:0] \V2/V1/V1/v3 ;
 wire [3:0] \V2/V1/V1/v4 ;
 wire [3:0] \V2/V1/V2/s1 ;
 wire [3:0] \V2/V1/V2/s2 ;
 wire [3:0] \V2/V1/V2/v1 ;
 wire [3:0] \V2/V1/V2/v2 ;
 wire [3:0] \V2/V1/V2/v3 ;
 wire [3:0] \V2/V1/V2/v4 ;
 wire [3:0] \V2/V1/V3/s1 ;
 wire [3:0] \V2/V1/V3/s2 ;
 wire [3:0] \V2/V1/V3/v1 ;
 wire [3:0] \V2/V1/V3/v2 ;
 wire [3:0] \V2/V1/V3/v3 ;
 wire [3:0] \V2/V1/V3/v4 ;
 wire [3:0] \V2/V1/V4/s1 ;
 wire [3:0] \V2/V1/V4/s2 ;
 wire [3:0] \V2/V1/V4/v1 ;
 wire [3:0] \V2/V1/V4/v2 ;
 wire [3:0] \V2/V1/V4/v3 ;
 wire [3:0] \V2/V1/V4/v4 ;
 wire [7:0] \V2/V1/s1 ;
 wire [7:0] \V2/V1/s2 ;
 wire [7:0] \V2/V1/v1 ;
 wire [7:0] \V2/V1/v2 ;
 wire [7:0] \V2/V1/v3 ;
 wire [7:0] \V2/V1/v4 ;
 wire [3:0] \V2/V2/V1/s1 ;
 wire [3:0] \V2/V2/V1/s2 ;
 wire [3:0] \V2/V2/V1/v1 ;
 wire [3:0] \V2/V2/V1/v2 ;
 wire [3:0] \V2/V2/V1/v3 ;
 wire [3:0] \V2/V2/V1/v4 ;
 wire [3:0] \V2/V2/V2/s1 ;
 wire [3:0] \V2/V2/V2/s2 ;
 wire [3:0] \V2/V2/V2/v1 ;
 wire [3:0] \V2/V2/V2/v2 ;
 wire [3:0] \V2/V2/V2/v3 ;
 wire [3:0] \V2/V2/V2/v4 ;
 wire [3:0] \V2/V2/V3/s1 ;
 wire [3:0] \V2/V2/V3/s2 ;
 wire [3:0] \V2/V2/V3/v1 ;
 wire [3:0] \V2/V2/V3/v2 ;
 wire [3:0] \V2/V2/V3/v3 ;
 wire [3:0] \V2/V2/V3/v4 ;
 wire [3:0] \V2/V2/V4/s1 ;
 wire [3:0] \V2/V2/V4/s2 ;
 wire [3:0] \V2/V2/V4/v1 ;
 wire [3:0] \V2/V2/V4/v2 ;
 wire [3:0] \V2/V2/V4/v3 ;
 wire [3:0] \V2/V2/V4/v4 ;
 wire [7:0] \V2/V2/s1 ;
 wire [7:0] \V2/V2/s2 ;
 wire [7:0] \V2/V2/v1 ;
 wire [7:0] \V2/V2/v2 ;
 wire [7:0] \V2/V2/v3 ;
 wire [7:0] \V2/V2/v4 ;
 wire [3:0] \V2/V3/V1/s1 ;
 wire [3:0] \V2/V3/V1/s2 ;
 wire [3:0] \V2/V3/V1/v1 ;
 wire [3:0] \V2/V3/V1/v2 ;
 wire [3:0] \V2/V3/V1/v3 ;
 wire [3:0] \V2/V3/V1/v4 ;
 wire [3:0] \V2/V3/V2/s1 ;
 wire [3:0] \V2/V3/V2/s2 ;
 wire [3:0] \V2/V3/V2/v1 ;
 wire [3:0] \V2/V3/V2/v2 ;
 wire [3:0] \V2/V3/V2/v3 ;
 wire [3:0] \V2/V3/V2/v4 ;
 wire [3:0] \V2/V3/V3/s1 ;
 wire [3:0] \V2/V3/V3/s2 ;
 wire [3:0] \V2/V3/V3/v1 ;
 wire [3:0] \V2/V3/V3/v2 ;
 wire [3:0] \V2/V3/V3/v3 ;
 wire [3:0] \V2/V3/V3/v4 ;
 wire [3:0] \V2/V3/V4/s1 ;
 wire [3:0] \V2/V3/V4/s2 ;
 wire [3:0] \V2/V3/V4/v1 ;
 wire [3:0] \V2/V3/V4/v2 ;
 wire [3:0] \V2/V3/V4/v3 ;
 wire [3:0] \V2/V3/V4/v4 ;
 wire [7:0] \V2/V3/s1 ;
 wire [7:0] \V2/V3/s2 ;
 wire [7:0] \V2/V3/v1 ;
 wire [7:0] \V2/V3/v2 ;
 wire [7:0] \V2/V3/v3 ;
 wire [7:0] \V2/V3/v4 ;
 wire [3:0] \V2/V4/V1/s1 ;
 wire [3:0] \V2/V4/V1/s2 ;
 wire [3:0] \V2/V4/V1/v1 ;
 wire [3:0] \V2/V4/V1/v2 ;
 wire [3:0] \V2/V4/V1/v3 ;
 wire [3:0] \V2/V4/V1/v4 ;
 wire [3:0] \V2/V4/V2/s1 ;
 wire [3:0] \V2/V4/V2/s2 ;
 wire [3:0] \V2/V4/V2/v1 ;
 wire [3:0] \V2/V4/V2/v2 ;
 wire [3:0] \V2/V4/V2/v3 ;
 wire [3:0] \V2/V4/V2/v4 ;
 wire [3:0] \V2/V4/V3/s1 ;
 wire [3:0] \V2/V4/V3/s2 ;
 wire [3:0] \V2/V4/V3/v1 ;
 wire [3:0] \V2/V4/V3/v2 ;
 wire [3:0] \V2/V4/V3/v3 ;
 wire [3:0] \V2/V4/V3/v4 ;
 wire [3:0] \V2/V4/V4/s1 ;
 wire [3:0] \V2/V4/V4/s2 ;
 wire [3:0] \V2/V4/V4/v1 ;
 wire [3:0] \V2/V4/V4/v2 ;
 wire [3:0] \V2/V4/V4/v3 ;
 wire [3:0] \V2/V4/V4/v4 ;
 wire [7:0] \V2/V4/s1 ;
 wire [7:0] \V2/V4/s2 ;
 wire [7:0] \V2/V4/v1 ;
 wire [7:0] \V2/V4/v2 ;
 wire [7:0] \V2/V4/v3 ;
 wire [7:0] \V2/V4/v4 ;
 wire [15:0] \V2/s1 ;
 wire [15:0] \V2/s2 ;
 wire [15:0] \V2/v1 ;
 wire [15:0] \V2/v2 ;
 wire [15:0] \V2/v3 ;
 wire [15:0] \V2/v4 ;
 wire [3:0] \V3/V1/V1/s1 ;
 wire [3:0] \V3/V1/V1/s2 ;
 wire [3:0] \V3/V1/V1/v1 ;
 wire [3:0] \V3/V1/V1/v2 ;
 wire [3:0] \V3/V1/V1/v3 ;
 wire [3:0] \V3/V1/V1/v4 ;
 wire [3:0] \V3/V1/V2/s1 ;
 wire [3:0] \V3/V1/V2/s2 ;
 wire [3:0] \V3/V1/V2/v1 ;
 wire [3:0] \V3/V1/V2/v2 ;
 wire [3:0] \V3/V1/V2/v3 ;
 wire [3:0] \V3/V1/V2/v4 ;
 wire [3:0] \V3/V1/V3/s1 ;
 wire [3:0] \V3/V1/V3/s2 ;
 wire [3:0] \V3/V1/V3/v1 ;
 wire [3:0] \V3/V1/V3/v2 ;
 wire [3:0] \V3/V1/V3/v3 ;
 wire [3:0] \V3/V1/V3/v4 ;
 wire [3:0] \V3/V1/V4/s1 ;
 wire [3:0] \V3/V1/V4/s2 ;
 wire [3:0] \V3/V1/V4/v1 ;
 wire [3:0] \V3/V1/V4/v2 ;
 wire [3:0] \V3/V1/V4/v3 ;
 wire [3:0] \V3/V1/V4/v4 ;
 wire [7:0] \V3/V1/s1 ;
 wire [7:0] \V3/V1/s2 ;
 wire [7:0] \V3/V1/v1 ;
 wire [7:0] \V3/V1/v2 ;
 wire [7:0] \V3/V1/v3 ;
 wire [7:0] \V3/V1/v4 ;
 wire [3:0] \V3/V2/V1/s1 ;
 wire [3:0] \V3/V2/V1/s2 ;
 wire [3:0] \V3/V2/V1/v1 ;
 wire [3:0] \V3/V2/V1/v2 ;
 wire [3:0] \V3/V2/V1/v3 ;
 wire [3:0] \V3/V2/V1/v4 ;
 wire [3:0] \V3/V2/V2/s1 ;
 wire [3:0] \V3/V2/V2/s2 ;
 wire [3:0] \V3/V2/V2/v1 ;
 wire [3:0] \V3/V2/V2/v2 ;
 wire [3:0] \V3/V2/V2/v3 ;
 wire [3:0] \V3/V2/V2/v4 ;
 wire [3:0] \V3/V2/V3/s1 ;
 wire [3:0] \V3/V2/V3/s2 ;
 wire [3:0] \V3/V2/V3/v1 ;
 wire [3:0] \V3/V2/V3/v2 ;
 wire [3:0] \V3/V2/V3/v3 ;
 wire [3:0] \V3/V2/V3/v4 ;
 wire [3:0] \V3/V2/V4/s1 ;
 wire [3:0] \V3/V2/V4/s2 ;
 wire [3:0] \V3/V2/V4/v1 ;
 wire [3:0] \V3/V2/V4/v2 ;
 wire [3:0] \V3/V2/V4/v3 ;
 wire [3:0] \V3/V2/V4/v4 ;
 wire [7:0] \V3/V2/s1 ;
 wire [7:0] \V3/V2/s2 ;
 wire [7:0] \V3/V2/v1 ;
 wire [7:0] \V3/V2/v2 ;
 wire [7:0] \V3/V2/v3 ;
 wire [7:0] \V3/V2/v4 ;
 wire [3:0] \V3/V3/V1/s1 ;
 wire [3:0] \V3/V3/V1/s2 ;
 wire [3:0] \V3/V3/V1/v1 ;
 wire [3:0] \V3/V3/V1/v2 ;
 wire [3:0] \V3/V3/V1/v3 ;
 wire [3:0] \V3/V3/V1/v4 ;
 wire [3:0] \V3/V3/V2/s1 ;
 wire [3:0] \V3/V3/V2/s2 ;
 wire [3:0] \V3/V3/V2/v1 ;
 wire [3:0] \V3/V3/V2/v2 ;
 wire [3:0] \V3/V3/V2/v3 ;
 wire [3:0] \V3/V3/V2/v4 ;
 wire [3:0] \V3/V3/V3/s1 ;
 wire [3:0] \V3/V3/V3/s2 ;
 wire [3:0] \V3/V3/V3/v1 ;
 wire [3:0] \V3/V3/V3/v2 ;
 wire [3:0] \V3/V3/V3/v3 ;
 wire [3:0] \V3/V3/V3/v4 ;
 wire [3:0] \V3/V3/V4/s1 ;
 wire [3:0] \V3/V3/V4/s2 ;
 wire [3:0] \V3/V3/V4/v1 ;
 wire [3:0] \V3/V3/V4/v2 ;
 wire [3:0] \V3/V3/V4/v3 ;
 wire [3:0] \V3/V3/V4/v4 ;
 wire [7:0] \V3/V3/s1 ;
 wire [7:0] \V3/V3/s2 ;
 wire [7:0] \V3/V3/v1 ;
 wire [7:0] \V3/V3/v2 ;
 wire [7:0] \V3/V3/v3 ;
 wire [7:0] \V3/V3/v4 ;
 wire [3:0] \V3/V4/V1/s1 ;
 wire [3:0] \V3/V4/V1/s2 ;
 wire [3:0] \V3/V4/V1/v1 ;
 wire [3:0] \V3/V4/V1/v2 ;
 wire [3:0] \V3/V4/V1/v3 ;
 wire [3:0] \V3/V4/V1/v4 ;
 wire [3:0] \V3/V4/V2/s1 ;
 wire [3:0] \V3/V4/V2/s2 ;
 wire [3:0] \V3/V4/V2/v1 ;
 wire [3:0] \V3/V4/V2/v2 ;
 wire [3:0] \V3/V4/V2/v3 ;
 wire [3:0] \V3/V4/V2/v4 ;
 wire [3:0] \V3/V4/V3/s1 ;
 wire [3:0] \V3/V4/V3/s2 ;
 wire [3:0] \V3/V4/V3/v1 ;
 wire [3:0] \V3/V4/V3/v2 ;
 wire [3:0] \V3/V4/V3/v3 ;
 wire [3:0] \V3/V4/V3/v4 ;
 wire [3:0] \V3/V4/V4/s1 ;
 wire [3:0] \V3/V4/V4/s2 ;
 wire [3:0] \V3/V4/V4/v1 ;
 wire [3:0] \V3/V4/V4/v2 ;
 wire [3:0] \V3/V4/V4/v3 ;
 wire [3:0] \V3/V4/V4/v4 ;
 wire [7:0] \V3/V4/s1 ;
 wire [7:0] \V3/V4/s2 ;
 wire [7:0] \V3/V4/v1 ;
 wire [7:0] \V3/V4/v2 ;
 wire [7:0] \V3/V4/v3 ;
 wire [7:0] \V3/V4/v4 ;
 wire [15:0] \V3/s1 ;
 wire [15:0] \V3/s2 ;
 wire [15:0] \V3/v1 ;
 wire [15:0] \V3/v2 ;
 wire [15:0] \V3/v3 ;
 wire [15:0] \V3/v4 ;
 wire [3:0] \V4/V1/V1/s1 ;
 wire [3:0] \V4/V1/V1/s2 ;
 wire [3:0] \V4/V1/V1/v1 ;
 wire [3:0] \V4/V1/V1/v2 ;
 wire [3:0] \V4/V1/V1/v3 ;
 wire [3:0] \V4/V1/V1/v4 ;
 wire [3:0] \V4/V1/V2/s1 ;
 wire [3:0] \V4/V1/V2/s2 ;
 wire [3:0] \V4/V1/V2/v1 ;
 wire [3:0] \V4/V1/V2/v2 ;
 wire [3:0] \V4/V1/V2/v3 ;
 wire [3:0] \V4/V1/V2/v4 ;
 wire [3:0] \V4/V1/V3/s1 ;
 wire [3:0] \V4/V1/V3/s2 ;
 wire [3:0] \V4/V1/V3/v1 ;
 wire [3:0] \V4/V1/V3/v2 ;
 wire [3:0] \V4/V1/V3/v3 ;
 wire [3:0] \V4/V1/V3/v4 ;
 wire [3:0] \V4/V1/V4/s1 ;
 wire [3:0] \V4/V1/V4/s2 ;
 wire [3:0] \V4/V1/V4/v1 ;
 wire [3:0] \V4/V1/V4/v2 ;
 wire [3:0] \V4/V1/V4/v3 ;
 wire [3:0] \V4/V1/V4/v4 ;
 wire [7:0] \V4/V1/s1 ;
 wire [7:0] \V4/V1/s2 ;
 wire [7:0] \V4/V1/v1 ;
 wire [7:0] \V4/V1/v2 ;
 wire [7:0] \V4/V1/v3 ;
 wire [7:0] \V4/V1/v4 ;
 wire [3:0] \V4/V2/V1/s1 ;
 wire [3:0] \V4/V2/V1/s2 ;
 wire [3:0] \V4/V2/V1/v1 ;
 wire [3:0] \V4/V2/V1/v2 ;
 wire [3:0] \V4/V2/V1/v3 ;
 wire [3:0] \V4/V2/V1/v4 ;
 wire [3:0] \V4/V2/V2/s1 ;
 wire [3:0] \V4/V2/V2/s2 ;
 wire [3:0] \V4/V2/V2/v1 ;
 wire [3:0] \V4/V2/V2/v2 ;
 wire [3:0] \V4/V2/V2/v3 ;
 wire [3:0] \V4/V2/V2/v4 ;
 wire [3:0] \V4/V2/V3/s1 ;
 wire [3:0] \V4/V2/V3/s2 ;
 wire [3:0] \V4/V2/V3/v1 ;
 wire [3:0] \V4/V2/V3/v2 ;
 wire [3:0] \V4/V2/V3/v3 ;
 wire [3:0] \V4/V2/V3/v4 ;
 wire [3:0] \V4/V2/V4/s1 ;
 wire [3:0] \V4/V2/V4/s2 ;
 wire [3:0] \V4/V2/V4/v1 ;
 wire [3:0] \V4/V2/V4/v2 ;
 wire [3:0] \V4/V2/V4/v3 ;
 wire [3:0] \V4/V2/V4/v4 ;
 wire [7:0] \V4/V2/s1 ;
 wire [7:0] \V4/V2/s2 ;
 wire [7:0] \V4/V2/v1 ;
 wire [7:0] \V4/V2/v2 ;
 wire [7:0] \V4/V2/v3 ;
 wire [7:0] \V4/V2/v4 ;
 wire [3:0] \V4/V3/V1/s1 ;
 wire [3:0] \V4/V3/V1/s2 ;
 wire [3:0] \V4/V3/V1/v1 ;
 wire [3:0] \V4/V3/V1/v2 ;
 wire [3:0] \V4/V3/V1/v3 ;
 wire [3:0] \V4/V3/V1/v4 ;
 wire [3:0] \V4/V3/V2/s1 ;
 wire [3:0] \V4/V3/V2/s2 ;
 wire [3:0] \V4/V3/V2/v1 ;
 wire [3:0] \V4/V3/V2/v2 ;
 wire [3:0] \V4/V3/V2/v3 ;
 wire [3:0] \V4/V3/V2/v4 ;
 wire [3:0] \V4/V3/V3/s1 ;
 wire [3:0] \V4/V3/V3/s2 ;
 wire [3:0] \V4/V3/V3/v1 ;
 wire [3:0] \V4/V3/V3/v2 ;
 wire [3:0] \V4/V3/V3/v3 ;
 wire [3:0] \V4/V3/V3/v4 ;
 wire [3:0] \V4/V3/V4/s1 ;
 wire [3:0] \V4/V3/V4/s2 ;
 wire [3:0] \V4/V3/V4/v1 ;
 wire [3:0] \V4/V3/V4/v2 ;
 wire [3:0] \V4/V3/V4/v3 ;
 wire [3:0] \V4/V3/V4/v4 ;
 wire [7:0] \V4/V3/s1 ;
 wire [7:0] \V4/V3/s2 ;
 wire [7:0] \V4/V3/v1 ;
 wire [7:0] \V4/V3/v2 ;
 wire [7:0] \V4/V3/v3 ;
 wire [7:0] \V4/V3/v4 ;
 wire [3:0] \V4/V4/V1/s1 ;
 wire [3:0] \V4/V4/V1/s2 ;
 wire [3:0] \V4/V4/V1/v1 ;
 wire [3:0] \V4/V4/V1/v2 ;
 wire [3:0] \V4/V4/V1/v3 ;
 wire [3:0] \V4/V4/V1/v4 ;
 wire [3:0] \V4/V4/V2/s1 ;
 wire [3:0] \V4/V4/V2/s2 ;
 wire [3:0] \V4/V4/V2/v1 ;
 wire [3:0] \V4/V4/V2/v2 ;
 wire [3:0] \V4/V4/V2/v3 ;
 wire [3:0] \V4/V4/V2/v4 ;
 wire [3:0] \V4/V4/V3/s1 ;
 wire [3:0] \V4/V4/V3/s2 ;
 wire [3:0] \V4/V4/V3/v1 ;
 wire [3:0] \V4/V4/V3/v2 ;
 wire [3:0] \V4/V4/V3/v3 ;
 wire [3:0] \V4/V4/V3/v4 ;
 wire [3:0] \V4/V4/V4/s1 ;
 wire [3:0] \V4/V4/V4/s2 ;
 wire [3:0] \V4/V4/V4/v1 ;
 wire [3:0] \V4/V4/V4/v2 ;
 wire [3:0] \V4/V4/V4/v3 ;
 wire [3:0] \V4/V4/V4/v4 ;
 wire [7:0] \V4/V4/s1 ;
 wire [7:0] \V4/V4/s2 ;
 wire [7:0] \V4/V4/v1 ;
 wire [7:0] \V4/V4/v2 ;
 wire [7:0] \V4/V4/v3 ;
 wire [7:0] \V4/V4/v4 ;
 wire [15:0] \V4/s1 ;
 wire [15:0] \V4/s2 ;
 wire [15:0] \V4/v1 ;
 wire [15:0] \V4/v2 ;
 wire [15:0] \V4/v3 ;
 wire [15:0] \V4/v4 ;
 wire [31:0] s1;
 wire [31:0] s2;
 wire [31:0] v1;
 wire [31:0] v2;
 wire [31:0] v3;
 wire [31:0] v4;

 AND2_X1 \A1/A1/A1/A1/M1/M1/_0_  (.A1(v2[0]),
    .A2(v3[0]),
    .ZN(\A1/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M1/M1/_1_  (.A(v2[0]),
    .B(v3[0]),
    .Z(\A1/A1/A1/A1/M1/s1 ));
 AND2_X1 \A1/A1/A1/A1/M1/M2/_0_  (.A1(\A1/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A1/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M1/M2/_1_  (.A(\A1/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(s1[0]));
 OR2_X1 \A1/A1/A1/A1/M1/_0_  (.A1(\A1/A1/A1/A1/M1/c1 ),
    .A2(\A1/A1/A1/A1/M1/c2 ),
    .ZN(\A1/A1/A1/A1/c1 ));
 AND2_X1 \A1/A1/A1/A1/M2/M1/_0_  (.A1(v2[1]),
    .A2(v3[1]),
    .ZN(\A1/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M2/M1/_1_  (.A(v2[1]),
    .B(v3[1]),
    .Z(\A1/A1/A1/A1/M2/s1 ));
 AND2_X1 \A1/A1/A1/A1/M2/M2/_0_  (.A1(\A1/A1/A1/A1/M2/s1 ),
    .A2(\A1/A1/A1/A1/c1 ),
    .ZN(\A1/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M2/M2/_1_  (.A(\A1/A1/A1/A1/M2/s1 ),
    .B(\A1/A1/A1/A1/c1 ),
    .Z(s1[1]));
 OR2_X1 \A1/A1/A1/A1/M2/_0_  (.A1(\A1/A1/A1/A1/M2/c1 ),
    .A2(\A1/A1/A1/A1/M2/c2 ),
    .ZN(\A1/A1/A1/A1/c2 ));
 AND2_X1 \A1/A1/A1/A1/M3/M1/_0_  (.A1(v2[2]),
    .A2(v3[2]),
    .ZN(\A1/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M3/M1/_1_  (.A(v2[2]),
    .B(v3[2]),
    .Z(\A1/A1/A1/A1/M3/s1 ));
 AND2_X1 \A1/A1/A1/A1/M3/M2/_0_  (.A1(\A1/A1/A1/A1/M3/s1 ),
    .A2(\A1/A1/A1/A1/c2 ),
    .ZN(\A1/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M3/M2/_1_  (.A(\A1/A1/A1/A1/M3/s1 ),
    .B(\A1/A1/A1/A1/c2 ),
    .Z(s1[2]));
 OR2_X1 \A1/A1/A1/A1/M3/_0_  (.A1(\A1/A1/A1/A1/M3/c1 ),
    .A2(\A1/A1/A1/A1/M3/c2 ),
    .ZN(\A1/A1/A1/A1/c3 ));
 AND2_X1 \A1/A1/A1/A1/M4/M1/_0_  (.A1(v2[3]),
    .A2(v3[3]),
    .ZN(\A1/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M4/M1/_1_  (.A(v2[3]),
    .B(v3[3]),
    .Z(\A1/A1/A1/A1/M4/s1 ));
 AND2_X1 \A1/A1/A1/A1/M4/M2/_0_  (.A1(\A1/A1/A1/A1/M4/s1 ),
    .A2(\A1/A1/A1/A1/c3 ),
    .ZN(\A1/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M4/M2/_1_  (.A(\A1/A1/A1/A1/M4/s1 ),
    .B(\A1/A1/A1/A1/c3 ),
    .Z(s1[3]));
 OR2_X1 \A1/A1/A1/A1/M4/_0_  (.A1(\A1/A1/A1/A1/M4/c1 ),
    .A2(\A1/A1/A1/A1/M4/c2 ),
    .ZN(\A1/A1/A1/c1 ));
 AND2_X1 \A1/A1/A1/A2/M1/M1/_0_  (.A1(v2[4]),
    .A2(v3[4]),
    .ZN(\A1/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M1/M1/_1_  (.A(v2[4]),
    .B(v3[4]),
    .Z(\A1/A1/A1/A2/M1/s1 ));
 AND2_X1 \A1/A1/A1/A2/M1/M2/_0_  (.A1(\A1/A1/A1/A2/M1/s1 ),
    .A2(\A1/A1/A1/c1 ),
    .ZN(\A1/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M1/M2/_1_  (.A(\A1/A1/A1/A2/M1/s1 ),
    .B(\A1/A1/A1/c1 ),
    .Z(s1[4]));
 OR2_X1 \A1/A1/A1/A2/M1/_0_  (.A1(\A1/A1/A1/A2/M1/c1 ),
    .A2(\A1/A1/A1/A2/M1/c2 ),
    .ZN(\A1/A1/A1/A2/c1 ));
 AND2_X1 \A1/A1/A1/A2/M2/M1/_0_  (.A1(v2[5]),
    .A2(v3[5]),
    .ZN(\A1/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M2/M1/_1_  (.A(v2[5]),
    .B(v3[5]),
    .Z(\A1/A1/A1/A2/M2/s1 ));
 AND2_X1 \A1/A1/A1/A2/M2/M2/_0_  (.A1(\A1/A1/A1/A2/M2/s1 ),
    .A2(\A1/A1/A1/A2/c1 ),
    .ZN(\A1/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M2/M2/_1_  (.A(\A1/A1/A1/A2/M2/s1 ),
    .B(\A1/A1/A1/A2/c1 ),
    .Z(s1[5]));
 OR2_X1 \A1/A1/A1/A2/M2/_0_  (.A1(\A1/A1/A1/A2/M2/c1 ),
    .A2(\A1/A1/A1/A2/M2/c2 ),
    .ZN(\A1/A1/A1/A2/c2 ));
 AND2_X1 \A1/A1/A1/A2/M3/M1/_0_  (.A1(v2[6]),
    .A2(v3[6]),
    .ZN(\A1/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M3/M1/_1_  (.A(v2[6]),
    .B(v3[6]),
    .Z(\A1/A1/A1/A2/M3/s1 ));
 AND2_X1 \A1/A1/A1/A2/M3/M2/_0_  (.A1(\A1/A1/A1/A2/M3/s1 ),
    .A2(\A1/A1/A1/A2/c2 ),
    .ZN(\A1/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M3/M2/_1_  (.A(\A1/A1/A1/A2/M3/s1 ),
    .B(\A1/A1/A1/A2/c2 ),
    .Z(s1[6]));
 OR2_X1 \A1/A1/A1/A2/M3/_0_  (.A1(\A1/A1/A1/A2/M3/c1 ),
    .A2(\A1/A1/A1/A2/M3/c2 ),
    .ZN(\A1/A1/A1/A2/c3 ));
 AND2_X1 \A1/A1/A1/A2/M4/M1/_0_  (.A1(v2[7]),
    .A2(v3[7]),
    .ZN(\A1/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M4/M1/_1_  (.A(v2[7]),
    .B(v3[7]),
    .Z(\A1/A1/A1/A2/M4/s1 ));
 AND2_X1 \A1/A1/A1/A2/M4/M2/_0_  (.A1(\A1/A1/A1/A2/M4/s1 ),
    .A2(\A1/A1/A1/A2/c3 ),
    .ZN(\A1/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M4/M2/_1_  (.A(\A1/A1/A1/A2/M4/s1 ),
    .B(\A1/A1/A1/A2/c3 ),
    .Z(s1[7]));
 OR2_X1 \A1/A1/A1/A2/M4/_0_  (.A1(\A1/A1/A1/A2/M4/c1 ),
    .A2(\A1/A1/A1/A2/M4/c2 ),
    .ZN(\A1/A1/c1 ));
 AND2_X1 \A1/A1/A2/A1/M1/M1/_0_  (.A1(v2[8]),
    .A2(v3[8]),
    .ZN(\A1/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M1/M1/_1_  (.A(v2[8]),
    .B(v3[8]),
    .Z(\A1/A1/A2/A1/M1/s1 ));
 AND2_X1 \A1/A1/A2/A1/M1/M2/_0_  (.A1(\A1/A1/A2/A1/M1/s1 ),
    .A2(\A1/A1/c1 ),
    .ZN(\A1/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M1/M2/_1_  (.A(\A1/A1/A2/A1/M1/s1 ),
    .B(\A1/A1/c1 ),
    .Z(s1[8]));
 OR2_X1 \A1/A1/A2/A1/M1/_0_  (.A1(\A1/A1/A2/A1/M1/c1 ),
    .A2(\A1/A1/A2/A1/M1/c2 ),
    .ZN(\A1/A1/A2/A1/c1 ));
 AND2_X1 \A1/A1/A2/A1/M2/M1/_0_  (.A1(v2[9]),
    .A2(v3[9]),
    .ZN(\A1/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M2/M1/_1_  (.A(v2[9]),
    .B(v3[9]),
    .Z(\A1/A1/A2/A1/M2/s1 ));
 AND2_X1 \A1/A1/A2/A1/M2/M2/_0_  (.A1(\A1/A1/A2/A1/M2/s1 ),
    .A2(\A1/A1/A2/A1/c1 ),
    .ZN(\A1/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M2/M2/_1_  (.A(\A1/A1/A2/A1/M2/s1 ),
    .B(\A1/A1/A2/A1/c1 ),
    .Z(s1[9]));
 OR2_X1 \A1/A1/A2/A1/M2/_0_  (.A1(\A1/A1/A2/A1/M2/c1 ),
    .A2(\A1/A1/A2/A1/M2/c2 ),
    .ZN(\A1/A1/A2/A1/c2 ));
 AND2_X1 \A1/A1/A2/A1/M3/M1/_0_  (.A1(v2[10]),
    .A2(v3[10]),
    .ZN(\A1/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M3/M1/_1_  (.A(v2[10]),
    .B(v3[10]),
    .Z(\A1/A1/A2/A1/M3/s1 ));
 AND2_X1 \A1/A1/A2/A1/M3/M2/_0_  (.A1(\A1/A1/A2/A1/M3/s1 ),
    .A2(\A1/A1/A2/A1/c2 ),
    .ZN(\A1/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M3/M2/_1_  (.A(\A1/A1/A2/A1/M3/s1 ),
    .B(\A1/A1/A2/A1/c2 ),
    .Z(s1[10]));
 OR2_X1 \A1/A1/A2/A1/M3/_0_  (.A1(\A1/A1/A2/A1/M3/c1 ),
    .A2(\A1/A1/A2/A1/M3/c2 ),
    .ZN(\A1/A1/A2/A1/c3 ));
 AND2_X1 \A1/A1/A2/A1/M4/M1/_0_  (.A1(v2[11]),
    .A2(v3[11]),
    .ZN(\A1/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M4/M1/_1_  (.A(v2[11]),
    .B(v3[11]),
    .Z(\A1/A1/A2/A1/M4/s1 ));
 AND2_X1 \A1/A1/A2/A1/M4/M2/_0_  (.A1(\A1/A1/A2/A1/M4/s1 ),
    .A2(\A1/A1/A2/A1/c3 ),
    .ZN(\A1/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M4/M2/_1_  (.A(\A1/A1/A2/A1/M4/s1 ),
    .B(\A1/A1/A2/A1/c3 ),
    .Z(s1[11]));
 OR2_X1 \A1/A1/A2/A1/M4/_0_  (.A1(\A1/A1/A2/A1/M4/c1 ),
    .A2(\A1/A1/A2/A1/M4/c2 ),
    .ZN(\A1/A1/A2/c1 ));
 AND2_X1 \A1/A1/A2/A2/M1/M1/_0_  (.A1(v2[12]),
    .A2(v3[12]),
    .ZN(\A1/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M1/M1/_1_  (.A(v2[12]),
    .B(v3[12]),
    .Z(\A1/A1/A2/A2/M1/s1 ));
 AND2_X1 \A1/A1/A2/A2/M1/M2/_0_  (.A1(\A1/A1/A2/A2/M1/s1 ),
    .A2(\A1/A1/A2/c1 ),
    .ZN(\A1/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M1/M2/_1_  (.A(\A1/A1/A2/A2/M1/s1 ),
    .B(\A1/A1/A2/c1 ),
    .Z(s1[12]));
 OR2_X1 \A1/A1/A2/A2/M1/_0_  (.A1(\A1/A1/A2/A2/M1/c1 ),
    .A2(\A1/A1/A2/A2/M1/c2 ),
    .ZN(\A1/A1/A2/A2/c1 ));
 AND2_X1 \A1/A1/A2/A2/M2/M1/_0_  (.A1(v2[13]),
    .A2(v3[13]),
    .ZN(\A1/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M2/M1/_1_  (.A(v2[13]),
    .B(v3[13]),
    .Z(\A1/A1/A2/A2/M2/s1 ));
 AND2_X1 \A1/A1/A2/A2/M2/M2/_0_  (.A1(\A1/A1/A2/A2/M2/s1 ),
    .A2(\A1/A1/A2/A2/c1 ),
    .ZN(\A1/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M2/M2/_1_  (.A(\A1/A1/A2/A2/M2/s1 ),
    .B(\A1/A1/A2/A2/c1 ),
    .Z(s1[13]));
 OR2_X1 \A1/A1/A2/A2/M2/_0_  (.A1(\A1/A1/A2/A2/M2/c1 ),
    .A2(\A1/A1/A2/A2/M2/c2 ),
    .ZN(\A1/A1/A2/A2/c2 ));
 AND2_X1 \A1/A1/A2/A2/M3/M1/_0_  (.A1(v2[14]),
    .A2(v3[14]),
    .ZN(\A1/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M3/M1/_1_  (.A(v2[14]),
    .B(v3[14]),
    .Z(\A1/A1/A2/A2/M3/s1 ));
 AND2_X1 \A1/A1/A2/A2/M3/M2/_0_  (.A1(\A1/A1/A2/A2/M3/s1 ),
    .A2(\A1/A1/A2/A2/c2 ),
    .ZN(\A1/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M3/M2/_1_  (.A(\A1/A1/A2/A2/M3/s1 ),
    .B(\A1/A1/A2/A2/c2 ),
    .Z(s1[14]));
 OR2_X1 \A1/A1/A2/A2/M3/_0_  (.A1(\A1/A1/A2/A2/M3/c1 ),
    .A2(\A1/A1/A2/A2/M3/c2 ),
    .ZN(\A1/A1/A2/A2/c3 ));
 AND2_X1 \A1/A1/A2/A2/M4/M1/_0_  (.A1(v2[15]),
    .A2(v3[15]),
    .ZN(\A1/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M4/M1/_1_  (.A(v2[15]),
    .B(v3[15]),
    .Z(\A1/A1/A2/A2/M4/s1 ));
 AND2_X1 \A1/A1/A2/A2/M4/M2/_0_  (.A1(\A1/A1/A2/A2/M4/s1 ),
    .A2(\A1/A1/A2/A2/c3 ),
    .ZN(\A1/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M4/M2/_1_  (.A(\A1/A1/A2/A2/M4/s1 ),
    .B(\A1/A1/A2/A2/c3 ),
    .Z(s1[15]));
 OR2_X1 \A1/A1/A2/A2/M4/_0_  (.A1(\A1/A1/A2/A2/M4/c1 ),
    .A2(\A1/A1/A2/A2/M4/c2 ),
    .ZN(\A1/c1 ));
 AND2_X1 \A1/A2/A1/A1/M1/M1/_0_  (.A1(v2[16]),
    .A2(v3[16]),
    .ZN(\A1/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M1/M1/_1_  (.A(v2[16]),
    .B(v3[16]),
    .Z(\A1/A2/A1/A1/M1/s1 ));
 AND2_X1 \A1/A2/A1/A1/M1/M2/_0_  (.A1(\A1/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A1/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M1/M2/_1_  (.A(\A1/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(s1[16]));
 OR2_X1 \A1/A2/A1/A1/M1/_0_  (.A1(\A1/A2/A1/A1/M1/c1 ),
    .A2(\A1/A2/A1/A1/M1/c2 ),
    .ZN(\A1/A2/A1/A1/c1 ));
 AND2_X1 \A1/A2/A1/A1/M2/M1/_0_  (.A1(v2[17]),
    .A2(v3[17]),
    .ZN(\A1/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M2/M1/_1_  (.A(v2[17]),
    .B(v3[17]),
    .Z(\A1/A2/A1/A1/M2/s1 ));
 AND2_X1 \A1/A2/A1/A1/M2/M2/_0_  (.A1(\A1/A2/A1/A1/M2/s1 ),
    .A2(\A1/A2/A1/A1/c1 ),
    .ZN(\A1/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M2/M2/_1_  (.A(\A1/A2/A1/A1/M2/s1 ),
    .B(\A1/A2/A1/A1/c1 ),
    .Z(s1[17]));
 OR2_X1 \A1/A2/A1/A1/M2/_0_  (.A1(\A1/A2/A1/A1/M2/c1 ),
    .A2(\A1/A2/A1/A1/M2/c2 ),
    .ZN(\A1/A2/A1/A1/c2 ));
 AND2_X1 \A1/A2/A1/A1/M3/M1/_0_  (.A1(v2[18]),
    .A2(v3[18]),
    .ZN(\A1/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M3/M1/_1_  (.A(v2[18]),
    .B(v3[18]),
    .Z(\A1/A2/A1/A1/M3/s1 ));
 AND2_X1 \A1/A2/A1/A1/M3/M2/_0_  (.A1(\A1/A2/A1/A1/M3/s1 ),
    .A2(\A1/A2/A1/A1/c2 ),
    .ZN(\A1/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M3/M2/_1_  (.A(\A1/A2/A1/A1/M3/s1 ),
    .B(\A1/A2/A1/A1/c2 ),
    .Z(s1[18]));
 OR2_X1 \A1/A2/A1/A1/M3/_0_  (.A1(\A1/A2/A1/A1/M3/c1 ),
    .A2(\A1/A2/A1/A1/M3/c2 ),
    .ZN(\A1/A2/A1/A1/c3 ));
 AND2_X1 \A1/A2/A1/A1/M4/M1/_0_  (.A1(v2[19]),
    .A2(v3[19]),
    .ZN(\A1/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M4/M1/_1_  (.A(v2[19]),
    .B(v3[19]),
    .Z(\A1/A2/A1/A1/M4/s1 ));
 AND2_X1 \A1/A2/A1/A1/M4/M2/_0_  (.A1(\A1/A2/A1/A1/M4/s1 ),
    .A2(\A1/A2/A1/A1/c3 ),
    .ZN(\A1/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M4/M2/_1_  (.A(\A1/A2/A1/A1/M4/s1 ),
    .B(\A1/A2/A1/A1/c3 ),
    .Z(s1[19]));
 OR2_X1 \A1/A2/A1/A1/M4/_0_  (.A1(\A1/A2/A1/A1/M4/c1 ),
    .A2(\A1/A2/A1/A1/M4/c2 ),
    .ZN(\A1/A2/A1/c1 ));
 AND2_X1 \A1/A2/A1/A2/M1/M1/_0_  (.A1(v2[20]),
    .A2(v3[20]),
    .ZN(\A1/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M1/M1/_1_  (.A(v2[20]),
    .B(v3[20]),
    .Z(\A1/A2/A1/A2/M1/s1 ));
 AND2_X1 \A1/A2/A1/A2/M1/M2/_0_  (.A1(\A1/A2/A1/A2/M1/s1 ),
    .A2(\A1/A2/A1/c1 ),
    .ZN(\A1/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M1/M2/_1_  (.A(\A1/A2/A1/A2/M1/s1 ),
    .B(\A1/A2/A1/c1 ),
    .Z(s1[20]));
 OR2_X1 \A1/A2/A1/A2/M1/_0_  (.A1(\A1/A2/A1/A2/M1/c1 ),
    .A2(\A1/A2/A1/A2/M1/c2 ),
    .ZN(\A1/A2/A1/A2/c1 ));
 AND2_X1 \A1/A2/A1/A2/M2/M1/_0_  (.A1(v2[21]),
    .A2(v3[21]),
    .ZN(\A1/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M2/M1/_1_  (.A(v2[21]),
    .B(v3[21]),
    .Z(\A1/A2/A1/A2/M2/s1 ));
 AND2_X1 \A1/A2/A1/A2/M2/M2/_0_  (.A1(\A1/A2/A1/A2/M2/s1 ),
    .A2(\A1/A2/A1/A2/c1 ),
    .ZN(\A1/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M2/M2/_1_  (.A(\A1/A2/A1/A2/M2/s1 ),
    .B(\A1/A2/A1/A2/c1 ),
    .Z(s1[21]));
 OR2_X1 \A1/A2/A1/A2/M2/_0_  (.A1(\A1/A2/A1/A2/M2/c1 ),
    .A2(\A1/A2/A1/A2/M2/c2 ),
    .ZN(\A1/A2/A1/A2/c2 ));
 AND2_X1 \A1/A2/A1/A2/M3/M1/_0_  (.A1(v2[22]),
    .A2(v3[22]),
    .ZN(\A1/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M3/M1/_1_  (.A(v2[22]),
    .B(v3[22]),
    .Z(\A1/A2/A1/A2/M3/s1 ));
 AND2_X1 \A1/A2/A1/A2/M3/M2/_0_  (.A1(\A1/A2/A1/A2/M3/s1 ),
    .A2(\A1/A2/A1/A2/c2 ),
    .ZN(\A1/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M3/M2/_1_  (.A(\A1/A2/A1/A2/M3/s1 ),
    .B(\A1/A2/A1/A2/c2 ),
    .Z(s1[22]));
 OR2_X1 \A1/A2/A1/A2/M3/_0_  (.A1(\A1/A2/A1/A2/M3/c1 ),
    .A2(\A1/A2/A1/A2/M3/c2 ),
    .ZN(\A1/A2/A1/A2/c3 ));
 AND2_X1 \A1/A2/A1/A2/M4/M1/_0_  (.A1(v2[23]),
    .A2(v3[23]),
    .ZN(\A1/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M4/M1/_1_  (.A(v2[23]),
    .B(v3[23]),
    .Z(\A1/A2/A1/A2/M4/s1 ));
 AND2_X1 \A1/A2/A1/A2/M4/M2/_0_  (.A1(\A1/A2/A1/A2/M4/s1 ),
    .A2(\A1/A2/A1/A2/c3 ),
    .ZN(\A1/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M4/M2/_1_  (.A(\A1/A2/A1/A2/M4/s1 ),
    .B(\A1/A2/A1/A2/c3 ),
    .Z(s1[23]));
 OR2_X1 \A1/A2/A1/A2/M4/_0_  (.A1(\A1/A2/A1/A2/M4/c1 ),
    .A2(\A1/A2/A1/A2/M4/c2 ),
    .ZN(\A1/A2/c1 ));
 AND2_X1 \A1/A2/A2/A1/M1/M1/_0_  (.A1(v2[24]),
    .A2(v3[24]),
    .ZN(\A1/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M1/M1/_1_  (.A(v2[24]),
    .B(v3[24]),
    .Z(\A1/A2/A2/A1/M1/s1 ));
 AND2_X1 \A1/A2/A2/A1/M1/M2/_0_  (.A1(\A1/A2/A2/A1/M1/s1 ),
    .A2(\A1/A2/c1 ),
    .ZN(\A1/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M1/M2/_1_  (.A(\A1/A2/A2/A1/M1/s1 ),
    .B(\A1/A2/c1 ),
    .Z(s1[24]));
 OR2_X1 \A1/A2/A2/A1/M1/_0_  (.A1(\A1/A2/A2/A1/M1/c1 ),
    .A2(\A1/A2/A2/A1/M1/c2 ),
    .ZN(\A1/A2/A2/A1/c1 ));
 AND2_X1 \A1/A2/A2/A1/M2/M1/_0_  (.A1(v2[25]),
    .A2(v3[25]),
    .ZN(\A1/A2/A2/A1/M2/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M2/M1/_1_  (.A(v2[25]),
    .B(v3[25]),
    .Z(\A1/A2/A2/A1/M2/s1 ));
 AND2_X1 \A1/A2/A2/A1/M2/M2/_0_  (.A1(\A1/A2/A2/A1/M2/s1 ),
    .A2(\A1/A2/A2/A1/c1 ),
    .ZN(\A1/A2/A2/A1/M2/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M2/M2/_1_  (.A(\A1/A2/A2/A1/M2/s1 ),
    .B(\A1/A2/A2/A1/c1 ),
    .Z(s1[25]));
 OR2_X1 \A1/A2/A2/A1/M2/_0_  (.A1(\A1/A2/A2/A1/M2/c1 ),
    .A2(\A1/A2/A2/A1/M2/c2 ),
    .ZN(\A1/A2/A2/A1/c2 ));
 AND2_X1 \A1/A2/A2/A1/M3/M1/_0_  (.A1(v2[26]),
    .A2(v3[26]),
    .ZN(\A1/A2/A2/A1/M3/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M3/M1/_1_  (.A(v2[26]),
    .B(v3[26]),
    .Z(\A1/A2/A2/A1/M3/s1 ));
 AND2_X1 \A1/A2/A2/A1/M3/M2/_0_  (.A1(\A1/A2/A2/A1/M3/s1 ),
    .A2(\A1/A2/A2/A1/c2 ),
    .ZN(\A1/A2/A2/A1/M3/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M3/M2/_1_  (.A(\A1/A2/A2/A1/M3/s1 ),
    .B(\A1/A2/A2/A1/c2 ),
    .Z(s1[26]));
 OR2_X1 \A1/A2/A2/A1/M3/_0_  (.A1(\A1/A2/A2/A1/M3/c1 ),
    .A2(\A1/A2/A2/A1/M3/c2 ),
    .ZN(\A1/A2/A2/A1/c3 ));
 AND2_X1 \A1/A2/A2/A1/M4/M1/_0_  (.A1(v2[27]),
    .A2(v3[27]),
    .ZN(\A1/A2/A2/A1/M4/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M4/M1/_1_  (.A(v2[27]),
    .B(v3[27]),
    .Z(\A1/A2/A2/A1/M4/s1 ));
 AND2_X1 \A1/A2/A2/A1/M4/M2/_0_  (.A1(\A1/A2/A2/A1/M4/s1 ),
    .A2(\A1/A2/A2/A1/c3 ),
    .ZN(\A1/A2/A2/A1/M4/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M4/M2/_1_  (.A(\A1/A2/A2/A1/M4/s1 ),
    .B(\A1/A2/A2/A1/c3 ),
    .Z(s1[27]));
 OR2_X1 \A1/A2/A2/A1/M4/_0_  (.A1(\A1/A2/A2/A1/M4/c1 ),
    .A2(\A1/A2/A2/A1/M4/c2 ),
    .ZN(\A1/A2/A2/c1 ));
 AND2_X1 \A1/A2/A2/A2/M1/M1/_0_  (.A1(v2[28]),
    .A2(v3[28]),
    .ZN(\A1/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M1/M1/_1_  (.A(v2[28]),
    .B(v3[28]),
    .Z(\A1/A2/A2/A2/M1/s1 ));
 AND2_X1 \A1/A2/A2/A2/M1/M2/_0_  (.A1(\A1/A2/A2/A2/M1/s1 ),
    .A2(\A1/A2/A2/c1 ),
    .ZN(\A1/A2/A2/A2/M1/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M1/M2/_1_  (.A(\A1/A2/A2/A2/M1/s1 ),
    .B(\A1/A2/A2/c1 ),
    .Z(s1[28]));
 OR2_X1 \A1/A2/A2/A2/M1/_0_  (.A1(\A1/A2/A2/A2/M1/c1 ),
    .A2(\A1/A2/A2/A2/M1/c2 ),
    .ZN(\A1/A2/A2/A2/c1 ));
 AND2_X1 \A1/A2/A2/A2/M2/M1/_0_  (.A1(v2[29]),
    .A2(v3[29]),
    .ZN(\A1/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M2/M1/_1_  (.A(v2[29]),
    .B(v3[29]),
    .Z(\A1/A2/A2/A2/M2/s1 ));
 AND2_X1 \A1/A2/A2/A2/M2/M2/_0_  (.A1(\A1/A2/A2/A2/M2/s1 ),
    .A2(\A1/A2/A2/A2/c1 ),
    .ZN(\A1/A2/A2/A2/M2/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M2/M2/_1_  (.A(\A1/A2/A2/A2/M2/s1 ),
    .B(\A1/A2/A2/A2/c1 ),
    .Z(s1[29]));
 OR2_X1 \A1/A2/A2/A2/M2/_0_  (.A1(\A1/A2/A2/A2/M2/c1 ),
    .A2(\A1/A2/A2/A2/M2/c2 ),
    .ZN(\A1/A2/A2/A2/c2 ));
 AND2_X1 \A1/A2/A2/A2/M3/M1/_0_  (.A1(v2[30]),
    .A2(v3[30]),
    .ZN(\A1/A2/A2/A2/M3/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M3/M1/_1_  (.A(v2[30]),
    .B(v3[30]),
    .Z(\A1/A2/A2/A2/M3/s1 ));
 AND2_X1 \A1/A2/A2/A2/M3/M2/_0_  (.A1(\A1/A2/A2/A2/M3/s1 ),
    .A2(\A1/A2/A2/A2/c2 ),
    .ZN(\A1/A2/A2/A2/M3/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M3/M2/_1_  (.A(\A1/A2/A2/A2/M3/s1 ),
    .B(\A1/A2/A2/A2/c2 ),
    .Z(s1[30]));
 OR2_X1 \A1/A2/A2/A2/M3/_0_  (.A1(\A1/A2/A2/A2/M3/c1 ),
    .A2(\A1/A2/A2/A2/M3/c2 ),
    .ZN(\A1/A2/A2/A2/c3 ));
 AND2_X1 \A1/A2/A2/A2/M4/M1/_0_  (.A1(v2[31]),
    .A2(v3[31]),
    .ZN(\A1/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M4/M1/_1_  (.A(v2[31]),
    .B(v3[31]),
    .Z(\A1/A2/A2/A2/M4/s1 ));
 AND2_X1 \A1/A2/A2/A2/M4/M2/_0_  (.A1(\A1/A2/A2/A2/M4/s1 ),
    .A2(\A1/A2/A2/A2/c3 ),
    .ZN(\A1/A2/A2/A2/M4/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M4/M2/_1_  (.A(\A1/A2/A2/A2/M4/s1 ),
    .B(\A1/A2/A2/A2/c3 ),
    .Z(s1[31]));
 OR2_X1 \A1/A2/A2/A2/M4/_0_  (.A1(\A1/A2/A2/A2/M4/c1 ),
    .A2(\A1/A2/A2/A2/M4/c2 ),
    .ZN(c1));
 AND2_X1 \A2/A1/A1/A1/M1/M1/_0_  (.A1(s1[0]),
    .A2(v1[16]),
    .ZN(\A2/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M1/M1/_1_  (.A(s1[0]),
    .B(v1[16]),
    .Z(\A2/A1/A1/A1/M1/s1 ));
 AND2_X1 \A2/A1/A1/A1/M1/M2/_0_  (.A1(\A2/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A2/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M1/M2/_1_  (.A(\A2/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(s2[0]));
 OR2_X1 \A2/A1/A1/A1/M1/_0_  (.A1(\A2/A1/A1/A1/M1/c1 ),
    .A2(\A2/A1/A1/A1/M1/c2 ),
    .ZN(\A2/A1/A1/A1/c1 ));
 AND2_X1 \A2/A1/A1/A1/M2/M1/_0_  (.A1(s1[1]),
    .A2(v1[17]),
    .ZN(\A2/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M2/M1/_1_  (.A(s1[1]),
    .B(v1[17]),
    .Z(\A2/A1/A1/A1/M2/s1 ));
 AND2_X1 \A2/A1/A1/A1/M2/M2/_0_  (.A1(\A2/A1/A1/A1/M2/s1 ),
    .A2(\A2/A1/A1/A1/c1 ),
    .ZN(\A2/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M2/M2/_1_  (.A(\A2/A1/A1/A1/M2/s1 ),
    .B(\A2/A1/A1/A1/c1 ),
    .Z(s2[1]));
 OR2_X1 \A2/A1/A1/A1/M2/_0_  (.A1(\A2/A1/A1/A1/M2/c1 ),
    .A2(\A2/A1/A1/A1/M2/c2 ),
    .ZN(\A2/A1/A1/A1/c2 ));
 AND2_X1 \A2/A1/A1/A1/M3/M1/_0_  (.A1(s1[2]),
    .A2(v1[18]),
    .ZN(\A2/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M3/M1/_1_  (.A(s1[2]),
    .B(v1[18]),
    .Z(\A2/A1/A1/A1/M3/s1 ));
 AND2_X1 \A2/A1/A1/A1/M3/M2/_0_  (.A1(\A2/A1/A1/A1/M3/s1 ),
    .A2(\A2/A1/A1/A1/c2 ),
    .ZN(\A2/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M3/M2/_1_  (.A(\A2/A1/A1/A1/M3/s1 ),
    .B(\A2/A1/A1/A1/c2 ),
    .Z(s2[2]));
 OR2_X1 \A2/A1/A1/A1/M3/_0_  (.A1(\A2/A1/A1/A1/M3/c1 ),
    .A2(\A2/A1/A1/A1/M3/c2 ),
    .ZN(\A2/A1/A1/A1/c3 ));
 AND2_X1 \A2/A1/A1/A1/M4/M1/_0_  (.A1(s1[3]),
    .A2(v1[19]),
    .ZN(\A2/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M4/M1/_1_  (.A(s1[3]),
    .B(v1[19]),
    .Z(\A2/A1/A1/A1/M4/s1 ));
 AND2_X1 \A2/A1/A1/A1/M4/M2/_0_  (.A1(\A2/A1/A1/A1/M4/s1 ),
    .A2(\A2/A1/A1/A1/c3 ),
    .ZN(\A2/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M4/M2/_1_  (.A(\A2/A1/A1/A1/M4/s1 ),
    .B(\A2/A1/A1/A1/c3 ),
    .Z(s2[3]));
 OR2_X1 \A2/A1/A1/A1/M4/_0_  (.A1(\A2/A1/A1/A1/M4/c1 ),
    .A2(\A2/A1/A1/A1/M4/c2 ),
    .ZN(\A2/A1/A1/c1 ));
 AND2_X1 \A2/A1/A1/A2/M1/M1/_0_  (.A1(s1[4]),
    .A2(v1[20]),
    .ZN(\A2/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M1/M1/_1_  (.A(s1[4]),
    .B(v1[20]),
    .Z(\A2/A1/A1/A2/M1/s1 ));
 AND2_X1 \A2/A1/A1/A2/M1/M2/_0_  (.A1(\A2/A1/A1/A2/M1/s1 ),
    .A2(\A2/A1/A1/c1 ),
    .ZN(\A2/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M1/M2/_1_  (.A(\A2/A1/A1/A2/M1/s1 ),
    .B(\A2/A1/A1/c1 ),
    .Z(s2[4]));
 OR2_X1 \A2/A1/A1/A2/M1/_0_  (.A1(\A2/A1/A1/A2/M1/c1 ),
    .A2(\A2/A1/A1/A2/M1/c2 ),
    .ZN(\A2/A1/A1/A2/c1 ));
 AND2_X1 \A2/A1/A1/A2/M2/M1/_0_  (.A1(s1[5]),
    .A2(v1[21]),
    .ZN(\A2/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M2/M1/_1_  (.A(s1[5]),
    .B(v1[21]),
    .Z(\A2/A1/A1/A2/M2/s1 ));
 AND2_X1 \A2/A1/A1/A2/M2/M2/_0_  (.A1(\A2/A1/A1/A2/M2/s1 ),
    .A2(\A2/A1/A1/A2/c1 ),
    .ZN(\A2/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M2/M2/_1_  (.A(\A2/A1/A1/A2/M2/s1 ),
    .B(\A2/A1/A1/A2/c1 ),
    .Z(s2[5]));
 OR2_X1 \A2/A1/A1/A2/M2/_0_  (.A1(\A2/A1/A1/A2/M2/c1 ),
    .A2(\A2/A1/A1/A2/M2/c2 ),
    .ZN(\A2/A1/A1/A2/c2 ));
 AND2_X1 \A2/A1/A1/A2/M3/M1/_0_  (.A1(s1[6]),
    .A2(v1[22]),
    .ZN(\A2/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M3/M1/_1_  (.A(s1[6]),
    .B(v1[22]),
    .Z(\A2/A1/A1/A2/M3/s1 ));
 AND2_X1 \A2/A1/A1/A2/M3/M2/_0_  (.A1(\A2/A1/A1/A2/M3/s1 ),
    .A2(\A2/A1/A1/A2/c2 ),
    .ZN(\A2/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M3/M2/_1_  (.A(\A2/A1/A1/A2/M3/s1 ),
    .B(\A2/A1/A1/A2/c2 ),
    .Z(s2[6]));
 OR2_X1 \A2/A1/A1/A2/M3/_0_  (.A1(\A2/A1/A1/A2/M3/c1 ),
    .A2(\A2/A1/A1/A2/M3/c2 ),
    .ZN(\A2/A1/A1/A2/c3 ));
 AND2_X1 \A2/A1/A1/A2/M4/M1/_0_  (.A1(s1[7]),
    .A2(v1[23]),
    .ZN(\A2/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M4/M1/_1_  (.A(s1[7]),
    .B(v1[23]),
    .Z(\A2/A1/A1/A2/M4/s1 ));
 AND2_X1 \A2/A1/A1/A2/M4/M2/_0_  (.A1(\A2/A1/A1/A2/M4/s1 ),
    .A2(\A2/A1/A1/A2/c3 ),
    .ZN(\A2/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M4/M2/_1_  (.A(\A2/A1/A1/A2/M4/s1 ),
    .B(\A2/A1/A1/A2/c3 ),
    .Z(s2[7]));
 OR2_X1 \A2/A1/A1/A2/M4/_0_  (.A1(\A2/A1/A1/A2/M4/c1 ),
    .A2(\A2/A1/A1/A2/M4/c2 ),
    .ZN(\A2/A1/c1 ));
 AND2_X1 \A2/A1/A2/A1/M1/M1/_0_  (.A1(s1[8]),
    .A2(v1[24]),
    .ZN(\A2/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M1/M1/_1_  (.A(s1[8]),
    .B(v1[24]),
    .Z(\A2/A1/A2/A1/M1/s1 ));
 AND2_X1 \A2/A1/A2/A1/M1/M2/_0_  (.A1(\A2/A1/A2/A1/M1/s1 ),
    .A2(\A2/A1/c1 ),
    .ZN(\A2/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M1/M2/_1_  (.A(\A2/A1/A2/A1/M1/s1 ),
    .B(\A2/A1/c1 ),
    .Z(s2[8]));
 OR2_X1 \A2/A1/A2/A1/M1/_0_  (.A1(\A2/A1/A2/A1/M1/c1 ),
    .A2(\A2/A1/A2/A1/M1/c2 ),
    .ZN(\A2/A1/A2/A1/c1 ));
 AND2_X1 \A2/A1/A2/A1/M2/M1/_0_  (.A1(s1[9]),
    .A2(v1[25]),
    .ZN(\A2/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M2/M1/_1_  (.A(s1[9]),
    .B(v1[25]),
    .Z(\A2/A1/A2/A1/M2/s1 ));
 AND2_X1 \A2/A1/A2/A1/M2/M2/_0_  (.A1(\A2/A1/A2/A1/M2/s1 ),
    .A2(\A2/A1/A2/A1/c1 ),
    .ZN(\A2/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M2/M2/_1_  (.A(\A2/A1/A2/A1/M2/s1 ),
    .B(\A2/A1/A2/A1/c1 ),
    .Z(s2[9]));
 OR2_X1 \A2/A1/A2/A1/M2/_0_  (.A1(\A2/A1/A2/A1/M2/c1 ),
    .A2(\A2/A1/A2/A1/M2/c2 ),
    .ZN(\A2/A1/A2/A1/c2 ));
 AND2_X1 \A2/A1/A2/A1/M3/M1/_0_  (.A1(s1[10]),
    .A2(v1[26]),
    .ZN(\A2/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M3/M1/_1_  (.A(s1[10]),
    .B(v1[26]),
    .Z(\A2/A1/A2/A1/M3/s1 ));
 AND2_X1 \A2/A1/A2/A1/M3/M2/_0_  (.A1(\A2/A1/A2/A1/M3/s1 ),
    .A2(\A2/A1/A2/A1/c2 ),
    .ZN(\A2/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M3/M2/_1_  (.A(\A2/A1/A2/A1/M3/s1 ),
    .B(\A2/A1/A2/A1/c2 ),
    .Z(s2[10]));
 OR2_X1 \A2/A1/A2/A1/M3/_0_  (.A1(\A2/A1/A2/A1/M3/c1 ),
    .A2(\A2/A1/A2/A1/M3/c2 ),
    .ZN(\A2/A1/A2/A1/c3 ));
 AND2_X1 \A2/A1/A2/A1/M4/M1/_0_  (.A1(s1[11]),
    .A2(v1[27]),
    .ZN(\A2/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M4/M1/_1_  (.A(s1[11]),
    .B(v1[27]),
    .Z(\A2/A1/A2/A1/M4/s1 ));
 AND2_X1 \A2/A1/A2/A1/M4/M2/_0_  (.A1(\A2/A1/A2/A1/M4/s1 ),
    .A2(\A2/A1/A2/A1/c3 ),
    .ZN(\A2/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M4/M2/_1_  (.A(\A2/A1/A2/A1/M4/s1 ),
    .B(\A2/A1/A2/A1/c3 ),
    .Z(s2[11]));
 OR2_X1 \A2/A1/A2/A1/M4/_0_  (.A1(\A2/A1/A2/A1/M4/c1 ),
    .A2(\A2/A1/A2/A1/M4/c2 ),
    .ZN(\A2/A1/A2/c1 ));
 AND2_X1 \A2/A1/A2/A2/M1/M1/_0_  (.A1(s1[12]),
    .A2(v1[28]),
    .ZN(\A2/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M1/M1/_1_  (.A(s1[12]),
    .B(v1[28]),
    .Z(\A2/A1/A2/A2/M1/s1 ));
 AND2_X1 \A2/A1/A2/A2/M1/M2/_0_  (.A1(\A2/A1/A2/A2/M1/s1 ),
    .A2(\A2/A1/A2/c1 ),
    .ZN(\A2/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M1/M2/_1_  (.A(\A2/A1/A2/A2/M1/s1 ),
    .B(\A2/A1/A2/c1 ),
    .Z(s2[12]));
 OR2_X1 \A2/A1/A2/A2/M1/_0_  (.A1(\A2/A1/A2/A2/M1/c1 ),
    .A2(\A2/A1/A2/A2/M1/c2 ),
    .ZN(\A2/A1/A2/A2/c1 ));
 AND2_X1 \A2/A1/A2/A2/M2/M1/_0_  (.A1(s1[13]),
    .A2(v1[29]),
    .ZN(\A2/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M2/M1/_1_  (.A(s1[13]),
    .B(v1[29]),
    .Z(\A2/A1/A2/A2/M2/s1 ));
 AND2_X1 \A2/A1/A2/A2/M2/M2/_0_  (.A1(\A2/A1/A2/A2/M2/s1 ),
    .A2(\A2/A1/A2/A2/c1 ),
    .ZN(\A2/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M2/M2/_1_  (.A(\A2/A1/A2/A2/M2/s1 ),
    .B(\A2/A1/A2/A2/c1 ),
    .Z(s2[13]));
 OR2_X1 \A2/A1/A2/A2/M2/_0_  (.A1(\A2/A1/A2/A2/M2/c1 ),
    .A2(\A2/A1/A2/A2/M2/c2 ),
    .ZN(\A2/A1/A2/A2/c2 ));
 AND2_X1 \A2/A1/A2/A2/M3/M1/_0_  (.A1(s1[14]),
    .A2(v1[30]),
    .ZN(\A2/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M3/M1/_1_  (.A(s1[14]),
    .B(v1[30]),
    .Z(\A2/A1/A2/A2/M3/s1 ));
 AND2_X1 \A2/A1/A2/A2/M3/M2/_0_  (.A1(\A2/A1/A2/A2/M3/s1 ),
    .A2(\A2/A1/A2/A2/c2 ),
    .ZN(\A2/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M3/M2/_1_  (.A(\A2/A1/A2/A2/M3/s1 ),
    .B(\A2/A1/A2/A2/c2 ),
    .Z(s2[14]));
 OR2_X1 \A2/A1/A2/A2/M3/_0_  (.A1(\A2/A1/A2/A2/M3/c1 ),
    .A2(\A2/A1/A2/A2/M3/c2 ),
    .ZN(\A2/A1/A2/A2/c3 ));
 AND2_X1 \A2/A1/A2/A2/M4/M1/_0_  (.A1(s1[15]),
    .A2(v1[31]),
    .ZN(\A2/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M4/M1/_1_  (.A(s1[15]),
    .B(v1[31]),
    .Z(\A2/A1/A2/A2/M4/s1 ));
 AND2_X1 \A2/A1/A2/A2/M4/M2/_0_  (.A1(\A2/A1/A2/A2/M4/s1 ),
    .A2(\A2/A1/A2/A2/c3 ),
    .ZN(\A2/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M4/M2/_1_  (.A(\A2/A1/A2/A2/M4/s1 ),
    .B(\A2/A1/A2/A2/c3 ),
    .Z(s2[15]));
 OR2_X1 \A2/A1/A2/A2/M4/_0_  (.A1(\A2/A1/A2/A2/M4/c1 ),
    .A2(\A2/A1/A2/A2/M4/c2 ),
    .ZN(\A2/c1 ));
 AND2_X1 \A2/A2/A1/A1/M1/M1/_0_  (.A1(s1[16]),
    .A2(ground),
    .ZN(\A2/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M1/M1/_1_  (.A(s1[16]),
    .B(ground),
    .Z(\A2/A2/A1/A1/M1/s1 ));
 AND2_X1 \A2/A2/A1/A1/M1/M2/_0_  (.A1(\A2/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A2/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M1/M2/_1_  (.A(\A2/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(s2[16]));
 OR2_X1 \A2/A2/A1/A1/M1/_0_  (.A1(\A2/A2/A1/A1/M1/c1 ),
    .A2(\A2/A2/A1/A1/M1/c2 ),
    .ZN(\A2/A2/A1/A1/c1 ));
 AND2_X1 \A2/A2/A1/A1/M2/M1/_0_  (.A1(s1[17]),
    .A2(ground),
    .ZN(\A2/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M2/M1/_1_  (.A(s1[17]),
    .B(ground),
    .Z(\A2/A2/A1/A1/M2/s1 ));
 AND2_X1 \A2/A2/A1/A1/M2/M2/_0_  (.A1(\A2/A2/A1/A1/M2/s1 ),
    .A2(\A2/A2/A1/A1/c1 ),
    .ZN(\A2/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M2/M2/_1_  (.A(\A2/A2/A1/A1/M2/s1 ),
    .B(\A2/A2/A1/A1/c1 ),
    .Z(s2[17]));
 OR2_X1 \A2/A2/A1/A1/M2/_0_  (.A1(\A2/A2/A1/A1/M2/c1 ),
    .A2(\A2/A2/A1/A1/M2/c2 ),
    .ZN(\A2/A2/A1/A1/c2 ));
 AND2_X1 \A2/A2/A1/A1/M3/M1/_0_  (.A1(s1[18]),
    .A2(ground),
    .ZN(\A2/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M3/M1/_1_  (.A(s1[18]),
    .B(ground),
    .Z(\A2/A2/A1/A1/M3/s1 ));
 AND2_X1 \A2/A2/A1/A1/M3/M2/_0_  (.A1(\A2/A2/A1/A1/M3/s1 ),
    .A2(\A2/A2/A1/A1/c2 ),
    .ZN(\A2/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M3/M2/_1_  (.A(\A2/A2/A1/A1/M3/s1 ),
    .B(\A2/A2/A1/A1/c2 ),
    .Z(s2[18]));
 OR2_X1 \A2/A2/A1/A1/M3/_0_  (.A1(\A2/A2/A1/A1/M3/c1 ),
    .A2(\A2/A2/A1/A1/M3/c2 ),
    .ZN(\A2/A2/A1/A1/c3 ));
 AND2_X1 \A2/A2/A1/A1/M4/M1/_0_  (.A1(s1[19]),
    .A2(ground),
    .ZN(\A2/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M4/M1/_1_  (.A(s1[19]),
    .B(ground),
    .Z(\A2/A2/A1/A1/M4/s1 ));
 AND2_X1 \A2/A2/A1/A1/M4/M2/_0_  (.A1(\A2/A2/A1/A1/M4/s1 ),
    .A2(\A2/A2/A1/A1/c3 ),
    .ZN(\A2/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M4/M2/_1_  (.A(\A2/A2/A1/A1/M4/s1 ),
    .B(\A2/A2/A1/A1/c3 ),
    .Z(s2[19]));
 OR2_X1 \A2/A2/A1/A1/M4/_0_  (.A1(\A2/A2/A1/A1/M4/c1 ),
    .A2(\A2/A2/A1/A1/M4/c2 ),
    .ZN(\A2/A2/A1/c1 ));
 AND2_X1 \A2/A2/A1/A2/M1/M1/_0_  (.A1(s1[20]),
    .A2(ground),
    .ZN(\A2/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M1/M1/_1_  (.A(s1[20]),
    .B(ground),
    .Z(\A2/A2/A1/A2/M1/s1 ));
 AND2_X1 \A2/A2/A1/A2/M1/M2/_0_  (.A1(\A2/A2/A1/A2/M1/s1 ),
    .A2(\A2/A2/A1/c1 ),
    .ZN(\A2/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M1/M2/_1_  (.A(\A2/A2/A1/A2/M1/s1 ),
    .B(\A2/A2/A1/c1 ),
    .Z(s2[20]));
 OR2_X1 \A2/A2/A1/A2/M1/_0_  (.A1(\A2/A2/A1/A2/M1/c1 ),
    .A2(\A2/A2/A1/A2/M1/c2 ),
    .ZN(\A2/A2/A1/A2/c1 ));
 AND2_X1 \A2/A2/A1/A2/M2/M1/_0_  (.A1(s1[21]),
    .A2(ground),
    .ZN(\A2/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M2/M1/_1_  (.A(s1[21]),
    .B(ground),
    .Z(\A2/A2/A1/A2/M2/s1 ));
 AND2_X1 \A2/A2/A1/A2/M2/M2/_0_  (.A1(\A2/A2/A1/A2/M2/s1 ),
    .A2(\A2/A2/A1/A2/c1 ),
    .ZN(\A2/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M2/M2/_1_  (.A(\A2/A2/A1/A2/M2/s1 ),
    .B(\A2/A2/A1/A2/c1 ),
    .Z(s2[21]));
 OR2_X1 \A2/A2/A1/A2/M2/_0_  (.A1(\A2/A2/A1/A2/M2/c1 ),
    .A2(\A2/A2/A1/A2/M2/c2 ),
    .ZN(\A2/A2/A1/A2/c2 ));
 AND2_X1 \A2/A2/A1/A2/M3/M1/_0_  (.A1(s1[22]),
    .A2(ground),
    .ZN(\A2/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M3/M1/_1_  (.A(s1[22]),
    .B(ground),
    .Z(\A2/A2/A1/A2/M3/s1 ));
 AND2_X1 \A2/A2/A1/A2/M3/M2/_0_  (.A1(\A2/A2/A1/A2/M3/s1 ),
    .A2(\A2/A2/A1/A2/c2 ),
    .ZN(\A2/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M3/M2/_1_  (.A(\A2/A2/A1/A2/M3/s1 ),
    .B(\A2/A2/A1/A2/c2 ),
    .Z(s2[22]));
 OR2_X1 \A2/A2/A1/A2/M3/_0_  (.A1(\A2/A2/A1/A2/M3/c1 ),
    .A2(\A2/A2/A1/A2/M3/c2 ),
    .ZN(\A2/A2/A1/A2/c3 ));
 AND2_X1 \A2/A2/A1/A2/M4/M1/_0_  (.A1(s1[23]),
    .A2(ground),
    .ZN(\A2/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M4/M1/_1_  (.A(s1[23]),
    .B(ground),
    .Z(\A2/A2/A1/A2/M4/s1 ));
 AND2_X1 \A2/A2/A1/A2/M4/M2/_0_  (.A1(\A2/A2/A1/A2/M4/s1 ),
    .A2(\A2/A2/A1/A2/c3 ),
    .ZN(\A2/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M4/M2/_1_  (.A(\A2/A2/A1/A2/M4/s1 ),
    .B(\A2/A2/A1/A2/c3 ),
    .Z(s2[23]));
 OR2_X1 \A2/A2/A1/A2/M4/_0_  (.A1(\A2/A2/A1/A2/M4/c1 ),
    .A2(\A2/A2/A1/A2/M4/c2 ),
    .ZN(\A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A1/M1/M1/_0_  (.A1(s1[24]),
    .A2(ground),
    .ZN(\A2/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M1/M1/_1_  (.A(s1[24]),
    .B(ground),
    .Z(\A2/A2/A2/A1/M1/s1 ));
 AND2_X1 \A2/A2/A2/A1/M1/M2/_0_  (.A1(\A2/A2/A2/A1/M1/s1 ),
    .A2(\A2/A2/c1 ),
    .ZN(\A2/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M1/M2/_1_  (.A(\A2/A2/A2/A1/M1/s1 ),
    .B(\A2/A2/c1 ),
    .Z(s2[24]));
 OR2_X1 \A2/A2/A2/A1/M1/_0_  (.A1(\A2/A2/A2/A1/M1/c1 ),
    .A2(\A2/A2/A2/A1/M1/c2 ),
    .ZN(\A2/A2/A2/A1/c1 ));
 AND2_X1 \A2/A2/A2/A1/M2/M1/_0_  (.A1(s1[25]),
    .A2(ground),
    .ZN(\A2/A2/A2/A1/M2/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M2/M1/_1_  (.A(s1[25]),
    .B(ground),
    .Z(\A2/A2/A2/A1/M2/s1 ));
 AND2_X1 \A2/A2/A2/A1/M2/M2/_0_  (.A1(\A2/A2/A2/A1/M2/s1 ),
    .A2(\A2/A2/A2/A1/c1 ),
    .ZN(\A2/A2/A2/A1/M2/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M2/M2/_1_  (.A(\A2/A2/A2/A1/M2/s1 ),
    .B(\A2/A2/A2/A1/c1 ),
    .Z(s2[25]));
 OR2_X1 \A2/A2/A2/A1/M2/_0_  (.A1(\A2/A2/A2/A1/M2/c1 ),
    .A2(\A2/A2/A2/A1/M2/c2 ),
    .ZN(\A2/A2/A2/A1/c2 ));
 AND2_X1 \A2/A2/A2/A1/M3/M1/_0_  (.A1(s1[26]),
    .A2(ground),
    .ZN(\A2/A2/A2/A1/M3/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M3/M1/_1_  (.A(s1[26]),
    .B(ground),
    .Z(\A2/A2/A2/A1/M3/s1 ));
 AND2_X1 \A2/A2/A2/A1/M3/M2/_0_  (.A1(\A2/A2/A2/A1/M3/s1 ),
    .A2(\A2/A2/A2/A1/c2 ),
    .ZN(\A2/A2/A2/A1/M3/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M3/M2/_1_  (.A(\A2/A2/A2/A1/M3/s1 ),
    .B(\A2/A2/A2/A1/c2 ),
    .Z(s2[26]));
 OR2_X1 \A2/A2/A2/A1/M3/_0_  (.A1(\A2/A2/A2/A1/M3/c1 ),
    .A2(\A2/A2/A2/A1/M3/c2 ),
    .ZN(\A2/A2/A2/A1/c3 ));
 AND2_X1 \A2/A2/A2/A1/M4/M1/_0_  (.A1(s1[27]),
    .A2(ground),
    .ZN(\A2/A2/A2/A1/M4/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M4/M1/_1_  (.A(s1[27]),
    .B(ground),
    .Z(\A2/A2/A2/A1/M4/s1 ));
 AND2_X1 \A2/A2/A2/A1/M4/M2/_0_  (.A1(\A2/A2/A2/A1/M4/s1 ),
    .A2(\A2/A2/A2/A1/c3 ),
    .ZN(\A2/A2/A2/A1/M4/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M4/M2/_1_  (.A(\A2/A2/A2/A1/M4/s1 ),
    .B(\A2/A2/A2/A1/c3 ),
    .Z(s2[27]));
 OR2_X1 \A2/A2/A2/A1/M4/_0_  (.A1(\A2/A2/A2/A1/M4/c1 ),
    .A2(\A2/A2/A2/A1/M4/c2 ),
    .ZN(\A2/A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A2/M1/M1/_0_  (.A1(s1[28]),
    .A2(ground),
    .ZN(\A2/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M1/M1/_1_  (.A(s1[28]),
    .B(ground),
    .Z(\A2/A2/A2/A2/M1/s1 ));
 AND2_X1 \A2/A2/A2/A2/M1/M2/_0_  (.A1(\A2/A2/A2/A2/M1/s1 ),
    .A2(\A2/A2/A2/c1 ),
    .ZN(\A2/A2/A2/A2/M1/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M1/M2/_1_  (.A(\A2/A2/A2/A2/M1/s1 ),
    .B(\A2/A2/A2/c1 ),
    .Z(s2[28]));
 OR2_X1 \A2/A2/A2/A2/M1/_0_  (.A1(\A2/A2/A2/A2/M1/c1 ),
    .A2(\A2/A2/A2/A2/M1/c2 ),
    .ZN(\A2/A2/A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A2/M2/M1/_0_  (.A1(s1[29]),
    .A2(ground),
    .ZN(\A2/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M2/M1/_1_  (.A(s1[29]),
    .B(ground),
    .Z(\A2/A2/A2/A2/M2/s1 ));
 AND2_X1 \A2/A2/A2/A2/M2/M2/_0_  (.A1(\A2/A2/A2/A2/M2/s1 ),
    .A2(\A2/A2/A2/A2/c1 ),
    .ZN(\A2/A2/A2/A2/M2/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M2/M2/_1_  (.A(\A2/A2/A2/A2/M2/s1 ),
    .B(\A2/A2/A2/A2/c1 ),
    .Z(s2[29]));
 OR2_X1 \A2/A2/A2/A2/M2/_0_  (.A1(\A2/A2/A2/A2/M2/c1 ),
    .A2(\A2/A2/A2/A2/M2/c2 ),
    .ZN(\A2/A2/A2/A2/c2 ));
 AND2_X1 \A2/A2/A2/A2/M3/M1/_0_  (.A1(s1[30]),
    .A2(ground),
    .ZN(\A2/A2/A2/A2/M3/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M3/M1/_1_  (.A(s1[30]),
    .B(ground),
    .Z(\A2/A2/A2/A2/M3/s1 ));
 AND2_X1 \A2/A2/A2/A2/M3/M2/_0_  (.A1(\A2/A2/A2/A2/M3/s1 ),
    .A2(\A2/A2/A2/A2/c2 ),
    .ZN(\A2/A2/A2/A2/M3/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M3/M2/_1_  (.A(\A2/A2/A2/A2/M3/s1 ),
    .B(\A2/A2/A2/A2/c2 ),
    .Z(s2[30]));
 OR2_X1 \A2/A2/A2/A2/M3/_0_  (.A1(\A2/A2/A2/A2/M3/c1 ),
    .A2(\A2/A2/A2/A2/M3/c2 ),
    .ZN(\A2/A2/A2/A2/c3 ));
 AND2_X1 \A2/A2/A2/A2/M4/M1/_0_  (.A1(s1[31]),
    .A2(ground),
    .ZN(\A2/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M4/M1/_1_  (.A(s1[31]),
    .B(ground),
    .Z(\A2/A2/A2/A2/M4/s1 ));
 AND2_X1 \A2/A2/A2/A2/M4/M2/_0_  (.A1(\A2/A2/A2/A2/M4/s1 ),
    .A2(\A2/A2/A2/A2/c3 ),
    .ZN(\A2/A2/A2/A2/M4/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M4/M2/_1_  (.A(\A2/A2/A2/A2/M4/s1 ),
    .B(\A2/A2/A2/A2/c3 ),
    .Z(s2[31]));
 OR2_X1 \A2/A2/A2/A2/M4/_0_  (.A1(\A2/A2/A2/A2/M4/c1 ),
    .A2(\A2/A2/A2/A2/M4/c2 ),
    .ZN(c2));
 AND2_X1 \A3/A1/A1/A1/M1/M1/_0_  (.A1(v4[0]),
    .A2(s2[16]),
    .ZN(\A3/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M1/M1/_1_  (.A(v4[0]),
    .B(s2[16]),
    .Z(\A3/A1/A1/A1/M1/s1 ));
 AND2_X1 \A3/A1/A1/A1/M1/M2/_0_  (.A1(\A3/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A3/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M1/M2/_1_  (.A(\A3/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(Prod[32]));
 OR2_X1 \A3/A1/A1/A1/M1/_0_  (.A1(\A3/A1/A1/A1/M1/c1 ),
    .A2(\A3/A1/A1/A1/M1/c2 ),
    .ZN(\A3/A1/A1/A1/c1 ));
 AND2_X1 \A3/A1/A1/A1/M2/M1/_0_  (.A1(v4[1]),
    .A2(s2[17]),
    .ZN(\A3/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M2/M1/_1_  (.A(v4[1]),
    .B(s2[17]),
    .Z(\A3/A1/A1/A1/M2/s1 ));
 AND2_X1 \A3/A1/A1/A1/M2/M2/_0_  (.A1(\A3/A1/A1/A1/M2/s1 ),
    .A2(\A3/A1/A1/A1/c1 ),
    .ZN(\A3/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M2/M2/_1_  (.A(\A3/A1/A1/A1/M2/s1 ),
    .B(\A3/A1/A1/A1/c1 ),
    .Z(Prod[33]));
 OR2_X1 \A3/A1/A1/A1/M2/_0_  (.A1(\A3/A1/A1/A1/M2/c1 ),
    .A2(\A3/A1/A1/A1/M2/c2 ),
    .ZN(\A3/A1/A1/A1/c2 ));
 AND2_X1 \A3/A1/A1/A1/M3/M1/_0_  (.A1(v4[2]),
    .A2(s2[18]),
    .ZN(\A3/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M3/M1/_1_  (.A(v4[2]),
    .B(s2[18]),
    .Z(\A3/A1/A1/A1/M3/s1 ));
 AND2_X1 \A3/A1/A1/A1/M3/M2/_0_  (.A1(\A3/A1/A1/A1/M3/s1 ),
    .A2(\A3/A1/A1/A1/c2 ),
    .ZN(\A3/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M3/M2/_1_  (.A(\A3/A1/A1/A1/M3/s1 ),
    .B(\A3/A1/A1/A1/c2 ),
    .Z(Prod[34]));
 OR2_X1 \A3/A1/A1/A1/M3/_0_  (.A1(\A3/A1/A1/A1/M3/c1 ),
    .A2(\A3/A1/A1/A1/M3/c2 ),
    .ZN(\A3/A1/A1/A1/c3 ));
 AND2_X1 \A3/A1/A1/A1/M4/M1/_0_  (.A1(v4[3]),
    .A2(s2[19]),
    .ZN(\A3/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M4/M1/_1_  (.A(v4[3]),
    .B(s2[19]),
    .Z(\A3/A1/A1/A1/M4/s1 ));
 AND2_X1 \A3/A1/A1/A1/M4/M2/_0_  (.A1(\A3/A1/A1/A1/M4/s1 ),
    .A2(\A3/A1/A1/A1/c3 ),
    .ZN(\A3/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M4/M2/_1_  (.A(\A3/A1/A1/A1/M4/s1 ),
    .B(\A3/A1/A1/A1/c3 ),
    .Z(Prod[35]));
 OR2_X1 \A3/A1/A1/A1/M4/_0_  (.A1(\A3/A1/A1/A1/M4/c1 ),
    .A2(\A3/A1/A1/A1/M4/c2 ),
    .ZN(\A3/A1/A1/c1 ));
 AND2_X1 \A3/A1/A1/A2/M1/M1/_0_  (.A1(v4[4]),
    .A2(s2[20]),
    .ZN(\A3/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M1/M1/_1_  (.A(v4[4]),
    .B(s2[20]),
    .Z(\A3/A1/A1/A2/M1/s1 ));
 AND2_X1 \A3/A1/A1/A2/M1/M2/_0_  (.A1(\A3/A1/A1/A2/M1/s1 ),
    .A2(\A3/A1/A1/c1 ),
    .ZN(\A3/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M1/M2/_1_  (.A(\A3/A1/A1/A2/M1/s1 ),
    .B(\A3/A1/A1/c1 ),
    .Z(Prod[36]));
 OR2_X1 \A3/A1/A1/A2/M1/_0_  (.A1(\A3/A1/A1/A2/M1/c1 ),
    .A2(\A3/A1/A1/A2/M1/c2 ),
    .ZN(\A3/A1/A1/A2/c1 ));
 AND2_X1 \A3/A1/A1/A2/M2/M1/_0_  (.A1(v4[5]),
    .A2(s2[21]),
    .ZN(\A3/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M2/M1/_1_  (.A(v4[5]),
    .B(s2[21]),
    .Z(\A3/A1/A1/A2/M2/s1 ));
 AND2_X1 \A3/A1/A1/A2/M2/M2/_0_  (.A1(\A3/A1/A1/A2/M2/s1 ),
    .A2(\A3/A1/A1/A2/c1 ),
    .ZN(\A3/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M2/M2/_1_  (.A(\A3/A1/A1/A2/M2/s1 ),
    .B(\A3/A1/A1/A2/c1 ),
    .Z(Prod[37]));
 OR2_X1 \A3/A1/A1/A2/M2/_0_  (.A1(\A3/A1/A1/A2/M2/c1 ),
    .A2(\A3/A1/A1/A2/M2/c2 ),
    .ZN(\A3/A1/A1/A2/c2 ));
 AND2_X1 \A3/A1/A1/A2/M3/M1/_0_  (.A1(v4[6]),
    .A2(s2[22]),
    .ZN(\A3/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M3/M1/_1_  (.A(v4[6]),
    .B(s2[22]),
    .Z(\A3/A1/A1/A2/M3/s1 ));
 AND2_X1 \A3/A1/A1/A2/M3/M2/_0_  (.A1(\A3/A1/A1/A2/M3/s1 ),
    .A2(\A3/A1/A1/A2/c2 ),
    .ZN(\A3/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M3/M2/_1_  (.A(\A3/A1/A1/A2/M3/s1 ),
    .B(\A3/A1/A1/A2/c2 ),
    .Z(Prod[38]));
 OR2_X1 \A3/A1/A1/A2/M3/_0_  (.A1(\A3/A1/A1/A2/M3/c1 ),
    .A2(\A3/A1/A1/A2/M3/c2 ),
    .ZN(\A3/A1/A1/A2/c3 ));
 AND2_X1 \A3/A1/A1/A2/M4/M1/_0_  (.A1(v4[7]),
    .A2(s2[23]),
    .ZN(\A3/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M4/M1/_1_  (.A(v4[7]),
    .B(s2[23]),
    .Z(\A3/A1/A1/A2/M4/s1 ));
 AND2_X1 \A3/A1/A1/A2/M4/M2/_0_  (.A1(\A3/A1/A1/A2/M4/s1 ),
    .A2(\A3/A1/A1/A2/c3 ),
    .ZN(\A3/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M4/M2/_1_  (.A(\A3/A1/A1/A2/M4/s1 ),
    .B(\A3/A1/A1/A2/c3 ),
    .Z(Prod[39]));
 OR2_X1 \A3/A1/A1/A2/M4/_0_  (.A1(\A3/A1/A1/A2/M4/c1 ),
    .A2(\A3/A1/A1/A2/M4/c2 ),
    .ZN(\A3/A1/c1 ));
 AND2_X1 \A3/A1/A2/A1/M1/M1/_0_  (.A1(v4[8]),
    .A2(s2[24]),
    .ZN(\A3/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M1/M1/_1_  (.A(v4[8]),
    .B(s2[24]),
    .Z(\A3/A1/A2/A1/M1/s1 ));
 AND2_X1 \A3/A1/A2/A1/M1/M2/_0_  (.A1(\A3/A1/A2/A1/M1/s1 ),
    .A2(\A3/A1/c1 ),
    .ZN(\A3/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M1/M2/_1_  (.A(\A3/A1/A2/A1/M1/s1 ),
    .B(\A3/A1/c1 ),
    .Z(Prod[40]));
 OR2_X1 \A3/A1/A2/A1/M1/_0_  (.A1(\A3/A1/A2/A1/M1/c1 ),
    .A2(\A3/A1/A2/A1/M1/c2 ),
    .ZN(\A3/A1/A2/A1/c1 ));
 AND2_X1 \A3/A1/A2/A1/M2/M1/_0_  (.A1(v4[9]),
    .A2(s2[25]),
    .ZN(\A3/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M2/M1/_1_  (.A(v4[9]),
    .B(s2[25]),
    .Z(\A3/A1/A2/A1/M2/s1 ));
 AND2_X1 \A3/A1/A2/A1/M2/M2/_0_  (.A1(\A3/A1/A2/A1/M2/s1 ),
    .A2(\A3/A1/A2/A1/c1 ),
    .ZN(\A3/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M2/M2/_1_  (.A(\A3/A1/A2/A1/M2/s1 ),
    .B(\A3/A1/A2/A1/c1 ),
    .Z(Prod[41]));
 OR2_X1 \A3/A1/A2/A1/M2/_0_  (.A1(\A3/A1/A2/A1/M2/c1 ),
    .A2(\A3/A1/A2/A1/M2/c2 ),
    .ZN(\A3/A1/A2/A1/c2 ));
 AND2_X1 \A3/A1/A2/A1/M3/M1/_0_  (.A1(v4[10]),
    .A2(s2[26]),
    .ZN(\A3/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M3/M1/_1_  (.A(v4[10]),
    .B(s2[26]),
    .Z(\A3/A1/A2/A1/M3/s1 ));
 AND2_X1 \A3/A1/A2/A1/M3/M2/_0_  (.A1(\A3/A1/A2/A1/M3/s1 ),
    .A2(\A3/A1/A2/A1/c2 ),
    .ZN(\A3/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M3/M2/_1_  (.A(\A3/A1/A2/A1/M3/s1 ),
    .B(\A3/A1/A2/A1/c2 ),
    .Z(Prod[42]));
 OR2_X1 \A3/A1/A2/A1/M3/_0_  (.A1(\A3/A1/A2/A1/M3/c1 ),
    .A2(\A3/A1/A2/A1/M3/c2 ),
    .ZN(\A3/A1/A2/A1/c3 ));
 AND2_X1 \A3/A1/A2/A1/M4/M1/_0_  (.A1(v4[11]),
    .A2(s2[27]),
    .ZN(\A3/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M4/M1/_1_  (.A(v4[11]),
    .B(s2[27]),
    .Z(\A3/A1/A2/A1/M4/s1 ));
 AND2_X1 \A3/A1/A2/A1/M4/M2/_0_  (.A1(\A3/A1/A2/A1/M4/s1 ),
    .A2(\A3/A1/A2/A1/c3 ),
    .ZN(\A3/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M4/M2/_1_  (.A(\A3/A1/A2/A1/M4/s1 ),
    .B(\A3/A1/A2/A1/c3 ),
    .Z(Prod[43]));
 OR2_X1 \A3/A1/A2/A1/M4/_0_  (.A1(\A3/A1/A2/A1/M4/c1 ),
    .A2(\A3/A1/A2/A1/M4/c2 ),
    .ZN(\A3/A1/A2/c1 ));
 AND2_X1 \A3/A1/A2/A2/M1/M1/_0_  (.A1(v4[12]),
    .A2(s2[28]),
    .ZN(\A3/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M1/M1/_1_  (.A(v4[12]),
    .B(s2[28]),
    .Z(\A3/A1/A2/A2/M1/s1 ));
 AND2_X1 \A3/A1/A2/A2/M1/M2/_0_  (.A1(\A3/A1/A2/A2/M1/s1 ),
    .A2(\A3/A1/A2/c1 ),
    .ZN(\A3/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M1/M2/_1_  (.A(\A3/A1/A2/A2/M1/s1 ),
    .B(\A3/A1/A2/c1 ),
    .Z(Prod[44]));
 OR2_X1 \A3/A1/A2/A2/M1/_0_  (.A1(\A3/A1/A2/A2/M1/c1 ),
    .A2(\A3/A1/A2/A2/M1/c2 ),
    .ZN(\A3/A1/A2/A2/c1 ));
 AND2_X1 \A3/A1/A2/A2/M2/M1/_0_  (.A1(v4[13]),
    .A2(s2[29]),
    .ZN(\A3/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M2/M1/_1_  (.A(v4[13]),
    .B(s2[29]),
    .Z(\A3/A1/A2/A2/M2/s1 ));
 AND2_X1 \A3/A1/A2/A2/M2/M2/_0_  (.A1(\A3/A1/A2/A2/M2/s1 ),
    .A2(\A3/A1/A2/A2/c1 ),
    .ZN(\A3/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M2/M2/_1_  (.A(\A3/A1/A2/A2/M2/s1 ),
    .B(\A3/A1/A2/A2/c1 ),
    .Z(Prod[45]));
 OR2_X1 \A3/A1/A2/A2/M2/_0_  (.A1(\A3/A1/A2/A2/M2/c1 ),
    .A2(\A3/A1/A2/A2/M2/c2 ),
    .ZN(\A3/A1/A2/A2/c2 ));
 AND2_X1 \A3/A1/A2/A2/M3/M1/_0_  (.A1(v4[14]),
    .A2(s2[30]),
    .ZN(\A3/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M3/M1/_1_  (.A(v4[14]),
    .B(s2[30]),
    .Z(\A3/A1/A2/A2/M3/s1 ));
 AND2_X1 \A3/A1/A2/A2/M3/M2/_0_  (.A1(\A3/A1/A2/A2/M3/s1 ),
    .A2(\A3/A1/A2/A2/c2 ),
    .ZN(\A3/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M3/M2/_1_  (.A(\A3/A1/A2/A2/M3/s1 ),
    .B(\A3/A1/A2/A2/c2 ),
    .Z(Prod[46]));
 OR2_X2 \A3/A1/A2/A2/M3/_0_  (.A1(\A3/A1/A2/A2/M3/c1 ),
    .A2(\A3/A1/A2/A2/M3/c2 ),
    .ZN(\A3/A1/A2/A2/c3 ));
 AND2_X1 \A3/A1/A2/A2/M4/M1/_0_  (.A1(v4[15]),
    .A2(s2[31]),
    .ZN(\A3/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M4/M1/_1_  (.A(v4[15]),
    .B(s2[31]),
    .Z(\A3/A1/A2/A2/M4/s1 ));
 AND2_X1 \A3/A1/A2/A2/M4/M2/_0_  (.A1(\A3/A1/A2/A2/M4/s1 ),
    .A2(\A3/A1/A2/A2/c3 ),
    .ZN(\A3/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M4/M2/_1_  (.A(\A3/A1/A2/A2/M4/s1 ),
    .B(\A3/A1/A2/A2/c3 ),
    .Z(Prod[47]));
 OR2_X1 \A3/A1/A2/A2/M4/_0_  (.A1(\A3/A1/A2/A2/M4/c1 ),
    .A2(\A3/A1/A2/A2/M4/c2 ),
    .ZN(\A3/c1 ));
 AND2_X1 \A3/A2/A1/A1/M1/M1/_0_  (.A1(v4[16]),
    .A2(c3),
    .ZN(\A3/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M1/M1/_1_  (.A(v4[16]),
    .B(c3),
    .Z(\A3/A2/A1/A1/M1/s1 ));
 AND2_X1 \A3/A2/A1/A1/M1/M2/_0_  (.A1(\A3/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\A3/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M1/M2/_1_  (.A(\A3/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(Prod[48]));
 OR2_X1 \A3/A2/A1/A1/M1/_0_  (.A1(\A3/A2/A1/A1/M1/c1 ),
    .A2(\A3/A2/A1/A1/M1/c2 ),
    .ZN(\A3/A2/A1/A1/c1 ));
 AND2_X1 \A3/A2/A1/A1/M2/M1/_0_  (.A1(v4[17]),
    .A2(ground),
    .ZN(\A3/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M2/M1/_1_  (.A(v4[17]),
    .B(ground),
    .Z(\A3/A2/A1/A1/M2/s1 ));
 AND2_X1 \A3/A2/A1/A1/M2/M2/_0_  (.A1(\A3/A2/A1/A1/M2/s1 ),
    .A2(\A3/A2/A1/A1/c1 ),
    .ZN(\A3/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M2/M2/_1_  (.A(\A3/A2/A1/A1/M2/s1 ),
    .B(\A3/A2/A1/A1/c1 ),
    .Z(Prod[49]));
 OR2_X1 \A3/A2/A1/A1/M2/_0_  (.A1(\A3/A2/A1/A1/M2/c1 ),
    .A2(\A3/A2/A1/A1/M2/c2 ),
    .ZN(\A3/A2/A1/A1/c2 ));
 AND2_X1 \A3/A2/A1/A1/M3/M1/_0_  (.A1(v4[18]),
    .A2(ground),
    .ZN(\A3/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M3/M1/_1_  (.A(v4[18]),
    .B(ground),
    .Z(\A3/A2/A1/A1/M3/s1 ));
 AND2_X1 \A3/A2/A1/A1/M3/M2/_0_  (.A1(\A3/A2/A1/A1/M3/s1 ),
    .A2(\A3/A2/A1/A1/c2 ),
    .ZN(\A3/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M3/M2/_1_  (.A(\A3/A2/A1/A1/M3/s1 ),
    .B(\A3/A2/A1/A1/c2 ),
    .Z(Prod[50]));
 OR2_X1 \A3/A2/A1/A1/M3/_0_  (.A1(\A3/A2/A1/A1/M3/c1 ),
    .A2(\A3/A2/A1/A1/M3/c2 ),
    .ZN(\A3/A2/A1/A1/c3 ));
 AND2_X1 \A3/A2/A1/A1/M4/M1/_0_  (.A1(v4[19]),
    .A2(ground),
    .ZN(\A3/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M4/M1/_1_  (.A(v4[19]),
    .B(ground),
    .Z(\A3/A2/A1/A1/M4/s1 ));
 AND2_X1 \A3/A2/A1/A1/M4/M2/_0_  (.A1(\A3/A2/A1/A1/M4/s1 ),
    .A2(\A3/A2/A1/A1/c3 ),
    .ZN(\A3/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M4/M2/_1_  (.A(\A3/A2/A1/A1/M4/s1 ),
    .B(\A3/A2/A1/A1/c3 ),
    .Z(Prod[51]));
 OR2_X1 \A3/A2/A1/A1/M4/_0_  (.A1(\A3/A2/A1/A1/M4/c1 ),
    .A2(\A3/A2/A1/A1/M4/c2 ),
    .ZN(\A3/A2/A1/c1 ));
 AND2_X1 \A3/A2/A1/A2/M1/M1/_0_  (.A1(v4[20]),
    .A2(ground),
    .ZN(\A3/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M1/M1/_1_  (.A(v4[20]),
    .B(ground),
    .Z(\A3/A2/A1/A2/M1/s1 ));
 AND2_X1 \A3/A2/A1/A2/M1/M2/_0_  (.A1(\A3/A2/A1/A2/M1/s1 ),
    .A2(\A3/A2/A1/c1 ),
    .ZN(\A3/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M1/M2/_1_  (.A(\A3/A2/A1/A2/M1/s1 ),
    .B(\A3/A2/A1/c1 ),
    .Z(Prod[52]));
 OR2_X1 \A3/A2/A1/A2/M1/_0_  (.A1(\A3/A2/A1/A2/M1/c1 ),
    .A2(\A3/A2/A1/A2/M1/c2 ),
    .ZN(\A3/A2/A1/A2/c1 ));
 AND2_X1 \A3/A2/A1/A2/M2/M1/_0_  (.A1(v4[21]),
    .A2(ground),
    .ZN(\A3/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M2/M1/_1_  (.A(v4[21]),
    .B(ground),
    .Z(\A3/A2/A1/A2/M2/s1 ));
 AND2_X1 \A3/A2/A1/A2/M2/M2/_0_  (.A1(\A3/A2/A1/A2/M2/s1 ),
    .A2(\A3/A2/A1/A2/c1 ),
    .ZN(\A3/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M2/M2/_1_  (.A(\A3/A2/A1/A2/M2/s1 ),
    .B(\A3/A2/A1/A2/c1 ),
    .Z(Prod[53]));
 OR2_X1 \A3/A2/A1/A2/M2/_0_  (.A1(\A3/A2/A1/A2/M2/c1 ),
    .A2(\A3/A2/A1/A2/M2/c2 ),
    .ZN(\A3/A2/A1/A2/c2 ));
 AND2_X1 \A3/A2/A1/A2/M3/M1/_0_  (.A1(v4[22]),
    .A2(ground),
    .ZN(\A3/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M3/M1/_1_  (.A(v4[22]),
    .B(ground),
    .Z(\A3/A2/A1/A2/M3/s1 ));
 AND2_X1 \A3/A2/A1/A2/M3/M2/_0_  (.A1(\A3/A2/A1/A2/M3/s1 ),
    .A2(\A3/A2/A1/A2/c2 ),
    .ZN(\A3/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M3/M2/_1_  (.A(\A3/A2/A1/A2/M3/s1 ),
    .B(\A3/A2/A1/A2/c2 ),
    .Z(Prod[54]));
 OR2_X1 \A3/A2/A1/A2/M3/_0_  (.A1(\A3/A2/A1/A2/M3/c1 ),
    .A2(\A3/A2/A1/A2/M3/c2 ),
    .ZN(\A3/A2/A1/A2/c3 ));
 AND2_X1 \A3/A2/A1/A2/M4/M1/_0_  (.A1(v4[23]),
    .A2(ground),
    .ZN(\A3/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M4/M1/_1_  (.A(v4[23]),
    .B(ground),
    .Z(\A3/A2/A1/A2/M4/s1 ));
 AND2_X1 \A3/A2/A1/A2/M4/M2/_0_  (.A1(\A3/A2/A1/A2/M4/s1 ),
    .A2(\A3/A2/A1/A2/c3 ),
    .ZN(\A3/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M4/M2/_1_  (.A(\A3/A2/A1/A2/M4/s1 ),
    .B(\A3/A2/A1/A2/c3 ),
    .Z(Prod[55]));
 OR2_X1 \A3/A2/A1/A2/M4/_0_  (.A1(\A3/A2/A1/A2/M4/c1 ),
    .A2(\A3/A2/A1/A2/M4/c2 ),
    .ZN(\A3/A2/c1 ));
 AND2_X1 \A3/A2/A2/A1/M1/M1/_0_  (.A1(v4[24]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A3/A2/A2/A1/M1/M1/_1_  (.A(v4[24]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M1/s1 ));
 AND2_X1 \A3/A2/A2/A1/M1/M2/_0_  (.A1(\A3/A2/A2/A1/M1/s1 ),
    .A2(\A3/A2/c1 ),
    .ZN(\A3/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A3/A2/A2/A1/M1/M2/_1_  (.A(\A3/A2/A2/A1/M1/s1 ),
    .B(\A3/A2/c1 ),
    .Z(Prod[56]));
 OR2_X1 \A3/A2/A2/A1/M1/_0_  (.A1(\A3/A2/A2/A1/M1/c1 ),
    .A2(\A3/A2/A2/A1/M1/c2 ),
    .ZN(\A3/A2/A2/A1/c1 ));
 AND2_X1 \A3/A2/A2/A1/M2/M1/_0_  (.A1(v4[25]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M2/c1 ));
 XOR2_X1 \A3/A2/A2/A1/M2/M1/_1_  (.A(v4[25]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M2/s1 ));
 AND2_X1 \A3/A2/A2/A1/M2/M2/_0_  (.A1(\A3/A2/A2/A1/M2/s1 ),
    .A2(\A3/A2/A2/A1/c1 ),
    .ZN(\A3/A2/A2/A1/M2/c2 ));
 XOR2_X1 \A3/A2/A2/A1/M2/M2/_1_  (.A(\A3/A2/A2/A1/M2/s1 ),
    .B(\A3/A2/A2/A1/c1 ),
    .Z(Prod[57]));
 OR2_X1 \A3/A2/A2/A1/M2/_0_  (.A1(\A3/A2/A2/A1/M2/c1 ),
    .A2(\A3/A2/A2/A1/M2/c2 ),
    .ZN(\A3/A2/A2/A1/c2 ));
 AND2_X1 \A3/A2/A2/A1/M3/M1/_0_  (.A1(v4[26]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M3/c1 ));
 XOR2_X1 \A3/A2/A2/A1/M3/M1/_1_  (.A(v4[26]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M3/s1 ));
 AND2_X1 \A3/A2/A2/A1/M3/M2/_0_  (.A1(\A3/A2/A2/A1/M3/s1 ),
    .A2(\A3/A2/A2/A1/c2 ),
    .ZN(\A3/A2/A2/A1/M3/c2 ));
 XOR2_X1 \A3/A2/A2/A1/M3/M2/_1_  (.A(\A3/A2/A2/A1/M3/s1 ),
    .B(\A3/A2/A2/A1/c2 ),
    .Z(Prod[58]));
 OR2_X1 \A3/A2/A2/A1/M3/_0_  (.A1(\A3/A2/A2/A1/M3/c1 ),
    .A2(\A3/A2/A2/A1/M3/c2 ),
    .ZN(\A3/A2/A2/A1/c3 ));
 AND2_X1 \A3/A2/A2/A1/M4/M1/_0_  (.A1(v4[27]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M4/c1 ));
 XOR2_X1 \A3/A2/A2/A1/M4/M1/_1_  (.A(v4[27]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M4/s1 ));
 AND2_X1 \A3/A2/A2/A1/M4/M2/_0_  (.A1(\A3/A2/A2/A1/M4/s1 ),
    .A2(\A3/A2/A2/A1/c3 ),
    .ZN(\A3/A2/A2/A1/M4/c2 ));
 XOR2_X1 \A3/A2/A2/A1/M4/M2/_1_  (.A(\A3/A2/A2/A1/M4/s1 ),
    .B(\A3/A2/A2/A1/c3 ),
    .Z(Prod[59]));
 OR2_X1 \A3/A2/A2/A1/M4/_0_  (.A1(\A3/A2/A2/A1/M4/c1 ),
    .A2(\A3/A2/A2/A1/M4/c2 ),
    .ZN(\A3/A2/A2/c1 ));
 AND2_X1 \A3/A2/A2/A2/M1/M1/_0_  (.A1(v4[28]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M1/M1/_1_  (.A(v4[28]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M1/s1 ));
 AND2_X1 \A3/A2/A2/A2/M1/M2/_0_  (.A1(\A3/A2/A2/A2/M1/s1 ),
    .A2(\A3/A2/A2/c1 ),
    .ZN(\A3/A2/A2/A2/M1/c2 ));
 XOR2_X1 \A3/A2/A2/A2/M1/M2/_1_  (.A(\A3/A2/A2/A2/M1/s1 ),
    .B(\A3/A2/A2/c1 ),
    .Z(Prod[60]));
 OR2_X1 \A3/A2/A2/A2/M1/_0_  (.A1(\A3/A2/A2/A2/M1/c1 ),
    .A2(\A3/A2/A2/A2/M1/c2 ),
    .ZN(\A3/A2/A2/A2/c1 ));
 AND2_X1 \A3/A2/A2/A2/M2/M1/_0_  (.A1(v4[29]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M2/M1/_1_  (.A(v4[29]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M2/s1 ));
 AND2_X1 \A3/A2/A2/A2/M2/M2/_0_  (.A1(\A3/A2/A2/A2/M2/s1 ),
    .A2(\A3/A2/A2/A2/c1 ),
    .ZN(\A3/A2/A2/A2/M2/c2 ));
 XOR2_X1 \A3/A2/A2/A2/M2/M2/_1_  (.A(\A3/A2/A2/A2/M2/s1 ),
    .B(\A3/A2/A2/A2/c1 ),
    .Z(Prod[61]));
 OR2_X1 \A3/A2/A2/A2/M2/_0_  (.A1(\A3/A2/A2/A2/M2/c1 ),
    .A2(\A3/A2/A2/A2/M2/c2 ),
    .ZN(\A3/A2/A2/A2/c2 ));
 AND2_X1 \A3/A2/A2/A2/M3/M1/_0_  (.A1(v4[30]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M3/c1 ));
 XOR2_X1 \A3/A2/A2/A2/M3/M1/_1_  (.A(v4[30]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M3/s1 ));
 AND2_X1 \A3/A2/A2/A2/M3/M2/_0_  (.A1(\A3/A2/A2/A2/M3/s1 ),
    .A2(\A3/A2/A2/A2/c2 ),
    .ZN(\A3/A2/A2/A2/M3/c2 ));
 XOR2_X1 \A3/A2/A2/A2/M3/M2/_1_  (.A(\A3/A2/A2/A2/M3/s1 ),
    .B(\A3/A2/A2/A2/c2 ),
    .Z(Prod[62]));
 OR2_X1 \A3/A2/A2/A2/M3/_0_  (.A1(\A3/A2/A2/A2/M3/c1 ),
    .A2(\A3/A2/A2/A2/M3/c2 ),
    .ZN(\A3/A2/A2/A2/c3 ));
 AND2_X1 \A3/A2/A2/A2/M4/M1/_0_  (.A1(v4[31]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M4/M1/_1_  (.A(v4[31]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M4/s1 ));
 AND2_X1 \A3/A2/A2/A2/M4/M2/_0_  (.A1(\A3/A2/A2/A2/M4/s1 ),
    .A2(\A3/A2/A2/A2/c3 ),
    .ZN(\A3/A2/A2/A2/M4/c2 ));
 XOR2_X1 \A3/A2/A2/A2/M4/M2/_1_  (.A(\A3/A2/A2/A2/M4/s1 ),
    .B(\A3/A2/A2/A2/c3 ),
    .Z(Prod[63]));
 OR2_X1 \A3/A2/A2/A2/M4/_0_  (.A1(\A3/A2/A2/A2/M4/c1 ),
    .A2(\A3/A2/A2/A2/M4/c2 ),
    .ZN(overflow));
 AND2_X1 \V1/A1/A1/A1/M1/M1/_0_  (.A1(\V1/v2 [0]),
    .A2(\V1/v3 [0]),
    .ZN(\V1/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M1/M1/_1_  (.A(\V1/v2 [0]),
    .B(\V1/v3 [0]),
    .Z(\V1/A1/A1/A1/M1/s1 ));
 AND2_X1 \V1/A1/A1/A1/M1/M2/_0_  (.A1(\V1/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M1/M2/_1_  (.A(\V1/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/s1 [0]));
 OR2_X1 \V1/A1/A1/A1/M1/_0_  (.A1(\V1/A1/A1/A1/M1/c1 ),
    .A2(\V1/A1/A1/A1/M1/c2 ),
    .ZN(\V1/A1/A1/A1/c1 ));
 AND2_X1 \V1/A1/A1/A1/M2/M1/_0_  (.A1(\V1/v2 [1]),
    .A2(\V1/v3 [1]),
    .ZN(\V1/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M2/M1/_1_  (.A(\V1/v2 [1]),
    .B(\V1/v3 [1]),
    .Z(\V1/A1/A1/A1/M2/s1 ));
 AND2_X1 \V1/A1/A1/A1/M2/M2/_0_  (.A1(\V1/A1/A1/A1/M2/s1 ),
    .A2(\V1/A1/A1/A1/c1 ),
    .ZN(\V1/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M2/M2/_1_  (.A(\V1/A1/A1/A1/M2/s1 ),
    .B(\V1/A1/A1/A1/c1 ),
    .Z(\V1/s1 [1]));
 OR2_X1 \V1/A1/A1/A1/M2/_0_  (.A1(\V1/A1/A1/A1/M2/c1 ),
    .A2(\V1/A1/A1/A1/M2/c2 ),
    .ZN(\V1/A1/A1/A1/c2 ));
 AND2_X1 \V1/A1/A1/A1/M3/M1/_0_  (.A1(\V1/v2 [2]),
    .A2(\V1/v3 [2]),
    .ZN(\V1/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M3/M1/_1_  (.A(\V1/v2 [2]),
    .B(\V1/v3 [2]),
    .Z(\V1/A1/A1/A1/M3/s1 ));
 AND2_X1 \V1/A1/A1/A1/M3/M2/_0_  (.A1(\V1/A1/A1/A1/M3/s1 ),
    .A2(\V1/A1/A1/A1/c2 ),
    .ZN(\V1/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M3/M2/_1_  (.A(\V1/A1/A1/A1/M3/s1 ),
    .B(\V1/A1/A1/A1/c2 ),
    .Z(\V1/s1 [2]));
 OR2_X1 \V1/A1/A1/A1/M3/_0_  (.A1(\V1/A1/A1/A1/M3/c1 ),
    .A2(\V1/A1/A1/A1/M3/c2 ),
    .ZN(\V1/A1/A1/A1/c3 ));
 AND2_X1 \V1/A1/A1/A1/M4/M1/_0_  (.A1(\V1/v2 [3]),
    .A2(\V1/v3 [3]),
    .ZN(\V1/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M4/M1/_1_  (.A(\V1/v2 [3]),
    .B(\V1/v3 [3]),
    .Z(\V1/A1/A1/A1/M4/s1 ));
 AND2_X1 \V1/A1/A1/A1/M4/M2/_0_  (.A1(\V1/A1/A1/A1/M4/s1 ),
    .A2(\V1/A1/A1/A1/c3 ),
    .ZN(\V1/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M4/M2/_1_  (.A(\V1/A1/A1/A1/M4/s1 ),
    .B(\V1/A1/A1/A1/c3 ),
    .Z(\V1/s1 [3]));
 OR2_X1 \V1/A1/A1/A1/M4/_0_  (.A1(\V1/A1/A1/A1/M4/c1 ),
    .A2(\V1/A1/A1/A1/M4/c2 ),
    .ZN(\V1/A1/A1/c1 ));
 AND2_X1 \V1/A1/A1/A2/M1/M1/_0_  (.A1(\V1/v2 [4]),
    .A2(\V1/v3 [4]),
    .ZN(\V1/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M1/M1/_1_  (.A(\V1/v2 [4]),
    .B(\V1/v3 [4]),
    .Z(\V1/A1/A1/A2/M1/s1 ));
 AND2_X1 \V1/A1/A1/A2/M1/M2/_0_  (.A1(\V1/A1/A1/A2/M1/s1 ),
    .A2(\V1/A1/A1/c1 ),
    .ZN(\V1/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M1/M2/_1_  (.A(\V1/A1/A1/A2/M1/s1 ),
    .B(\V1/A1/A1/c1 ),
    .Z(\V1/s1 [4]));
 OR2_X1 \V1/A1/A1/A2/M1/_0_  (.A1(\V1/A1/A1/A2/M1/c1 ),
    .A2(\V1/A1/A1/A2/M1/c2 ),
    .ZN(\V1/A1/A1/A2/c1 ));
 AND2_X1 \V1/A1/A1/A2/M2/M1/_0_  (.A1(\V1/v2 [5]),
    .A2(\V1/v3 [5]),
    .ZN(\V1/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M2/M1/_1_  (.A(\V1/v2 [5]),
    .B(\V1/v3 [5]),
    .Z(\V1/A1/A1/A2/M2/s1 ));
 AND2_X1 \V1/A1/A1/A2/M2/M2/_0_  (.A1(\V1/A1/A1/A2/M2/s1 ),
    .A2(\V1/A1/A1/A2/c1 ),
    .ZN(\V1/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M2/M2/_1_  (.A(\V1/A1/A1/A2/M2/s1 ),
    .B(\V1/A1/A1/A2/c1 ),
    .Z(\V1/s1 [5]));
 OR2_X1 \V1/A1/A1/A2/M2/_0_  (.A1(\V1/A1/A1/A2/M2/c1 ),
    .A2(\V1/A1/A1/A2/M2/c2 ),
    .ZN(\V1/A1/A1/A2/c2 ));
 AND2_X1 \V1/A1/A1/A2/M3/M1/_0_  (.A1(\V1/v2 [6]),
    .A2(\V1/v3 [6]),
    .ZN(\V1/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M3/M1/_1_  (.A(\V1/v2 [6]),
    .B(\V1/v3 [6]),
    .Z(\V1/A1/A1/A2/M3/s1 ));
 AND2_X1 \V1/A1/A1/A2/M3/M2/_0_  (.A1(\V1/A1/A1/A2/M3/s1 ),
    .A2(\V1/A1/A1/A2/c2 ),
    .ZN(\V1/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M3/M2/_1_  (.A(\V1/A1/A1/A2/M3/s1 ),
    .B(\V1/A1/A1/A2/c2 ),
    .Z(\V1/s1 [6]));
 OR2_X1 \V1/A1/A1/A2/M3/_0_  (.A1(\V1/A1/A1/A2/M3/c1 ),
    .A2(\V1/A1/A1/A2/M3/c2 ),
    .ZN(\V1/A1/A1/A2/c3 ));
 AND2_X1 \V1/A1/A1/A2/M4/M1/_0_  (.A1(\V1/v2 [7]),
    .A2(\V1/v3 [7]),
    .ZN(\V1/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M4/M1/_1_  (.A(\V1/v2 [7]),
    .B(\V1/v3 [7]),
    .Z(\V1/A1/A1/A2/M4/s1 ));
 AND2_X1 \V1/A1/A1/A2/M4/M2/_0_  (.A1(\V1/A1/A1/A2/M4/s1 ),
    .A2(\V1/A1/A1/A2/c3 ),
    .ZN(\V1/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M4/M2/_1_  (.A(\V1/A1/A1/A2/M4/s1 ),
    .B(\V1/A1/A1/A2/c3 ),
    .Z(\V1/s1 [7]));
 OR2_X1 \V1/A1/A1/A2/M4/_0_  (.A1(\V1/A1/A1/A2/M4/c1 ),
    .A2(\V1/A1/A1/A2/M4/c2 ),
    .ZN(\V1/A1/c1 ));
 AND2_X1 \V1/A1/A2/A1/M1/M1/_0_  (.A1(\V1/v2 [8]),
    .A2(\V1/v3 [8]),
    .ZN(\V1/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M1/M1/_1_  (.A(\V1/v2 [8]),
    .B(\V1/v3 [8]),
    .Z(\V1/A1/A2/A1/M1/s1 ));
 AND2_X1 \V1/A1/A2/A1/M1/M2/_0_  (.A1(\V1/A1/A2/A1/M1/s1 ),
    .A2(\V1/A1/c1 ),
    .ZN(\V1/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M1/M2/_1_  (.A(\V1/A1/A2/A1/M1/s1 ),
    .B(\V1/A1/c1 ),
    .Z(\V1/s1 [8]));
 OR2_X1 \V1/A1/A2/A1/M1/_0_  (.A1(\V1/A1/A2/A1/M1/c1 ),
    .A2(\V1/A1/A2/A1/M1/c2 ),
    .ZN(\V1/A1/A2/A1/c1 ));
 AND2_X1 \V1/A1/A2/A1/M2/M1/_0_  (.A1(\V1/v2 [9]),
    .A2(\V1/v3 [9]),
    .ZN(\V1/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M2/M1/_1_  (.A(\V1/v2 [9]),
    .B(\V1/v3 [9]),
    .Z(\V1/A1/A2/A1/M2/s1 ));
 AND2_X1 \V1/A1/A2/A1/M2/M2/_0_  (.A1(\V1/A1/A2/A1/M2/s1 ),
    .A2(\V1/A1/A2/A1/c1 ),
    .ZN(\V1/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M2/M2/_1_  (.A(\V1/A1/A2/A1/M2/s1 ),
    .B(\V1/A1/A2/A1/c1 ),
    .Z(\V1/s1 [9]));
 OR2_X1 \V1/A1/A2/A1/M2/_0_  (.A1(\V1/A1/A2/A1/M2/c1 ),
    .A2(\V1/A1/A2/A1/M2/c2 ),
    .ZN(\V1/A1/A2/A1/c2 ));
 AND2_X1 \V1/A1/A2/A1/M3/M1/_0_  (.A1(\V1/v2 [10]),
    .A2(\V1/v3 [10]),
    .ZN(\V1/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M3/M1/_1_  (.A(\V1/v2 [10]),
    .B(\V1/v3 [10]),
    .Z(\V1/A1/A2/A1/M3/s1 ));
 AND2_X1 \V1/A1/A2/A1/M3/M2/_0_  (.A1(\V1/A1/A2/A1/M3/s1 ),
    .A2(\V1/A1/A2/A1/c2 ),
    .ZN(\V1/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M3/M2/_1_  (.A(\V1/A1/A2/A1/M3/s1 ),
    .B(\V1/A1/A2/A1/c2 ),
    .Z(\V1/s1 [10]));
 OR2_X1 \V1/A1/A2/A1/M3/_0_  (.A1(\V1/A1/A2/A1/M3/c1 ),
    .A2(\V1/A1/A2/A1/M3/c2 ),
    .ZN(\V1/A1/A2/A1/c3 ));
 AND2_X1 \V1/A1/A2/A1/M4/M1/_0_  (.A1(\V1/v2 [11]),
    .A2(\V1/v3 [11]),
    .ZN(\V1/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M4/M1/_1_  (.A(\V1/v2 [11]),
    .B(\V1/v3 [11]),
    .Z(\V1/A1/A2/A1/M4/s1 ));
 AND2_X1 \V1/A1/A2/A1/M4/M2/_0_  (.A1(\V1/A1/A2/A1/M4/s1 ),
    .A2(\V1/A1/A2/A1/c3 ),
    .ZN(\V1/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M4/M2/_1_  (.A(\V1/A1/A2/A1/M4/s1 ),
    .B(\V1/A1/A2/A1/c3 ),
    .Z(\V1/s1 [11]));
 OR2_X1 \V1/A1/A2/A1/M4/_0_  (.A1(\V1/A1/A2/A1/M4/c1 ),
    .A2(\V1/A1/A2/A1/M4/c2 ),
    .ZN(\V1/A1/A2/c1 ));
 AND2_X1 \V1/A1/A2/A2/M1/M1/_0_  (.A1(\V1/v2 [12]),
    .A2(\V1/v3 [12]),
    .ZN(\V1/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M1/M1/_1_  (.A(\V1/v2 [12]),
    .B(\V1/v3 [12]),
    .Z(\V1/A1/A2/A2/M1/s1 ));
 AND2_X1 \V1/A1/A2/A2/M1/M2/_0_  (.A1(\V1/A1/A2/A2/M1/s1 ),
    .A2(\V1/A1/A2/c1 ),
    .ZN(\V1/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M1/M2/_1_  (.A(\V1/A1/A2/A2/M1/s1 ),
    .B(\V1/A1/A2/c1 ),
    .Z(\V1/s1 [12]));
 OR2_X1 \V1/A1/A2/A2/M1/_0_  (.A1(\V1/A1/A2/A2/M1/c1 ),
    .A2(\V1/A1/A2/A2/M1/c2 ),
    .ZN(\V1/A1/A2/A2/c1 ));
 AND2_X1 \V1/A1/A2/A2/M2/M1/_0_  (.A1(\V1/v2 [13]),
    .A2(\V1/v3 [13]),
    .ZN(\V1/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M2/M1/_1_  (.A(\V1/v2 [13]),
    .B(\V1/v3 [13]),
    .Z(\V1/A1/A2/A2/M2/s1 ));
 AND2_X1 \V1/A1/A2/A2/M2/M2/_0_  (.A1(\V1/A1/A2/A2/M2/s1 ),
    .A2(\V1/A1/A2/A2/c1 ),
    .ZN(\V1/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M2/M2/_1_  (.A(\V1/A1/A2/A2/M2/s1 ),
    .B(\V1/A1/A2/A2/c1 ),
    .Z(\V1/s1 [13]));
 OR2_X1 \V1/A1/A2/A2/M2/_0_  (.A1(\V1/A1/A2/A2/M2/c1 ),
    .A2(\V1/A1/A2/A2/M2/c2 ),
    .ZN(\V1/A1/A2/A2/c2 ));
 AND2_X1 \V1/A1/A2/A2/M3/M1/_0_  (.A1(\V1/v2 [14]),
    .A2(\V1/v3 [14]),
    .ZN(\V1/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M3/M1/_1_  (.A(\V1/v2 [14]),
    .B(\V1/v3 [14]),
    .Z(\V1/A1/A2/A2/M3/s1 ));
 AND2_X1 \V1/A1/A2/A2/M3/M2/_0_  (.A1(\V1/A1/A2/A2/M3/s1 ),
    .A2(\V1/A1/A2/A2/c2 ),
    .ZN(\V1/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M3/M2/_1_  (.A(\V1/A1/A2/A2/M3/s1 ),
    .B(\V1/A1/A2/A2/c2 ),
    .Z(\V1/s1 [14]));
 OR2_X1 \V1/A1/A2/A2/M3/_0_  (.A1(\V1/A1/A2/A2/M3/c1 ),
    .A2(\V1/A1/A2/A2/M3/c2 ),
    .ZN(\V1/A1/A2/A2/c3 ));
 AND2_X1 \V1/A1/A2/A2/M4/M1/_0_  (.A1(\V1/v2 [15]),
    .A2(\V1/v3 [15]),
    .ZN(\V1/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M4/M1/_1_  (.A(\V1/v2 [15]),
    .B(\V1/v3 [15]),
    .Z(\V1/A1/A2/A2/M4/s1 ));
 AND2_X1 \V1/A1/A2/A2/M4/M2/_0_  (.A1(\V1/A1/A2/A2/M4/s1 ),
    .A2(\V1/A1/A2/A2/c3 ),
    .ZN(\V1/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M4/M2/_1_  (.A(\V1/A1/A2/A2/M4/s1 ),
    .B(\V1/A1/A2/A2/c3 ),
    .Z(\V1/s1 [15]));
 OR2_X1 \V1/A1/A2/A2/M4/_0_  (.A1(\V1/A1/A2/A2/M4/c1 ),
    .A2(\V1/A1/A2/A2/M4/c2 ),
    .ZN(\V1/c1 ));
 AND2_X1 \V1/A2/A1/A1/M1/M1/_0_  (.A1(\V1/s1 [0]),
    .A2(\V1/v1 [8]),
    .ZN(\V1/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M1/M1/_1_  (.A(\V1/s1 [0]),
    .B(\V1/v1 [8]),
    .Z(\V1/A2/A1/A1/M1/s1 ));
 AND2_X1 \V1/A2/A1/A1/M1/M2/_0_  (.A1(\V1/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M1/M2/_1_  (.A(\V1/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v1[8]));
 OR2_X1 \V1/A2/A1/A1/M1/_0_  (.A1(\V1/A2/A1/A1/M1/c1 ),
    .A2(\V1/A2/A1/A1/M1/c2 ),
    .ZN(\V1/A2/A1/A1/c1 ));
 AND2_X1 \V1/A2/A1/A1/M2/M1/_0_  (.A1(\V1/s1 [1]),
    .A2(\V1/v1 [9]),
    .ZN(\V1/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M2/M1/_1_  (.A(\V1/s1 [1]),
    .B(\V1/v1 [9]),
    .Z(\V1/A2/A1/A1/M2/s1 ));
 AND2_X1 \V1/A2/A1/A1/M2/M2/_0_  (.A1(\V1/A2/A1/A1/M2/s1 ),
    .A2(\V1/A2/A1/A1/c1 ),
    .ZN(\V1/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M2/M2/_1_  (.A(\V1/A2/A1/A1/M2/s1 ),
    .B(\V1/A2/A1/A1/c1 ),
    .Z(v1[9]));
 OR2_X1 \V1/A2/A1/A1/M2/_0_  (.A1(\V1/A2/A1/A1/M2/c1 ),
    .A2(\V1/A2/A1/A1/M2/c2 ),
    .ZN(\V1/A2/A1/A1/c2 ));
 AND2_X1 \V1/A2/A1/A1/M3/M1/_0_  (.A1(\V1/s1 [2]),
    .A2(\V1/v1 [10]),
    .ZN(\V1/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M3/M1/_1_  (.A(\V1/s1 [2]),
    .B(\V1/v1 [10]),
    .Z(\V1/A2/A1/A1/M3/s1 ));
 AND2_X1 \V1/A2/A1/A1/M3/M2/_0_  (.A1(\V1/A2/A1/A1/M3/s1 ),
    .A2(\V1/A2/A1/A1/c2 ),
    .ZN(\V1/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M3/M2/_1_  (.A(\V1/A2/A1/A1/M3/s1 ),
    .B(\V1/A2/A1/A1/c2 ),
    .Z(v1[10]));
 OR2_X1 \V1/A2/A1/A1/M3/_0_  (.A1(\V1/A2/A1/A1/M3/c1 ),
    .A2(\V1/A2/A1/A1/M3/c2 ),
    .ZN(\V1/A2/A1/A1/c3 ));
 AND2_X1 \V1/A2/A1/A1/M4/M1/_0_  (.A1(\V1/s1 [3]),
    .A2(\V1/v1 [11]),
    .ZN(\V1/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M4/M1/_1_  (.A(\V1/s1 [3]),
    .B(\V1/v1 [11]),
    .Z(\V1/A2/A1/A1/M4/s1 ));
 AND2_X1 \V1/A2/A1/A1/M4/M2/_0_  (.A1(\V1/A2/A1/A1/M4/s1 ),
    .A2(\V1/A2/A1/A1/c3 ),
    .ZN(\V1/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M4/M2/_1_  (.A(\V1/A2/A1/A1/M4/s1 ),
    .B(\V1/A2/A1/A1/c3 ),
    .Z(v1[11]));
 OR2_X1 \V1/A2/A1/A1/M4/_0_  (.A1(\V1/A2/A1/A1/M4/c1 ),
    .A2(\V1/A2/A1/A1/M4/c2 ),
    .ZN(\V1/A2/A1/c1 ));
 AND2_X1 \V1/A2/A1/A2/M1/M1/_0_  (.A1(\V1/s1 [4]),
    .A2(\V1/v1 [12]),
    .ZN(\V1/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M1/M1/_1_  (.A(\V1/s1 [4]),
    .B(\V1/v1 [12]),
    .Z(\V1/A2/A1/A2/M1/s1 ));
 AND2_X1 \V1/A2/A1/A2/M1/M2/_0_  (.A1(\V1/A2/A1/A2/M1/s1 ),
    .A2(\V1/A2/A1/c1 ),
    .ZN(\V1/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M1/M2/_1_  (.A(\V1/A2/A1/A2/M1/s1 ),
    .B(\V1/A2/A1/c1 ),
    .Z(v1[12]));
 OR2_X2 \V1/A2/A1/A2/M1/_0_  (.A1(\V1/A2/A1/A2/M1/c1 ),
    .A2(\V1/A2/A1/A2/M1/c2 ),
    .ZN(\V1/A2/A1/A2/c1 ));
 AND2_X1 \V1/A2/A1/A2/M2/M1/_0_  (.A1(\V1/s1 [5]),
    .A2(\V1/v1 [13]),
    .ZN(\V1/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M2/M1/_1_  (.A(\V1/s1 [5]),
    .B(\V1/v1 [13]),
    .Z(\V1/A2/A1/A2/M2/s1 ));
 AND2_X1 \V1/A2/A1/A2/M2/M2/_0_  (.A1(\V1/A2/A1/A2/M2/s1 ),
    .A2(\V1/A2/A1/A2/c1 ),
    .ZN(\V1/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M2/M2/_1_  (.A(\V1/A2/A1/A2/M2/s1 ),
    .B(\V1/A2/A1/A2/c1 ),
    .Z(v1[13]));
 OR2_X1 \V1/A2/A1/A2/M2/_0_  (.A1(\V1/A2/A1/A2/M2/c1 ),
    .A2(\V1/A2/A1/A2/M2/c2 ),
    .ZN(\V1/A2/A1/A2/c2 ));
 AND2_X1 \V1/A2/A1/A2/M3/M1/_0_  (.A1(\V1/s1 [6]),
    .A2(\V1/v1 [14]),
    .ZN(\V1/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M3/M1/_1_  (.A(\V1/s1 [6]),
    .B(\V1/v1 [14]),
    .Z(\V1/A2/A1/A2/M3/s1 ));
 AND2_X1 \V1/A2/A1/A2/M3/M2/_0_  (.A1(\V1/A2/A1/A2/M3/s1 ),
    .A2(\V1/A2/A1/A2/c2 ),
    .ZN(\V1/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M3/M2/_1_  (.A(\V1/A2/A1/A2/M3/s1 ),
    .B(\V1/A2/A1/A2/c2 ),
    .Z(v1[14]));
 OR2_X1 \V1/A2/A1/A2/M3/_0_  (.A1(\V1/A2/A1/A2/M3/c1 ),
    .A2(\V1/A2/A1/A2/M3/c2 ),
    .ZN(\V1/A2/A1/A2/c3 ));
 AND2_X1 \V1/A2/A1/A2/M4/M1/_0_  (.A1(\V1/s1 [7]),
    .A2(\V1/v1 [15]),
    .ZN(\V1/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M4/M1/_1_  (.A(\V1/s1 [7]),
    .B(\V1/v1 [15]),
    .Z(\V1/A2/A1/A2/M4/s1 ));
 AND2_X1 \V1/A2/A1/A2/M4/M2/_0_  (.A1(\V1/A2/A1/A2/M4/s1 ),
    .A2(\V1/A2/A1/A2/c3 ),
    .ZN(\V1/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M4/M2/_1_  (.A(\V1/A2/A1/A2/M4/s1 ),
    .B(\V1/A2/A1/A2/c3 ),
    .Z(v1[15]));
 OR2_X2 \V1/A2/A1/A2/M4/_0_  (.A1(\V1/A2/A1/A2/M4/c1 ),
    .A2(\V1/A2/A1/A2/M4/c2 ),
    .ZN(\V1/A2/c1 ));
 AND2_X1 \V1/A2/A2/A1/M1/M1/_0_  (.A1(\V1/s1 [8]),
    .A2(ground),
    .ZN(\V1/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M1/M1/_1_  (.A(\V1/s1 [8]),
    .B(ground),
    .Z(\V1/A2/A2/A1/M1/s1 ));
 AND2_X1 \V1/A2/A2/A1/M1/M2/_0_  (.A1(\V1/A2/A2/A1/M1/s1 ),
    .A2(\V1/A2/c1 ),
    .ZN(\V1/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M1/M2/_1_  (.A(\V1/A2/A2/A1/M1/s1 ),
    .B(\V1/A2/c1 ),
    .Z(\V1/s2 [8]));
 OR2_X1 \V1/A2/A2/A1/M1/_0_  (.A1(\V1/A2/A2/A1/M1/c1 ),
    .A2(\V1/A2/A2/A1/M1/c2 ),
    .ZN(\V1/A2/A2/A1/c1 ));
 AND2_X1 \V1/A2/A2/A1/M2/M1/_0_  (.A1(\V1/s1 [9]),
    .A2(ground),
    .ZN(\V1/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M2/M1/_1_  (.A(\V1/s1 [9]),
    .B(ground),
    .Z(\V1/A2/A2/A1/M2/s1 ));
 AND2_X1 \V1/A2/A2/A1/M2/M2/_0_  (.A1(\V1/A2/A2/A1/M2/s1 ),
    .A2(\V1/A2/A2/A1/c1 ),
    .ZN(\V1/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M2/M2/_1_  (.A(\V1/A2/A2/A1/M2/s1 ),
    .B(\V1/A2/A2/A1/c1 ),
    .Z(\V1/s2 [9]));
 OR2_X1 \V1/A2/A2/A1/M2/_0_  (.A1(\V1/A2/A2/A1/M2/c1 ),
    .A2(\V1/A2/A2/A1/M2/c2 ),
    .ZN(\V1/A2/A2/A1/c2 ));
 AND2_X1 \V1/A2/A2/A1/M3/M1/_0_  (.A1(\V1/s1 [10]),
    .A2(ground),
    .ZN(\V1/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M3/M1/_1_  (.A(\V1/s1 [10]),
    .B(ground),
    .Z(\V1/A2/A2/A1/M3/s1 ));
 AND2_X1 \V1/A2/A2/A1/M3/M2/_0_  (.A1(\V1/A2/A2/A1/M3/s1 ),
    .A2(\V1/A2/A2/A1/c2 ),
    .ZN(\V1/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M3/M2/_1_  (.A(\V1/A2/A2/A1/M3/s1 ),
    .B(\V1/A2/A2/A1/c2 ),
    .Z(\V1/s2 [10]));
 OR2_X1 \V1/A2/A2/A1/M3/_0_  (.A1(\V1/A2/A2/A1/M3/c1 ),
    .A2(\V1/A2/A2/A1/M3/c2 ),
    .ZN(\V1/A2/A2/A1/c3 ));
 AND2_X1 \V1/A2/A2/A1/M4/M1/_0_  (.A1(\V1/s1 [11]),
    .A2(ground),
    .ZN(\V1/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M4/M1/_1_  (.A(\V1/s1 [11]),
    .B(ground),
    .Z(\V1/A2/A2/A1/M4/s1 ));
 AND2_X1 \V1/A2/A2/A1/M4/M2/_0_  (.A1(\V1/A2/A2/A1/M4/s1 ),
    .A2(\V1/A2/A2/A1/c3 ),
    .ZN(\V1/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M4/M2/_1_  (.A(\V1/A2/A2/A1/M4/s1 ),
    .B(\V1/A2/A2/A1/c3 ),
    .Z(\V1/s2 [11]));
 OR2_X1 \V1/A2/A2/A1/M4/_0_  (.A1(\V1/A2/A2/A1/M4/c1 ),
    .A2(\V1/A2/A2/A1/M4/c2 ),
    .ZN(\V1/A2/A2/c1 ));
 AND2_X1 \V1/A2/A2/A2/M1/M1/_0_  (.A1(\V1/s1 [12]),
    .A2(ground),
    .ZN(\V1/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M1/M1/_1_  (.A(\V1/s1 [12]),
    .B(ground),
    .Z(\V1/A2/A2/A2/M1/s1 ));
 AND2_X1 \V1/A2/A2/A2/M1/M2/_0_  (.A1(\V1/A2/A2/A2/M1/s1 ),
    .A2(\V1/A2/A2/c1 ),
    .ZN(\V1/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M1/M2/_1_  (.A(\V1/A2/A2/A2/M1/s1 ),
    .B(\V1/A2/A2/c1 ),
    .Z(\V1/s2 [12]));
 OR2_X1 \V1/A2/A2/A2/M1/_0_  (.A1(\V1/A2/A2/A2/M1/c1 ),
    .A2(\V1/A2/A2/A2/M1/c2 ),
    .ZN(\V1/A2/A2/A2/c1 ));
 AND2_X1 \V1/A2/A2/A2/M2/M1/_0_  (.A1(\V1/s1 [13]),
    .A2(ground),
    .ZN(\V1/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M2/M1/_1_  (.A(\V1/s1 [13]),
    .B(ground),
    .Z(\V1/A2/A2/A2/M2/s1 ));
 AND2_X1 \V1/A2/A2/A2/M2/M2/_0_  (.A1(\V1/A2/A2/A2/M2/s1 ),
    .A2(\V1/A2/A2/A2/c1 ),
    .ZN(\V1/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M2/M2/_1_  (.A(\V1/A2/A2/A2/M2/s1 ),
    .B(\V1/A2/A2/A2/c1 ),
    .Z(\V1/s2 [13]));
 OR2_X1 \V1/A2/A2/A2/M2/_0_  (.A1(\V1/A2/A2/A2/M2/c1 ),
    .A2(\V1/A2/A2/A2/M2/c2 ),
    .ZN(\V1/A2/A2/A2/c2 ));
 AND2_X1 \V1/A2/A2/A2/M3/M1/_0_  (.A1(\V1/s1 [14]),
    .A2(ground),
    .ZN(\V1/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M3/M1/_1_  (.A(\V1/s1 [14]),
    .B(ground),
    .Z(\V1/A2/A2/A2/M3/s1 ));
 AND2_X1 \V1/A2/A2/A2/M3/M2/_0_  (.A1(\V1/A2/A2/A2/M3/s1 ),
    .A2(\V1/A2/A2/A2/c2 ),
    .ZN(\V1/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M3/M2/_1_  (.A(\V1/A2/A2/A2/M3/s1 ),
    .B(\V1/A2/A2/A2/c2 ),
    .Z(\V1/s2 [14]));
 OR2_X1 \V1/A2/A2/A2/M3/_0_  (.A1(\V1/A2/A2/A2/M3/c1 ),
    .A2(\V1/A2/A2/A2/M3/c2 ),
    .ZN(\V1/A2/A2/A2/c3 ));
 AND2_X1 \V1/A2/A2/A2/M4/M1/_0_  (.A1(\V1/s1 [15]),
    .A2(ground),
    .ZN(\V1/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M4/M1/_1_  (.A(\V1/s1 [15]),
    .B(ground),
    .Z(\V1/A2/A2/A2/M4/s1 ));
 AND2_X1 \V1/A2/A2/A2/M4/M2/_0_  (.A1(\V1/A2/A2/A2/M4/s1 ),
    .A2(\V1/A2/A2/A2/c3 ),
    .ZN(\V1/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M4/M2/_1_  (.A(\V1/A2/A2/A2/M4/s1 ),
    .B(\V1/A2/A2/A2/c3 ),
    .Z(\V1/s2 [15]));
 OR2_X1 \V1/A2/A2/A2/M4/_0_  (.A1(\V1/A2/A2/A2/M4/c1 ),
    .A2(\V1/A2/A2/A2/M4/c2 ),
    .ZN(\V1/c2 ));
 AND2_X1 \V1/A3/A1/A1/M1/M1/_0_  (.A1(\V1/v4 [0]),
    .A2(\V1/s2 [8]),
    .ZN(\V1/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M1/M1/_1_  (.A(\V1/v4 [0]),
    .B(\V1/s2 [8]),
    .Z(\V1/A3/A1/A1/M1/s1 ));
 AND2_X1 \V1/A3/A1/A1/M1/M2/_0_  (.A1(\V1/A3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M1/M2/_1_  (.A(\V1/A3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v1[16]));
 OR2_X1 \V1/A3/A1/A1/M1/_0_  (.A1(\V1/A3/A1/A1/M1/c1 ),
    .A2(\V1/A3/A1/A1/M1/c2 ),
    .ZN(\V1/A3/A1/A1/c1 ));
 AND2_X1 \V1/A3/A1/A1/M2/M1/_0_  (.A1(\V1/v4 [1]),
    .A2(\V1/s2 [9]),
    .ZN(\V1/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M2/M1/_1_  (.A(\V1/v4 [1]),
    .B(\V1/s2 [9]),
    .Z(\V1/A3/A1/A1/M2/s1 ));
 AND2_X1 \V1/A3/A1/A1/M2/M2/_0_  (.A1(\V1/A3/A1/A1/M2/s1 ),
    .A2(\V1/A3/A1/A1/c1 ),
    .ZN(\V1/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M2/M2/_1_  (.A(\V1/A3/A1/A1/M2/s1 ),
    .B(\V1/A3/A1/A1/c1 ),
    .Z(v1[17]));
 OR2_X1 \V1/A3/A1/A1/M2/_0_  (.A1(\V1/A3/A1/A1/M2/c1 ),
    .A2(\V1/A3/A1/A1/M2/c2 ),
    .ZN(\V1/A3/A1/A1/c2 ));
 AND2_X1 \V1/A3/A1/A1/M3/M1/_0_  (.A1(\V1/v4 [2]),
    .A2(\V1/s2 [10]),
    .ZN(\V1/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M3/M1/_1_  (.A(\V1/v4 [2]),
    .B(\V1/s2 [10]),
    .Z(\V1/A3/A1/A1/M3/s1 ));
 AND2_X1 \V1/A3/A1/A1/M3/M2/_0_  (.A1(\V1/A3/A1/A1/M3/s1 ),
    .A2(\V1/A3/A1/A1/c2 ),
    .ZN(\V1/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M3/M2/_1_  (.A(\V1/A3/A1/A1/M3/s1 ),
    .B(\V1/A3/A1/A1/c2 ),
    .Z(v1[18]));
 OR2_X1 \V1/A3/A1/A1/M3/_0_  (.A1(\V1/A3/A1/A1/M3/c1 ),
    .A2(\V1/A3/A1/A1/M3/c2 ),
    .ZN(\V1/A3/A1/A1/c3 ));
 AND2_X1 \V1/A3/A1/A1/M4/M1/_0_  (.A1(\V1/v4 [3]),
    .A2(\V1/s2 [11]),
    .ZN(\V1/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M4/M1/_1_  (.A(\V1/v4 [3]),
    .B(\V1/s2 [11]),
    .Z(\V1/A3/A1/A1/M4/s1 ));
 AND2_X1 \V1/A3/A1/A1/M4/M2/_0_  (.A1(\V1/A3/A1/A1/M4/s1 ),
    .A2(\V1/A3/A1/A1/c3 ),
    .ZN(\V1/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M4/M2/_1_  (.A(\V1/A3/A1/A1/M4/s1 ),
    .B(\V1/A3/A1/A1/c3 ),
    .Z(v1[19]));
 OR2_X1 \V1/A3/A1/A1/M4/_0_  (.A1(\V1/A3/A1/A1/M4/c1 ),
    .A2(\V1/A3/A1/A1/M4/c2 ),
    .ZN(\V1/A3/A1/c1 ));
 AND2_X1 \V1/A3/A1/A2/M1/M1/_0_  (.A1(\V1/v4 [4]),
    .A2(\V1/s2 [12]),
    .ZN(\V1/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M1/M1/_1_  (.A(\V1/v4 [4]),
    .B(\V1/s2 [12]),
    .Z(\V1/A3/A1/A2/M1/s1 ));
 AND2_X1 \V1/A3/A1/A2/M1/M2/_0_  (.A1(\V1/A3/A1/A2/M1/s1 ),
    .A2(\V1/A3/A1/c1 ),
    .ZN(\V1/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M1/M2/_1_  (.A(\V1/A3/A1/A2/M1/s1 ),
    .B(\V1/A3/A1/c1 ),
    .Z(v1[20]));
 OR2_X1 \V1/A3/A1/A2/M1/_0_  (.A1(\V1/A3/A1/A2/M1/c1 ),
    .A2(\V1/A3/A1/A2/M1/c2 ),
    .ZN(\V1/A3/A1/A2/c1 ));
 AND2_X1 \V1/A3/A1/A2/M2/M1/_0_  (.A1(\V1/v4 [5]),
    .A2(\V1/s2 [13]),
    .ZN(\V1/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M2/M1/_1_  (.A(\V1/v4 [5]),
    .B(\V1/s2 [13]),
    .Z(\V1/A3/A1/A2/M2/s1 ));
 AND2_X1 \V1/A3/A1/A2/M2/M2/_0_  (.A1(\V1/A3/A1/A2/M2/s1 ),
    .A2(\V1/A3/A1/A2/c1 ),
    .ZN(\V1/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M2/M2/_1_  (.A(\V1/A3/A1/A2/M2/s1 ),
    .B(\V1/A3/A1/A2/c1 ),
    .Z(v1[21]));
 OR2_X1 \V1/A3/A1/A2/M2/_0_  (.A1(\V1/A3/A1/A2/M2/c1 ),
    .A2(\V1/A3/A1/A2/M2/c2 ),
    .ZN(\V1/A3/A1/A2/c2 ));
 AND2_X1 \V1/A3/A1/A2/M3/M1/_0_  (.A1(\V1/v4 [6]),
    .A2(\V1/s2 [14]),
    .ZN(\V1/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M3/M1/_1_  (.A(\V1/v4 [6]),
    .B(\V1/s2 [14]),
    .Z(\V1/A3/A1/A2/M3/s1 ));
 AND2_X1 \V1/A3/A1/A2/M3/M2/_0_  (.A1(\V1/A3/A1/A2/M3/s1 ),
    .A2(\V1/A3/A1/A2/c2 ),
    .ZN(\V1/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M3/M2/_1_  (.A(\V1/A3/A1/A2/M3/s1 ),
    .B(\V1/A3/A1/A2/c2 ),
    .Z(v1[22]));
 OR2_X1 \V1/A3/A1/A2/M3/_0_  (.A1(\V1/A3/A1/A2/M3/c1 ),
    .A2(\V1/A3/A1/A2/M3/c2 ),
    .ZN(\V1/A3/A1/A2/c3 ));
 AND2_X1 \V1/A3/A1/A2/M4/M1/_0_  (.A1(\V1/v4 [7]),
    .A2(\V1/s2 [15]),
    .ZN(\V1/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M4/M1/_1_  (.A(\V1/v4 [7]),
    .B(\V1/s2 [15]),
    .Z(\V1/A3/A1/A2/M4/s1 ));
 AND2_X1 \V1/A3/A1/A2/M4/M2/_0_  (.A1(\V1/A3/A1/A2/M4/s1 ),
    .A2(\V1/A3/A1/A2/c3 ),
    .ZN(\V1/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M4/M2/_1_  (.A(\V1/A3/A1/A2/M4/s1 ),
    .B(\V1/A3/A1/A2/c3 ),
    .Z(v1[23]));
 OR2_X1 \V1/A3/A1/A2/M4/_0_  (.A1(\V1/A3/A1/A2/M4/c1 ),
    .A2(\V1/A3/A1/A2/M4/c2 ),
    .ZN(\V1/A3/c1 ));
 AND2_X1 \V1/A3/A2/A1/M1/M1/_0_  (.A1(\V1/v4 [8]),
    .A2(\V1/c3 ),
    .ZN(\V1/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M1/M1/_1_  (.A(\V1/v4 [8]),
    .B(\V1/c3 ),
    .Z(\V1/A3/A2/A1/M1/s1 ));
 AND2_X1 \V1/A3/A2/A1/M1/M2/_0_  (.A1(\V1/A3/A2/A1/M1/s1 ),
    .A2(\V1/A3/c1 ),
    .ZN(\V1/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M1/M2/_1_  (.A(\V1/A3/A2/A1/M1/s1 ),
    .B(\V1/A3/c1 ),
    .Z(v1[24]));
 OR2_X1 \V1/A3/A2/A1/M1/_0_  (.A1(\V1/A3/A2/A1/M1/c1 ),
    .A2(\V1/A3/A2/A1/M1/c2 ),
    .ZN(\V1/A3/A2/A1/c1 ));
 AND2_X1 \V1/A3/A2/A1/M2/M1/_0_  (.A1(\V1/v4 [9]),
    .A2(ground),
    .ZN(\V1/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M2/M1/_1_  (.A(\V1/v4 [9]),
    .B(ground),
    .Z(\V1/A3/A2/A1/M2/s1 ));
 AND2_X1 \V1/A3/A2/A1/M2/M2/_0_  (.A1(\V1/A3/A2/A1/M2/s1 ),
    .A2(\V1/A3/A2/A1/c1 ),
    .ZN(\V1/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M2/M2/_1_  (.A(\V1/A3/A2/A1/M2/s1 ),
    .B(\V1/A3/A2/A1/c1 ),
    .Z(v1[25]));
 OR2_X1 \V1/A3/A2/A1/M2/_0_  (.A1(\V1/A3/A2/A1/M2/c1 ),
    .A2(\V1/A3/A2/A1/M2/c2 ),
    .ZN(\V1/A3/A2/A1/c2 ));
 AND2_X1 \V1/A3/A2/A1/M3/M1/_0_  (.A1(\V1/v4 [10]),
    .A2(ground),
    .ZN(\V1/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M3/M1/_1_  (.A(\V1/v4 [10]),
    .B(ground),
    .Z(\V1/A3/A2/A1/M3/s1 ));
 AND2_X1 \V1/A3/A2/A1/M3/M2/_0_  (.A1(\V1/A3/A2/A1/M3/s1 ),
    .A2(\V1/A3/A2/A1/c2 ),
    .ZN(\V1/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M3/M2/_1_  (.A(\V1/A3/A2/A1/M3/s1 ),
    .B(\V1/A3/A2/A1/c2 ),
    .Z(v1[26]));
 OR2_X1 \V1/A3/A2/A1/M3/_0_  (.A1(\V1/A3/A2/A1/M3/c1 ),
    .A2(\V1/A3/A2/A1/M3/c2 ),
    .ZN(\V1/A3/A2/A1/c3 ));
 AND2_X1 \V1/A3/A2/A1/M4/M1/_0_  (.A1(\V1/v4 [11]),
    .A2(ground),
    .ZN(\V1/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M4/M1/_1_  (.A(\V1/v4 [11]),
    .B(ground),
    .Z(\V1/A3/A2/A1/M4/s1 ));
 AND2_X1 \V1/A3/A2/A1/M4/M2/_0_  (.A1(\V1/A3/A2/A1/M4/s1 ),
    .A2(\V1/A3/A2/A1/c3 ),
    .ZN(\V1/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M4/M2/_1_  (.A(\V1/A3/A2/A1/M4/s1 ),
    .B(\V1/A3/A2/A1/c3 ),
    .Z(v1[27]));
 OR2_X1 \V1/A3/A2/A1/M4/_0_  (.A1(\V1/A3/A2/A1/M4/c1 ),
    .A2(\V1/A3/A2/A1/M4/c2 ),
    .ZN(\V1/A3/A2/c1 ));
 AND2_X1 \V1/A3/A2/A2/M1/M1/_0_  (.A1(\V1/v4 [12]),
    .A2(ground),
    .ZN(\V1/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M1/M1/_1_  (.A(\V1/v4 [12]),
    .B(ground),
    .Z(\V1/A3/A2/A2/M1/s1 ));
 AND2_X1 \V1/A3/A2/A2/M1/M2/_0_  (.A1(\V1/A3/A2/A2/M1/s1 ),
    .A2(\V1/A3/A2/c1 ),
    .ZN(\V1/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M1/M2/_1_  (.A(\V1/A3/A2/A2/M1/s1 ),
    .B(\V1/A3/A2/c1 ),
    .Z(v1[28]));
 OR2_X1 \V1/A3/A2/A2/M1/_0_  (.A1(\V1/A3/A2/A2/M1/c1 ),
    .A2(\V1/A3/A2/A2/M1/c2 ),
    .ZN(\V1/A3/A2/A2/c1 ));
 AND2_X1 \V1/A3/A2/A2/M2/M1/_0_  (.A1(\V1/v4 [13]),
    .A2(ground),
    .ZN(\V1/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M2/M1/_1_  (.A(\V1/v4 [13]),
    .B(ground),
    .Z(\V1/A3/A2/A2/M2/s1 ));
 AND2_X1 \V1/A3/A2/A2/M2/M2/_0_  (.A1(\V1/A3/A2/A2/M2/s1 ),
    .A2(\V1/A3/A2/A2/c1 ),
    .ZN(\V1/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M2/M2/_1_  (.A(\V1/A3/A2/A2/M2/s1 ),
    .B(\V1/A3/A2/A2/c1 ),
    .Z(v1[29]));
 OR2_X1 \V1/A3/A2/A2/M2/_0_  (.A1(\V1/A3/A2/A2/M2/c1 ),
    .A2(\V1/A3/A2/A2/M2/c2 ),
    .ZN(\V1/A3/A2/A2/c2 ));
 AND2_X1 \V1/A3/A2/A2/M3/M1/_0_  (.A1(\V1/v4 [14]),
    .A2(ground),
    .ZN(\V1/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M3/M1/_1_  (.A(\V1/v4 [14]),
    .B(ground),
    .Z(\V1/A3/A2/A2/M3/s1 ));
 AND2_X1 \V1/A3/A2/A2/M3/M2/_0_  (.A1(\V1/A3/A2/A2/M3/s1 ),
    .A2(\V1/A3/A2/A2/c2 ),
    .ZN(\V1/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M3/M2/_1_  (.A(\V1/A3/A2/A2/M3/s1 ),
    .B(\V1/A3/A2/A2/c2 ),
    .Z(v1[30]));
 OR2_X1 \V1/A3/A2/A2/M3/_0_  (.A1(\V1/A3/A2/A2/M3/c1 ),
    .A2(\V1/A3/A2/A2/M3/c2 ),
    .ZN(\V1/A3/A2/A2/c3 ));
 AND2_X1 \V1/A3/A2/A2/M4/M1/_0_  (.A1(\V1/v4 [15]),
    .A2(ground),
    .ZN(\V1/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M4/M1/_1_  (.A(\V1/v4 [15]),
    .B(ground),
    .Z(\V1/A3/A2/A2/M4/s1 ));
 AND2_X1 \V1/A3/A2/A2/M4/M2/_0_  (.A1(\V1/A3/A2/A2/M4/s1 ),
    .A2(\V1/A3/A2/A2/c3 ),
    .ZN(\V1/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M4/M2/_1_  (.A(\V1/A3/A2/A2/M4/s1 ),
    .B(\V1/A3/A2/A2/c3 ),
    .Z(v1[31]));
 OR2_X1 \V1/A3/A2/A2/M4/_0_  (.A1(\V1/A3/A2/A2/M4/c1 ),
    .A2(\V1/A3/A2/A2/M4/c2 ),
    .ZN(\V1/overflow ));
 AND2_X1 \V1/V1/A1/A1/M1/M1/_0_  (.A1(\V1/V1/v2 [0]),
    .A2(\V1/V1/v3 [0]),
    .ZN(\V1/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M1/M1/_1_  (.A(\V1/V1/v2 [0]),
    .B(\V1/V1/v3 [0]),
    .Z(\V1/V1/A1/A1/M1/s1 ));
 AND2_X1 \V1/V1/A1/A1/M1/M2/_0_  (.A1(\V1/V1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M1/M2/_1_  (.A(\V1/V1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/s1 [0]));
 OR2_X1 \V1/V1/A1/A1/M1/_0_  (.A1(\V1/V1/A1/A1/M1/c1 ),
    .A2(\V1/V1/A1/A1/M1/c2 ),
    .ZN(\V1/V1/A1/A1/c1 ));
 AND2_X1 \V1/V1/A1/A1/M2/M1/_0_  (.A1(\V1/V1/v2 [1]),
    .A2(\V1/V1/v3 [1]),
    .ZN(\V1/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M2/M1/_1_  (.A(\V1/V1/v2 [1]),
    .B(\V1/V1/v3 [1]),
    .Z(\V1/V1/A1/A1/M2/s1 ));
 AND2_X1 \V1/V1/A1/A1/M2/M2/_0_  (.A1(\V1/V1/A1/A1/M2/s1 ),
    .A2(\V1/V1/A1/A1/c1 ),
    .ZN(\V1/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M2/M2/_1_  (.A(\V1/V1/A1/A1/M2/s1 ),
    .B(\V1/V1/A1/A1/c1 ),
    .Z(\V1/V1/s1 [1]));
 OR2_X1 \V1/V1/A1/A1/M2/_0_  (.A1(\V1/V1/A1/A1/M2/c1 ),
    .A2(\V1/V1/A1/A1/M2/c2 ),
    .ZN(\V1/V1/A1/A1/c2 ));
 AND2_X1 \V1/V1/A1/A1/M3/M1/_0_  (.A1(\V1/V1/v2 [2]),
    .A2(\V1/V1/v3 [2]),
    .ZN(\V1/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M3/M1/_1_  (.A(\V1/V1/v2 [2]),
    .B(\V1/V1/v3 [2]),
    .Z(\V1/V1/A1/A1/M3/s1 ));
 AND2_X1 \V1/V1/A1/A1/M3/M2/_0_  (.A1(\V1/V1/A1/A1/M3/s1 ),
    .A2(\V1/V1/A1/A1/c2 ),
    .ZN(\V1/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M3/M2/_1_  (.A(\V1/V1/A1/A1/M3/s1 ),
    .B(\V1/V1/A1/A1/c2 ),
    .Z(\V1/V1/s1 [2]));
 OR2_X1 \V1/V1/A1/A1/M3/_0_  (.A1(\V1/V1/A1/A1/M3/c1 ),
    .A2(\V1/V1/A1/A1/M3/c2 ),
    .ZN(\V1/V1/A1/A1/c3 ));
 AND2_X1 \V1/V1/A1/A1/M4/M1/_0_  (.A1(\V1/V1/v2 [3]),
    .A2(\V1/V1/v3 [3]),
    .ZN(\V1/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M4/M1/_1_  (.A(\V1/V1/v2 [3]),
    .B(\V1/V1/v3 [3]),
    .Z(\V1/V1/A1/A1/M4/s1 ));
 AND2_X1 \V1/V1/A1/A1/M4/M2/_0_  (.A1(\V1/V1/A1/A1/M4/s1 ),
    .A2(\V1/V1/A1/A1/c3 ),
    .ZN(\V1/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M4/M2/_1_  (.A(\V1/V1/A1/A1/M4/s1 ),
    .B(\V1/V1/A1/A1/c3 ),
    .Z(\V1/V1/s1 [3]));
 OR2_X1 \V1/V1/A1/A1/M4/_0_  (.A1(\V1/V1/A1/A1/M4/c1 ),
    .A2(\V1/V1/A1/A1/M4/c2 ),
    .ZN(\V1/V1/A1/c1 ));
 AND2_X1 \V1/V1/A1/A2/M1/M1/_0_  (.A1(\V1/V1/v2 [4]),
    .A2(\V1/V1/v3 [4]),
    .ZN(\V1/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M1/M1/_1_  (.A(\V1/V1/v2 [4]),
    .B(\V1/V1/v3 [4]),
    .Z(\V1/V1/A1/A2/M1/s1 ));
 AND2_X1 \V1/V1/A1/A2/M1/M2/_0_  (.A1(\V1/V1/A1/A2/M1/s1 ),
    .A2(\V1/V1/A1/c1 ),
    .ZN(\V1/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M1/M2/_1_  (.A(\V1/V1/A1/A2/M1/s1 ),
    .B(\V1/V1/A1/c1 ),
    .Z(\V1/V1/s1 [4]));
 OR2_X1 \V1/V1/A1/A2/M1/_0_  (.A1(\V1/V1/A1/A2/M1/c1 ),
    .A2(\V1/V1/A1/A2/M1/c2 ),
    .ZN(\V1/V1/A1/A2/c1 ));
 AND2_X1 \V1/V1/A1/A2/M2/M1/_0_  (.A1(\V1/V1/v2 [5]),
    .A2(\V1/V1/v3 [5]),
    .ZN(\V1/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M2/M1/_1_  (.A(\V1/V1/v2 [5]),
    .B(\V1/V1/v3 [5]),
    .Z(\V1/V1/A1/A2/M2/s1 ));
 AND2_X1 \V1/V1/A1/A2/M2/M2/_0_  (.A1(\V1/V1/A1/A2/M2/s1 ),
    .A2(\V1/V1/A1/A2/c1 ),
    .ZN(\V1/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M2/M2/_1_  (.A(\V1/V1/A1/A2/M2/s1 ),
    .B(\V1/V1/A1/A2/c1 ),
    .Z(\V1/V1/s1 [5]));
 OR2_X1 \V1/V1/A1/A2/M2/_0_  (.A1(\V1/V1/A1/A2/M2/c1 ),
    .A2(\V1/V1/A1/A2/M2/c2 ),
    .ZN(\V1/V1/A1/A2/c2 ));
 AND2_X1 \V1/V1/A1/A2/M3/M1/_0_  (.A1(\V1/V1/v2 [6]),
    .A2(\V1/V1/v3 [6]),
    .ZN(\V1/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M3/M1/_1_  (.A(\V1/V1/v2 [6]),
    .B(\V1/V1/v3 [6]),
    .Z(\V1/V1/A1/A2/M3/s1 ));
 AND2_X1 \V1/V1/A1/A2/M3/M2/_0_  (.A1(\V1/V1/A1/A2/M3/s1 ),
    .A2(\V1/V1/A1/A2/c2 ),
    .ZN(\V1/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M3/M2/_1_  (.A(\V1/V1/A1/A2/M3/s1 ),
    .B(\V1/V1/A1/A2/c2 ),
    .Z(\V1/V1/s1 [6]));
 OR2_X1 \V1/V1/A1/A2/M3/_0_  (.A1(\V1/V1/A1/A2/M3/c1 ),
    .A2(\V1/V1/A1/A2/M3/c2 ),
    .ZN(\V1/V1/A1/A2/c3 ));
 AND2_X1 \V1/V1/A1/A2/M4/M1/_0_  (.A1(\V1/V1/v2 [7]),
    .A2(\V1/V1/v3 [7]),
    .ZN(\V1/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M4/M1/_1_  (.A(\V1/V1/v2 [7]),
    .B(\V1/V1/v3 [7]),
    .Z(\V1/V1/A1/A2/M4/s1 ));
 AND2_X1 \V1/V1/A1/A2/M4/M2/_0_  (.A1(\V1/V1/A1/A2/M4/s1 ),
    .A2(\V1/V1/A1/A2/c3 ),
    .ZN(\V1/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M4/M2/_1_  (.A(\V1/V1/A1/A2/M4/s1 ),
    .B(\V1/V1/A1/A2/c3 ),
    .Z(\V1/V1/s1 [7]));
 OR2_X1 \V1/V1/A1/A2/M4/_0_  (.A1(\V1/V1/A1/A2/M4/c1 ),
    .A2(\V1/V1/A1/A2/M4/c2 ),
    .ZN(\V1/V1/c1 ));
 AND2_X1 \V1/V1/A2/A1/M1/M1/_0_  (.A1(\V1/V1/s1 [0]),
    .A2(\V1/V1/v1 [4]),
    .ZN(\V1/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M1/M1/_1_  (.A(\V1/V1/s1 [0]),
    .B(\V1/V1/v1 [4]),
    .Z(\V1/V1/A2/A1/M1/s1 ));
 AND2_X1 \V1/V1/A2/A1/M1/M2/_0_  (.A1(\V1/V1/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/A2/A1/M1/c2 ));
 XOR2_X1 \V1/V1/A2/A1/M1/M2/_1_  (.A(\V1/V1/A2/A1/M1/s1 ),
    .B(ground),
    .Z(v1[4]));
 OR2_X1 \V1/V1/A2/A1/M1/_0_  (.A1(\V1/V1/A2/A1/M1/c1 ),
    .A2(\V1/V1/A2/A1/M1/c2 ),
    .ZN(\V1/V1/A2/A1/c1 ));
 AND2_X1 \V1/V1/A2/A1/M2/M1/_0_  (.A1(\V1/V1/s1 [1]),
    .A2(\V1/V1/v1 [5]),
    .ZN(\V1/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M2/M1/_1_  (.A(\V1/V1/s1 [1]),
    .B(\V1/V1/v1 [5]),
    .Z(\V1/V1/A2/A1/M2/s1 ));
 AND2_X1 \V1/V1/A2/A1/M2/M2/_0_  (.A1(\V1/V1/A2/A1/M2/s1 ),
    .A2(\V1/V1/A2/A1/c1 ),
    .ZN(\V1/V1/A2/A1/M2/c2 ));
 XOR2_X1 \V1/V1/A2/A1/M2/M2/_1_  (.A(\V1/V1/A2/A1/M2/s1 ),
    .B(\V1/V1/A2/A1/c1 ),
    .Z(v1[5]));
 OR2_X1 \V1/V1/A2/A1/M2/_0_  (.A1(\V1/V1/A2/A1/M2/c1 ),
    .A2(\V1/V1/A2/A1/M2/c2 ),
    .ZN(\V1/V1/A2/A1/c2 ));
 AND2_X1 \V1/V1/A2/A1/M3/M1/_0_  (.A1(\V1/V1/s1 [2]),
    .A2(\V1/V1/v1 [6]),
    .ZN(\V1/V1/A2/A1/M3/c1 ));
 XOR2_X1 \V1/V1/A2/A1/M3/M1/_1_  (.A(\V1/V1/s1 [2]),
    .B(\V1/V1/v1 [6]),
    .Z(\V1/V1/A2/A1/M3/s1 ));
 AND2_X1 \V1/V1/A2/A1/M3/M2/_0_  (.A1(\V1/V1/A2/A1/M3/s1 ),
    .A2(\V1/V1/A2/A1/c2 ),
    .ZN(\V1/V1/A2/A1/M3/c2 ));
 XOR2_X1 \V1/V1/A2/A1/M3/M2/_1_  (.A(\V1/V1/A2/A1/M3/s1 ),
    .B(\V1/V1/A2/A1/c2 ),
    .Z(v1[6]));
 OR2_X1 \V1/V1/A2/A1/M3/_0_  (.A1(\V1/V1/A2/A1/M3/c1 ),
    .A2(\V1/V1/A2/A1/M3/c2 ),
    .ZN(\V1/V1/A2/A1/c3 ));
 AND2_X1 \V1/V1/A2/A1/M4/M1/_0_  (.A1(\V1/V1/s1 [3]),
    .A2(\V1/V1/v1 [7]),
    .ZN(\V1/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M4/M1/_1_  (.A(\V1/V1/s1 [3]),
    .B(\V1/V1/v1 [7]),
    .Z(\V1/V1/A2/A1/M4/s1 ));
 AND2_X1 \V1/V1/A2/A1/M4/M2/_0_  (.A1(\V1/V1/A2/A1/M4/s1 ),
    .A2(\V1/V1/A2/A1/c3 ),
    .ZN(\V1/V1/A2/A1/M4/c2 ));
 XOR2_X1 \V1/V1/A2/A1/M4/M2/_1_  (.A(\V1/V1/A2/A1/M4/s1 ),
    .B(\V1/V1/A2/A1/c3 ),
    .Z(v1[7]));
 OR2_X1 \V1/V1/A2/A1/M4/_0_  (.A1(\V1/V1/A2/A1/M4/c1 ),
    .A2(\V1/V1/A2/A1/M4/c2 ),
    .ZN(\V1/V1/A2/c1 ));
 AND2_X1 \V1/V1/A2/A2/M1/M1/_0_  (.A1(\V1/V1/s1 [4]),
    .A2(ground),
    .ZN(\V1/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M1/M1/_1_  (.A(\V1/V1/s1 [4]),
    .B(ground),
    .Z(\V1/V1/A2/A2/M1/s1 ));
 AND2_X1 \V1/V1/A2/A2/M1/M2/_0_  (.A1(\V1/V1/A2/A2/M1/s1 ),
    .A2(\V1/V1/A2/c1 ),
    .ZN(\V1/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M1/M2/_1_  (.A(\V1/V1/A2/A2/M1/s1 ),
    .B(\V1/V1/A2/c1 ),
    .Z(\V1/V1/s2 [4]));
 OR2_X1 \V1/V1/A2/A2/M1/_0_  (.A1(\V1/V1/A2/A2/M1/c1 ),
    .A2(\V1/V1/A2/A2/M1/c2 ),
    .ZN(\V1/V1/A2/A2/c1 ));
 AND2_X1 \V1/V1/A2/A2/M2/M1/_0_  (.A1(\V1/V1/s1 [5]),
    .A2(ground),
    .ZN(\V1/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M2/M1/_1_  (.A(\V1/V1/s1 [5]),
    .B(ground),
    .Z(\V1/V1/A2/A2/M2/s1 ));
 AND2_X1 \V1/V1/A2/A2/M2/M2/_0_  (.A1(\V1/V1/A2/A2/M2/s1 ),
    .A2(\V1/V1/A2/A2/c1 ),
    .ZN(\V1/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M2/M2/_1_  (.A(\V1/V1/A2/A2/M2/s1 ),
    .B(\V1/V1/A2/A2/c1 ),
    .Z(\V1/V1/s2 [5]));
 OR2_X1 \V1/V1/A2/A2/M2/_0_  (.A1(\V1/V1/A2/A2/M2/c1 ),
    .A2(\V1/V1/A2/A2/M2/c2 ),
    .ZN(\V1/V1/A2/A2/c2 ));
 AND2_X1 \V1/V1/A2/A2/M3/M1/_0_  (.A1(\V1/V1/s1 [6]),
    .A2(ground),
    .ZN(\V1/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M3/M1/_1_  (.A(\V1/V1/s1 [6]),
    .B(ground),
    .Z(\V1/V1/A2/A2/M3/s1 ));
 AND2_X1 \V1/V1/A2/A2/M3/M2/_0_  (.A1(\V1/V1/A2/A2/M3/s1 ),
    .A2(\V1/V1/A2/A2/c2 ),
    .ZN(\V1/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M3/M2/_1_  (.A(\V1/V1/A2/A2/M3/s1 ),
    .B(\V1/V1/A2/A2/c2 ),
    .Z(\V1/V1/s2 [6]));
 OR2_X1 \V1/V1/A2/A2/M3/_0_  (.A1(\V1/V1/A2/A2/M3/c1 ),
    .A2(\V1/V1/A2/A2/M3/c2 ),
    .ZN(\V1/V1/A2/A2/c3 ));
 AND2_X1 \V1/V1/A2/A2/M4/M1/_0_  (.A1(\V1/V1/s1 [7]),
    .A2(ground),
    .ZN(\V1/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M4/M1/_1_  (.A(\V1/V1/s1 [7]),
    .B(ground),
    .Z(\V1/V1/A2/A2/M4/s1 ));
 AND2_X1 \V1/V1/A2/A2/M4/M2/_0_  (.A1(\V1/V1/A2/A2/M4/s1 ),
    .A2(\V1/V1/A2/A2/c3 ),
    .ZN(\V1/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M4/M2/_1_  (.A(\V1/V1/A2/A2/M4/s1 ),
    .B(\V1/V1/A2/A2/c3 ),
    .Z(\V1/V1/s2 [7]));
 OR2_X1 \V1/V1/A2/A2/M4/_0_  (.A1(\V1/V1/A2/A2/M4/c1 ),
    .A2(\V1/V1/A2/A2/M4/c2 ),
    .ZN(\V1/V1/c2 ));
 AND2_X1 \V1/V1/A3/A1/M1/M1/_0_  (.A1(\V1/V1/v4 [0]),
    .A2(\V1/V1/s2 [4]),
    .ZN(\V1/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M1/M1/_1_  (.A(\V1/V1/v4 [0]),
    .B(\V1/V1/s2 [4]),
    .Z(\V1/V1/A3/A1/M1/s1 ));
 AND2_X1 \V1/V1/A3/A1/M1/M2/_0_  (.A1(\V1/V1/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M1/M2/_1_  (.A(\V1/V1/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v1 [8]));
 OR2_X1 \V1/V1/A3/A1/M1/_0_  (.A1(\V1/V1/A3/A1/M1/c1 ),
    .A2(\V1/V1/A3/A1/M1/c2 ),
    .ZN(\V1/V1/A3/A1/c1 ));
 AND2_X1 \V1/V1/A3/A1/M2/M1/_0_  (.A1(\V1/V1/v4 [1]),
    .A2(\V1/V1/s2 [5]),
    .ZN(\V1/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M2/M1/_1_  (.A(\V1/V1/v4 [1]),
    .B(\V1/V1/s2 [5]),
    .Z(\V1/V1/A3/A1/M2/s1 ));
 AND2_X1 \V1/V1/A3/A1/M2/M2/_0_  (.A1(\V1/V1/A3/A1/M2/s1 ),
    .A2(\V1/V1/A3/A1/c1 ),
    .ZN(\V1/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M2/M2/_1_  (.A(\V1/V1/A3/A1/M2/s1 ),
    .B(\V1/V1/A3/A1/c1 ),
    .Z(\V1/v1 [9]));
 OR2_X1 \V1/V1/A3/A1/M2/_0_  (.A1(\V1/V1/A3/A1/M2/c1 ),
    .A2(\V1/V1/A3/A1/M2/c2 ),
    .ZN(\V1/V1/A3/A1/c2 ));
 AND2_X1 \V1/V1/A3/A1/M3/M1/_0_  (.A1(\V1/V1/v4 [2]),
    .A2(\V1/V1/s2 [6]),
    .ZN(\V1/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M3/M1/_1_  (.A(\V1/V1/v4 [2]),
    .B(\V1/V1/s2 [6]),
    .Z(\V1/V1/A3/A1/M3/s1 ));
 AND2_X1 \V1/V1/A3/A1/M3/M2/_0_  (.A1(\V1/V1/A3/A1/M3/s1 ),
    .A2(\V1/V1/A3/A1/c2 ),
    .ZN(\V1/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M3/M2/_1_  (.A(\V1/V1/A3/A1/M3/s1 ),
    .B(\V1/V1/A3/A1/c2 ),
    .Z(\V1/v1 [10]));
 OR2_X1 \V1/V1/A3/A1/M3/_0_  (.A1(\V1/V1/A3/A1/M3/c1 ),
    .A2(\V1/V1/A3/A1/M3/c2 ),
    .ZN(\V1/V1/A3/A1/c3 ));
 AND2_X1 \V1/V1/A3/A1/M4/M1/_0_  (.A1(\V1/V1/v4 [3]),
    .A2(\V1/V1/s2 [7]),
    .ZN(\V1/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M4/M1/_1_  (.A(\V1/V1/v4 [3]),
    .B(\V1/V1/s2 [7]),
    .Z(\V1/V1/A3/A1/M4/s1 ));
 AND2_X1 \V1/V1/A3/A1/M4/M2/_0_  (.A1(\V1/V1/A3/A1/M4/s1 ),
    .A2(\V1/V1/A3/A1/c3 ),
    .ZN(\V1/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M4/M2/_1_  (.A(\V1/V1/A3/A1/M4/s1 ),
    .B(\V1/V1/A3/A1/c3 ),
    .Z(\V1/v1 [11]));
 OR2_X1 \V1/V1/A3/A1/M4/_0_  (.A1(\V1/V1/A3/A1/M4/c1 ),
    .A2(\V1/V1/A3/A1/M4/c2 ),
    .ZN(\V1/V1/A3/c1 ));
 AND2_X1 \V1/V1/A3/A2/M1/M1/_0_  (.A1(\V1/V1/v4 [4]),
    .A2(\V1/V1/c3 ),
    .ZN(\V1/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M1/M1/_1_  (.A(\V1/V1/v4 [4]),
    .B(\V1/V1/c3 ),
    .Z(\V1/V1/A3/A2/M1/s1 ));
 AND2_X1 \V1/V1/A3/A2/M1/M2/_0_  (.A1(\V1/V1/A3/A2/M1/s1 ),
    .A2(\V1/V1/A3/c1 ),
    .ZN(\V1/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M1/M2/_1_  (.A(\V1/V1/A3/A2/M1/s1 ),
    .B(\V1/V1/A3/c1 ),
    .Z(\V1/v1 [12]));
 OR2_X1 \V1/V1/A3/A2/M1/_0_  (.A1(\V1/V1/A3/A2/M1/c1 ),
    .A2(\V1/V1/A3/A2/M1/c2 ),
    .ZN(\V1/V1/A3/A2/c1 ));
 AND2_X1 \V1/V1/A3/A2/M2/M1/_0_  (.A1(\V1/V1/v4 [5]),
    .A2(ground),
    .ZN(\V1/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M2/M1/_1_  (.A(\V1/V1/v4 [5]),
    .B(ground),
    .Z(\V1/V1/A3/A2/M2/s1 ));
 AND2_X1 \V1/V1/A3/A2/M2/M2/_0_  (.A1(\V1/V1/A3/A2/M2/s1 ),
    .A2(\V1/V1/A3/A2/c1 ),
    .ZN(\V1/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M2/M2/_1_  (.A(\V1/V1/A3/A2/M2/s1 ),
    .B(\V1/V1/A3/A2/c1 ),
    .Z(\V1/v1 [13]));
 OR2_X1 \V1/V1/A3/A2/M2/_0_  (.A1(\V1/V1/A3/A2/M2/c1 ),
    .A2(\V1/V1/A3/A2/M2/c2 ),
    .ZN(\V1/V1/A3/A2/c2 ));
 AND2_X1 \V1/V1/A3/A2/M3/M1/_0_  (.A1(\V1/V1/v4 [6]),
    .A2(ground),
    .ZN(\V1/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M3/M1/_1_  (.A(\V1/V1/v4 [6]),
    .B(ground),
    .Z(\V1/V1/A3/A2/M3/s1 ));
 AND2_X1 \V1/V1/A3/A2/M3/M2/_0_  (.A1(\V1/V1/A3/A2/M3/s1 ),
    .A2(\V1/V1/A3/A2/c2 ),
    .ZN(\V1/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M3/M2/_1_  (.A(\V1/V1/A3/A2/M3/s1 ),
    .B(\V1/V1/A3/A2/c2 ),
    .Z(\V1/v1 [14]));
 OR2_X1 \V1/V1/A3/A2/M3/_0_  (.A1(\V1/V1/A3/A2/M3/c1 ),
    .A2(\V1/V1/A3/A2/M3/c2 ),
    .ZN(\V1/V1/A3/A2/c3 ));
 AND2_X1 \V1/V1/A3/A2/M4/M1/_0_  (.A1(\V1/V1/v4 [7]),
    .A2(ground),
    .ZN(\V1/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M4/M1/_1_  (.A(\V1/V1/v4 [7]),
    .B(ground),
    .Z(\V1/V1/A3/A2/M4/s1 ));
 AND2_X1 \V1/V1/A3/A2/M4/M2/_0_  (.A1(\V1/V1/A3/A2/M4/s1 ),
    .A2(\V1/V1/A3/A2/c3 ),
    .ZN(\V1/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M4/M2/_1_  (.A(\V1/V1/A3/A2/M4/s1 ),
    .B(\V1/V1/A3/A2/c3 ),
    .Z(\V1/v1 [15]));
 OR2_X1 \V1/V1/A3/A2/M4/_0_  (.A1(\V1/V1/A3/A2/M4/c1 ),
    .A2(\V1/V1/A3/A2/M4/c2 ),
    .ZN(\V1/V1/overflow ));
 AND2_X1 \V1/V1/V1/A1/M1/M1/_0_  (.A1(\V1/V1/V1/v2 [0]),
    .A2(\V1/V1/V1/v3 [0]),
    .ZN(\V1/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M1/M1/_1_  (.A(\V1/V1/V1/v2 [0]),
    .B(\V1/V1/V1/v3 [0]),
    .Z(\V1/V1/V1/A1/M1/s1 ));
 AND2_X1 \V1/V1/V1/A1/M1/M2/_0_  (.A1(\V1/V1/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M1/M2/_1_  (.A(\V1/V1/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/V1/s1 [0]));
 OR2_X1 \V1/V1/V1/A1/M1/_0_  (.A1(\V1/V1/V1/A1/M1/c1 ),
    .A2(\V1/V1/V1/A1/M1/c2 ),
    .ZN(\V1/V1/V1/A1/c1 ));
 AND2_X1 \V1/V1/V1/A1/M2/M1/_0_  (.A1(\V1/V1/V1/v2 [1]),
    .A2(\V1/V1/V1/v3 [1]),
    .ZN(\V1/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M2/M1/_1_  (.A(\V1/V1/V1/v2 [1]),
    .B(\V1/V1/V1/v3 [1]),
    .Z(\V1/V1/V1/A1/M2/s1 ));
 AND2_X2 \V1/V1/V1/A1/M2/M2/_0_  (.A1(\V1/V1/V1/A1/M2/s1 ),
    .A2(\V1/V1/V1/A1/c1 ),
    .ZN(\V1/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M2/M2/_1_  (.A(\V1/V1/V1/A1/M2/s1 ),
    .B(\V1/V1/V1/A1/c1 ),
    .Z(\V1/V1/V1/s1 [1]));
 OR2_X1 \V1/V1/V1/A1/M2/_0_  (.A1(\V1/V1/V1/A1/M2/c1 ),
    .A2(\V1/V1/V1/A1/M2/c2 ),
    .ZN(\V1/V1/V1/A1/c2 ));
 AND2_X1 \V1/V1/V1/A1/M3/M1/_0_  (.A1(\V1/V1/V1/v2 [2]),
    .A2(\V1/V1/V1/v3 [2]),
    .ZN(\V1/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M3/M1/_1_  (.A(\V1/V1/V1/v2 [2]),
    .B(\V1/V1/V1/v3 [2]),
    .Z(\V1/V1/V1/A1/M3/s1 ));
 AND2_X1 \V1/V1/V1/A1/M3/M2/_0_  (.A1(\V1/V1/V1/A1/M3/s1 ),
    .A2(\V1/V1/V1/A1/c2 ),
    .ZN(\V1/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M3/M2/_1_  (.A(\V1/V1/V1/A1/M3/s1 ),
    .B(\V1/V1/V1/A1/c2 ),
    .Z(\V1/V1/V1/s1 [2]));
 OR2_X1 \V1/V1/V1/A1/M3/_0_  (.A1(\V1/V1/V1/A1/M3/c1 ),
    .A2(\V1/V1/V1/A1/M3/c2 ),
    .ZN(\V1/V1/V1/A1/c3 ));
 AND2_X1 \V1/V1/V1/A1/M4/M1/_0_  (.A1(\V1/V1/V1/v2 [3]),
    .A2(\V1/V1/V1/v3 [3]),
    .ZN(\V1/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M4/M1/_1_  (.A(\V1/V1/V1/v2 [3]),
    .B(\V1/V1/V1/v3 [3]),
    .Z(\V1/V1/V1/A1/M4/s1 ));
 AND2_X1 \V1/V1/V1/A1/M4/M2/_0_  (.A1(\V1/V1/V1/A1/M4/s1 ),
    .A2(\V1/V1/V1/A1/c3 ),
    .ZN(\V1/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M4/M2/_1_  (.A(\V1/V1/V1/A1/M4/s1 ),
    .B(\V1/V1/V1/A1/c3 ),
    .Z(\V1/V1/V1/s1 [3]));
 OR2_X1 \V1/V1/V1/A1/M4/_0_  (.A1(\V1/V1/V1/A1/M4/c1 ),
    .A2(\V1/V1/V1/A1/M4/c2 ),
    .ZN(\V1/V1/V1/c1 ));
 AND2_X1 \V1/V1/V1/A2/M1/M1/_0_  (.A1(\V1/V1/V1/s1 [0]),
    .A2(\V1/V1/V1/v1 [2]),
    .ZN(\V1/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M1/M1/_1_  (.A(\V1/V1/V1/s1 [0]),
    .B(\V1/V1/V1/v1 [2]),
    .Z(\V1/V1/V1/A2/M1/s1 ));
 AND2_X1 \V1/V1/V1/A2/M1/M2/_0_  (.A1(\V1/V1/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M1/M2/_1_  (.A(\V1/V1/V1/A2/M1/s1 ),
    .B(ground),
    .Z(v1[2]));
 OR2_X1 \V1/V1/V1/A2/M1/_0_  (.A1(\V1/V1/V1/A2/M1/c1 ),
    .A2(\V1/V1/V1/A2/M1/c2 ),
    .ZN(\V1/V1/V1/A2/c1 ));
 AND2_X1 \V1/V1/V1/A2/M2/M1/_0_  (.A1(\V1/V1/V1/s1 [1]),
    .A2(\V1/V1/V1/v1 [3]),
    .ZN(\V1/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M2/M1/_1_  (.A(\V1/V1/V1/s1 [1]),
    .B(\V1/V1/V1/v1 [3]),
    .Z(\V1/V1/V1/A2/M2/s1 ));
 AND2_X1 \V1/V1/V1/A2/M2/M2/_0_  (.A1(\V1/V1/V1/A2/M2/s1 ),
    .A2(\V1/V1/V1/A2/c1 ),
    .ZN(\V1/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M2/M2/_1_  (.A(\V1/V1/V1/A2/M2/s1 ),
    .B(\V1/V1/V1/A2/c1 ),
    .Z(v1[3]));
 OR2_X2 \V1/V1/V1/A2/M2/_0_  (.A1(\V1/V1/V1/A2/M2/c1 ),
    .A2(\V1/V1/V1/A2/M2/c2 ),
    .ZN(\V1/V1/V1/A2/c2 ));
 AND2_X1 \V1/V1/V1/A2/M3/M1/_0_  (.A1(\V1/V1/V1/s1 [2]),
    .A2(ground),
    .ZN(\V1/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M3/M1/_1_  (.A(\V1/V1/V1/s1 [2]),
    .B(ground),
    .Z(\V1/V1/V1/A2/M3/s1 ));
 AND2_X1 \V1/V1/V1/A2/M3/M2/_0_  (.A1(\V1/V1/V1/A2/M3/s1 ),
    .A2(\V1/V1/V1/A2/c2 ),
    .ZN(\V1/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M3/M2/_1_  (.A(\V1/V1/V1/A2/M3/s1 ),
    .B(\V1/V1/V1/A2/c2 ),
    .Z(\V1/V1/V1/s2 [2]));
 OR2_X1 \V1/V1/V1/A2/M3/_0_  (.A1(\V1/V1/V1/A2/M3/c1 ),
    .A2(\V1/V1/V1/A2/M3/c2 ),
    .ZN(\V1/V1/V1/A2/c3 ));
 AND2_X1 \V1/V1/V1/A2/M4/M1/_0_  (.A1(\V1/V1/V1/s1 [3]),
    .A2(ground),
    .ZN(\V1/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M4/M1/_1_  (.A(\V1/V1/V1/s1 [3]),
    .B(ground),
    .Z(\V1/V1/V1/A2/M4/s1 ));
 AND2_X1 \V1/V1/V1/A2/M4/M2/_0_  (.A1(\V1/V1/V1/A2/M4/s1 ),
    .A2(\V1/V1/V1/A2/c3 ),
    .ZN(\V1/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M4/M2/_1_  (.A(\V1/V1/V1/A2/M4/s1 ),
    .B(\V1/V1/V1/A2/c3 ),
    .Z(\V1/V1/V1/s2 [3]));
 OR2_X1 \V1/V1/V1/A2/M4/_0_  (.A1(\V1/V1/V1/A2/M4/c1 ),
    .A2(\V1/V1/V1/A2/M4/c2 ),
    .ZN(\V1/V1/V1/c2 ));
 AND2_X1 \V1/V1/V1/A3/M1/M1/_0_  (.A1(\V1/V1/V1/v4 [0]),
    .A2(\V1/V1/V1/s2 [2]),
    .ZN(\V1/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M1/M1/_1_  (.A(\V1/V1/V1/v4 [0]),
    .B(\V1/V1/V1/s2 [2]),
    .Z(\V1/V1/V1/A3/M1/s1 ));
 AND2_X1 \V1/V1/V1/A3/M1/M2/_0_  (.A1(\V1/V1/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M1/M2/_1_  (.A(\V1/V1/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v1 [4]));
 OR2_X1 \V1/V1/V1/A3/M1/_0_  (.A1(\V1/V1/V1/A3/M1/c1 ),
    .A2(\V1/V1/V1/A3/M1/c2 ),
    .ZN(\V1/V1/V1/A3/c1 ));
 AND2_X1 \V1/V1/V1/A3/M2/M1/_0_  (.A1(\V1/V1/V1/v4 [1]),
    .A2(\V1/V1/V1/s2 [3]),
    .ZN(\V1/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M2/M1/_1_  (.A(\V1/V1/V1/v4 [1]),
    .B(\V1/V1/V1/s2 [3]),
    .Z(\V1/V1/V1/A3/M2/s1 ));
 AND2_X1 \V1/V1/V1/A3/M2/M2/_0_  (.A1(\V1/V1/V1/A3/M2/s1 ),
    .A2(\V1/V1/V1/A3/c1 ),
    .ZN(\V1/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M2/M2/_1_  (.A(\V1/V1/V1/A3/M2/s1 ),
    .B(\V1/V1/V1/A3/c1 ),
    .Z(\V1/V1/v1 [5]));
 OR2_X1 \V1/V1/V1/A3/M2/_0_  (.A1(\V1/V1/V1/A3/M2/c1 ),
    .A2(\V1/V1/V1/A3/M2/c2 ),
    .ZN(\V1/V1/V1/A3/c2 ));
 AND2_X1 \V1/V1/V1/A3/M3/M1/_0_  (.A1(\V1/V1/V1/v4 [2]),
    .A2(\V1/V1/V1/c3 ),
    .ZN(\V1/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M3/M1/_1_  (.A(\V1/V1/V1/v4 [2]),
    .B(\V1/V1/V1/c3 ),
    .Z(\V1/V1/V1/A3/M3/s1 ));
 AND2_X1 \V1/V1/V1/A3/M3/M2/_0_  (.A1(\V1/V1/V1/A3/M3/s1 ),
    .A2(\V1/V1/V1/A3/c2 ),
    .ZN(\V1/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M3/M2/_1_  (.A(\V1/V1/V1/A3/M3/s1 ),
    .B(\V1/V1/V1/A3/c2 ),
    .Z(\V1/V1/v1 [6]));
 OR2_X1 \V1/V1/V1/A3/M3/_0_  (.A1(\V1/V1/V1/A3/M3/c1 ),
    .A2(\V1/V1/V1/A3/M3/c2 ),
    .ZN(\V1/V1/V1/A3/c3 ));
 AND2_X1 \V1/V1/V1/A3/M4/M1/_0_  (.A1(\V1/V1/V1/v4 [3]),
    .A2(ground),
    .ZN(\V1/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M4/M1/_1_  (.A(\V1/V1/V1/v4 [3]),
    .B(ground),
    .Z(\V1/V1/V1/A3/M4/s1 ));
 AND2_X1 \V1/V1/V1/A3/M4/M2/_0_  (.A1(\V1/V1/V1/A3/M4/s1 ),
    .A2(\V1/V1/V1/A3/c3 ),
    .ZN(\V1/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M4/M2/_1_  (.A(\V1/V1/V1/A3/M4/s1 ),
    .B(\V1/V1/V1/A3/c3 ),
    .Z(\V1/V1/v1 [7]));
 OR2_X1 \V1/V1/V1/A3/M4/_0_  (.A1(\V1/V1/V1/A3/M4/c1 ),
    .A2(\V1/V1/V1/A3/M4/c2 ),
    .ZN(\V1/V1/V1/overflow ));
 AND2_X1 \V1/V1/V1/V1/HA1/_0_  (.A1(\V1/V1/V1/V1/w2 ),
    .A2(\V1/V1/V1/V1/w1 ),
    .ZN(\V1/V1/V1/V1/w4 ));
 XOR2_X2 \V1/V1/V1/V1/HA1/_1_  (.A(\V1/V1/V1/V1/w2 ),
    .B(\V1/V1/V1/V1/w1 ),
    .Z(v1[1]));
 AND2_X1 \V1/V1/V1/V1/HA2/_0_  (.A1(\V1/V1/V1/V1/w4 ),
    .A2(\V1/V1/V1/V1/w3 ),
    .ZN(\V1/V1/V1/v1 [3]));
 XOR2_X2 \V1/V1/V1/V1/HA2/_1_  (.A(\V1/V1/V1/V1/w4 ),
    .B(\V1/V1/V1/V1/w3 ),
    .Z(\V1/V1/V1/v1 [2]));
 AND2_X1 \V1/V1/V1/V1/_0_  (.A1(A[0]),
    .A2(B[0]),
    .ZN(v1[0]));
 AND2_X1 \V1/V1/V1/V1/_1_  (.A1(A[0]),
    .A2(B[1]),
    .ZN(\V1/V1/V1/V1/w1 ));
 AND2_X1 \V1/V1/V1/V1/_2_  (.A1(B[0]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V1/w2 ));
 AND2_X1 \V1/V1/V1/V1/_3_  (.A1(B[1]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V1/w3 ));
 AND2_X1 \V1/V1/V1/V2/HA1/_0_  (.A1(\V1/V1/V1/V2/w2 ),
    .A2(\V1/V1/V1/V2/w1 ),
    .ZN(\V1/V1/V1/V2/w4 ));
 XOR2_X2 \V1/V1/V1/V2/HA1/_1_  (.A(\V1/V1/V1/V2/w2 ),
    .B(\V1/V1/V1/V2/w1 ),
    .Z(\V1/V1/V1/v2 [1]));
 AND2_X1 \V1/V1/V1/V2/HA2/_0_  (.A1(\V1/V1/V1/V2/w4 ),
    .A2(\V1/V1/V1/V2/w3 ),
    .ZN(\V1/V1/V1/v2 [3]));
 XOR2_X2 \V1/V1/V1/V2/HA2/_1_  (.A(\V1/V1/V1/V2/w4 ),
    .B(\V1/V1/V1/V2/w3 ),
    .Z(\V1/V1/V1/v2 [2]));
 AND2_X1 \V1/V1/V1/V2/_0_  (.A1(A[2]),
    .A2(B[0]),
    .ZN(\V1/V1/V1/v2 [0]));
 AND2_X1 \V1/V1/V1/V2/_1_  (.A1(A[2]),
    .A2(B[1]),
    .ZN(\V1/V1/V1/V2/w1 ));
 AND2_X1 \V1/V1/V1/V2/_2_  (.A1(B[0]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V2/w2 ));
 AND2_X1 \V1/V1/V1/V2/_3_  (.A1(B[1]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V2/w3 ));
 AND2_X1 \V1/V1/V1/V3/HA1/_0_  (.A1(\V1/V1/V1/V3/w2 ),
    .A2(\V1/V1/V1/V3/w1 ),
    .ZN(\V1/V1/V1/V3/w4 ));
 XOR2_X2 \V1/V1/V1/V3/HA1/_1_  (.A(\V1/V1/V1/V3/w2 ),
    .B(\V1/V1/V1/V3/w1 ),
    .Z(\V1/V1/V1/v3 [1]));
 AND2_X1 \V1/V1/V1/V3/HA2/_0_  (.A1(\V1/V1/V1/V3/w4 ),
    .A2(\V1/V1/V1/V3/w3 ),
    .ZN(\V1/V1/V1/v3 [3]));
 XOR2_X2 \V1/V1/V1/V3/HA2/_1_  (.A(\V1/V1/V1/V3/w4 ),
    .B(\V1/V1/V1/V3/w3 ),
    .Z(\V1/V1/V1/v3 [2]));
 AND2_X1 \V1/V1/V1/V3/_0_  (.A1(A[0]),
    .A2(B[2]),
    .ZN(\V1/V1/V1/v3 [0]));
 AND2_X1 \V1/V1/V1/V3/_1_  (.A1(A[0]),
    .A2(B[3]),
    .ZN(\V1/V1/V1/V3/w1 ));
 AND2_X1 \V1/V1/V1/V3/_2_  (.A1(B[2]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V3/w2 ));
 AND2_X1 \V1/V1/V1/V3/_3_  (.A1(B[3]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V3/w3 ));
 AND2_X1 \V1/V1/V1/V4/HA1/_0_  (.A1(\V1/V1/V1/V4/w2 ),
    .A2(\V1/V1/V1/V4/w1 ),
    .ZN(\V1/V1/V1/V4/w4 ));
 XOR2_X2 \V1/V1/V1/V4/HA1/_1_  (.A(\V1/V1/V1/V4/w2 ),
    .B(\V1/V1/V1/V4/w1 ),
    .Z(\V1/V1/V1/v4 [1]));
 AND2_X1 \V1/V1/V1/V4/HA2/_0_  (.A1(\V1/V1/V1/V4/w4 ),
    .A2(\V1/V1/V1/V4/w3 ),
    .ZN(\V1/V1/V1/v4 [3]));
 XOR2_X2 \V1/V1/V1/V4/HA2/_1_  (.A(\V1/V1/V1/V4/w4 ),
    .B(\V1/V1/V1/V4/w3 ),
    .Z(\V1/V1/V1/v4 [2]));
 AND2_X1 \V1/V1/V1/V4/_0_  (.A1(A[2]),
    .A2(B[2]),
    .ZN(\V1/V1/V1/v4 [0]));
 AND2_X1 \V1/V1/V1/V4/_1_  (.A1(A[2]),
    .A2(B[3]),
    .ZN(\V1/V1/V1/V4/w1 ));
 AND2_X1 \V1/V1/V1/V4/_2_  (.A1(B[2]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V4/w2 ));
 AND2_X1 \V1/V1/V1/V4/_3_  (.A1(B[3]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V4/w3 ));
 OR2_X1 \V1/V1/V1/_0_  (.A1(\V1/V1/V1/c1 ),
    .A2(\V1/V1/V1/c2 ),
    .ZN(\V1/V1/V1/c3 ));
 AND2_X1 \V1/V1/V2/A1/M1/M1/_0_  (.A1(\V1/V1/V2/v2 [0]),
    .A2(\V1/V1/V2/v3 [0]),
    .ZN(\V1/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M1/M1/_1_  (.A(\V1/V1/V2/v2 [0]),
    .B(\V1/V1/V2/v3 [0]),
    .Z(\V1/V1/V2/A1/M1/s1 ));
 AND2_X1 \V1/V1/V2/A1/M1/M2/_0_  (.A1(\V1/V1/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M1/M2/_1_  (.A(\V1/V1/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/V2/s1 [0]));
 OR2_X1 \V1/V1/V2/A1/M1/_0_  (.A1(\V1/V1/V2/A1/M1/c1 ),
    .A2(\V1/V1/V2/A1/M1/c2 ),
    .ZN(\V1/V1/V2/A1/c1 ));
 AND2_X1 \V1/V1/V2/A1/M2/M1/_0_  (.A1(\V1/V1/V2/v2 [1]),
    .A2(\V1/V1/V2/v3 [1]),
    .ZN(\V1/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M2/M1/_1_  (.A(\V1/V1/V2/v2 [1]),
    .B(\V1/V1/V2/v3 [1]),
    .Z(\V1/V1/V2/A1/M2/s1 ));
 AND2_X1 \V1/V1/V2/A1/M2/M2/_0_  (.A1(\V1/V1/V2/A1/M2/s1 ),
    .A2(\V1/V1/V2/A1/c1 ),
    .ZN(\V1/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M2/M2/_1_  (.A(\V1/V1/V2/A1/M2/s1 ),
    .B(\V1/V1/V2/A1/c1 ),
    .Z(\V1/V1/V2/s1 [1]));
 OR2_X1 \V1/V1/V2/A1/M2/_0_  (.A1(\V1/V1/V2/A1/M2/c1 ),
    .A2(\V1/V1/V2/A1/M2/c2 ),
    .ZN(\V1/V1/V2/A1/c2 ));
 AND2_X1 \V1/V1/V2/A1/M3/M1/_0_  (.A1(\V1/V1/V2/v2 [2]),
    .A2(\V1/V1/V2/v3 [2]),
    .ZN(\V1/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M3/M1/_1_  (.A(\V1/V1/V2/v2 [2]),
    .B(\V1/V1/V2/v3 [2]),
    .Z(\V1/V1/V2/A1/M3/s1 ));
 AND2_X1 \V1/V1/V2/A1/M3/M2/_0_  (.A1(\V1/V1/V2/A1/M3/s1 ),
    .A2(\V1/V1/V2/A1/c2 ),
    .ZN(\V1/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M3/M2/_1_  (.A(\V1/V1/V2/A1/M3/s1 ),
    .B(\V1/V1/V2/A1/c2 ),
    .Z(\V1/V1/V2/s1 [2]));
 OR2_X1 \V1/V1/V2/A1/M3/_0_  (.A1(\V1/V1/V2/A1/M3/c1 ),
    .A2(\V1/V1/V2/A1/M3/c2 ),
    .ZN(\V1/V1/V2/A1/c3 ));
 AND2_X1 \V1/V1/V2/A1/M4/M1/_0_  (.A1(\V1/V1/V2/v2 [3]),
    .A2(\V1/V1/V2/v3 [3]),
    .ZN(\V1/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M4/M1/_1_  (.A(\V1/V1/V2/v2 [3]),
    .B(\V1/V1/V2/v3 [3]),
    .Z(\V1/V1/V2/A1/M4/s1 ));
 AND2_X1 \V1/V1/V2/A1/M4/M2/_0_  (.A1(\V1/V1/V2/A1/M4/s1 ),
    .A2(\V1/V1/V2/A1/c3 ),
    .ZN(\V1/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M4/M2/_1_  (.A(\V1/V1/V2/A1/M4/s1 ),
    .B(\V1/V1/V2/A1/c3 ),
    .Z(\V1/V1/V2/s1 [3]));
 OR2_X1 \V1/V1/V2/A1/M4/_0_  (.A1(\V1/V1/V2/A1/M4/c1 ),
    .A2(\V1/V1/V2/A1/M4/c2 ),
    .ZN(\V1/V1/V2/c1 ));
 AND2_X1 \V1/V1/V2/A2/M1/M1/_0_  (.A1(\V1/V1/V2/s1 [0]),
    .A2(\V1/V1/V2/v1 [2]),
    .ZN(\V1/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M1/M1/_1_  (.A(\V1/V1/V2/s1 [0]),
    .B(\V1/V1/V2/v1 [2]),
    .Z(\V1/V1/V2/A2/M1/s1 ));
 AND2_X1 \V1/V1/V2/A2/M1/M2/_0_  (.A1(\V1/V1/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M1/M2/_1_  (.A(\V1/V1/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v2 [2]));
 OR2_X1 \V1/V1/V2/A2/M1/_0_  (.A1(\V1/V1/V2/A2/M1/c1 ),
    .A2(\V1/V1/V2/A2/M1/c2 ),
    .ZN(\V1/V1/V2/A2/c1 ));
 AND2_X1 \V1/V1/V2/A2/M2/M1/_0_  (.A1(\V1/V1/V2/s1 [1]),
    .A2(\V1/V1/V2/v1 [3]),
    .ZN(\V1/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M2/M1/_1_  (.A(\V1/V1/V2/s1 [1]),
    .B(\V1/V1/V2/v1 [3]),
    .Z(\V1/V1/V2/A2/M2/s1 ));
 AND2_X1 \V1/V1/V2/A2/M2/M2/_0_  (.A1(\V1/V1/V2/A2/M2/s1 ),
    .A2(\V1/V1/V2/A2/c1 ),
    .ZN(\V1/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M2/M2/_1_  (.A(\V1/V1/V2/A2/M2/s1 ),
    .B(\V1/V1/V2/A2/c1 ),
    .Z(\V1/V1/v2 [3]));
 OR2_X1 \V1/V1/V2/A2/M2/_0_  (.A1(\V1/V1/V2/A2/M2/c1 ),
    .A2(\V1/V1/V2/A2/M2/c2 ),
    .ZN(\V1/V1/V2/A2/c2 ));
 AND2_X1 \V1/V1/V2/A2/M3/M1/_0_  (.A1(\V1/V1/V2/s1 [2]),
    .A2(ground),
    .ZN(\V1/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M3/M1/_1_  (.A(\V1/V1/V2/s1 [2]),
    .B(ground),
    .Z(\V1/V1/V2/A2/M3/s1 ));
 AND2_X1 \V1/V1/V2/A2/M3/M2/_0_  (.A1(\V1/V1/V2/A2/M3/s1 ),
    .A2(\V1/V1/V2/A2/c2 ),
    .ZN(\V1/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M3/M2/_1_  (.A(\V1/V1/V2/A2/M3/s1 ),
    .B(\V1/V1/V2/A2/c2 ),
    .Z(\V1/V1/V2/s2 [2]));
 OR2_X1 \V1/V1/V2/A2/M3/_0_  (.A1(\V1/V1/V2/A2/M3/c1 ),
    .A2(\V1/V1/V2/A2/M3/c2 ),
    .ZN(\V1/V1/V2/A2/c3 ));
 AND2_X1 \V1/V1/V2/A2/M4/M1/_0_  (.A1(\V1/V1/V2/s1 [3]),
    .A2(ground),
    .ZN(\V1/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M4/M1/_1_  (.A(\V1/V1/V2/s1 [3]),
    .B(ground),
    .Z(\V1/V1/V2/A2/M4/s1 ));
 AND2_X1 \V1/V1/V2/A2/M4/M2/_0_  (.A1(\V1/V1/V2/A2/M4/s1 ),
    .A2(\V1/V1/V2/A2/c3 ),
    .ZN(\V1/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M4/M2/_1_  (.A(\V1/V1/V2/A2/M4/s1 ),
    .B(\V1/V1/V2/A2/c3 ),
    .Z(\V1/V1/V2/s2 [3]));
 OR2_X1 \V1/V1/V2/A2/M4/_0_  (.A1(\V1/V1/V2/A2/M4/c1 ),
    .A2(\V1/V1/V2/A2/M4/c2 ),
    .ZN(\V1/V1/V2/c2 ));
 AND2_X1 \V1/V1/V2/A3/M1/M1/_0_  (.A1(\V1/V1/V2/v4 [0]),
    .A2(\V1/V1/V2/s2 [2]),
    .ZN(\V1/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M1/M1/_1_  (.A(\V1/V1/V2/v4 [0]),
    .B(\V1/V1/V2/s2 [2]),
    .Z(\V1/V1/V2/A3/M1/s1 ));
 AND2_X1 \V1/V1/V2/A3/M1/M2/_0_  (.A1(\V1/V1/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M1/M2/_1_  (.A(\V1/V1/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v2 [4]));
 OR2_X1 \V1/V1/V2/A3/M1/_0_  (.A1(\V1/V1/V2/A3/M1/c1 ),
    .A2(\V1/V1/V2/A3/M1/c2 ),
    .ZN(\V1/V1/V2/A3/c1 ));
 AND2_X1 \V1/V1/V2/A3/M2/M1/_0_  (.A1(\V1/V1/V2/v4 [1]),
    .A2(\V1/V1/V2/s2 [3]),
    .ZN(\V1/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M2/M1/_1_  (.A(\V1/V1/V2/v4 [1]),
    .B(\V1/V1/V2/s2 [3]),
    .Z(\V1/V1/V2/A3/M2/s1 ));
 AND2_X1 \V1/V1/V2/A3/M2/M2/_0_  (.A1(\V1/V1/V2/A3/M2/s1 ),
    .A2(\V1/V1/V2/A3/c1 ),
    .ZN(\V1/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M2/M2/_1_  (.A(\V1/V1/V2/A3/M2/s1 ),
    .B(\V1/V1/V2/A3/c1 ),
    .Z(\V1/V1/v2 [5]));
 OR2_X1 \V1/V1/V2/A3/M2/_0_  (.A1(\V1/V1/V2/A3/M2/c1 ),
    .A2(\V1/V1/V2/A3/M2/c2 ),
    .ZN(\V1/V1/V2/A3/c2 ));
 AND2_X1 \V1/V1/V2/A3/M3/M1/_0_  (.A1(\V1/V1/V2/v4 [2]),
    .A2(\V1/V1/V2/c3 ),
    .ZN(\V1/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M3/M1/_1_  (.A(\V1/V1/V2/v4 [2]),
    .B(\V1/V1/V2/c3 ),
    .Z(\V1/V1/V2/A3/M3/s1 ));
 AND2_X1 \V1/V1/V2/A3/M3/M2/_0_  (.A1(\V1/V1/V2/A3/M3/s1 ),
    .A2(\V1/V1/V2/A3/c2 ),
    .ZN(\V1/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M3/M2/_1_  (.A(\V1/V1/V2/A3/M3/s1 ),
    .B(\V1/V1/V2/A3/c2 ),
    .Z(\V1/V1/v2 [6]));
 OR2_X1 \V1/V1/V2/A3/M3/_0_  (.A1(\V1/V1/V2/A3/M3/c1 ),
    .A2(\V1/V1/V2/A3/M3/c2 ),
    .ZN(\V1/V1/V2/A3/c3 ));
 AND2_X1 \V1/V1/V2/A3/M4/M1/_0_  (.A1(\V1/V1/V2/v4 [3]),
    .A2(ground),
    .ZN(\V1/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M4/M1/_1_  (.A(\V1/V1/V2/v4 [3]),
    .B(ground),
    .Z(\V1/V1/V2/A3/M4/s1 ));
 AND2_X1 \V1/V1/V2/A3/M4/M2/_0_  (.A1(\V1/V1/V2/A3/M4/s1 ),
    .A2(\V1/V1/V2/A3/c3 ),
    .ZN(\V1/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M4/M2/_1_  (.A(\V1/V1/V2/A3/M4/s1 ),
    .B(\V1/V1/V2/A3/c3 ),
    .Z(\V1/V1/v2 [7]));
 OR2_X1 \V1/V1/V2/A3/M4/_0_  (.A1(\V1/V1/V2/A3/M4/c1 ),
    .A2(\V1/V1/V2/A3/M4/c2 ),
    .ZN(\V1/V1/V2/overflow ));
 AND2_X1 \V1/V1/V2/V1/HA1/_0_  (.A1(\V1/V1/V2/V1/w2 ),
    .A2(\V1/V1/V2/V1/w1 ),
    .ZN(\V1/V1/V2/V1/w4 ));
 XOR2_X2 \V1/V1/V2/V1/HA1/_1_  (.A(\V1/V1/V2/V1/w2 ),
    .B(\V1/V1/V2/V1/w1 ),
    .Z(\V1/V1/v2 [1]));
 AND2_X1 \V1/V1/V2/V1/HA2/_0_  (.A1(\V1/V1/V2/V1/w4 ),
    .A2(\V1/V1/V2/V1/w3 ),
    .ZN(\V1/V1/V2/v1 [3]));
 XOR2_X2 \V1/V1/V2/V1/HA2/_1_  (.A(\V1/V1/V2/V1/w4 ),
    .B(\V1/V1/V2/V1/w3 ),
    .Z(\V1/V1/V2/v1 [2]));
 AND2_X1 \V1/V1/V2/V1/_0_  (.A1(A[4]),
    .A2(B[0]),
    .ZN(\V1/V1/v2 [0]));
 AND2_X1 \V1/V1/V2/V1/_1_  (.A1(A[4]),
    .A2(B[1]),
    .ZN(\V1/V1/V2/V1/w1 ));
 AND2_X1 \V1/V1/V2/V1/_2_  (.A1(B[0]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V1/w2 ));
 AND2_X1 \V1/V1/V2/V1/_3_  (.A1(B[1]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V1/w3 ));
 AND2_X1 \V1/V1/V2/V2/HA1/_0_  (.A1(\V1/V1/V2/V2/w2 ),
    .A2(\V1/V1/V2/V2/w1 ),
    .ZN(\V1/V1/V2/V2/w4 ));
 XOR2_X2 \V1/V1/V2/V2/HA1/_1_  (.A(\V1/V1/V2/V2/w2 ),
    .B(\V1/V1/V2/V2/w1 ),
    .Z(\V1/V1/V2/v2 [1]));
 AND2_X1 \V1/V1/V2/V2/HA2/_0_  (.A1(\V1/V1/V2/V2/w4 ),
    .A2(\V1/V1/V2/V2/w3 ),
    .ZN(\V1/V1/V2/v2 [3]));
 XOR2_X2 \V1/V1/V2/V2/HA2/_1_  (.A(\V1/V1/V2/V2/w4 ),
    .B(\V1/V1/V2/V2/w3 ),
    .Z(\V1/V1/V2/v2 [2]));
 AND2_X1 \V1/V1/V2/V2/_0_  (.A1(A[6]),
    .A2(B[0]),
    .ZN(\V1/V1/V2/v2 [0]));
 AND2_X1 \V1/V1/V2/V2/_1_  (.A1(A[6]),
    .A2(B[1]),
    .ZN(\V1/V1/V2/V2/w1 ));
 AND2_X1 \V1/V1/V2/V2/_2_  (.A1(B[0]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V2/w2 ));
 AND2_X1 \V1/V1/V2/V2/_3_  (.A1(B[1]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V2/w3 ));
 AND2_X1 \V1/V1/V2/V3/HA1/_0_  (.A1(\V1/V1/V2/V3/w2 ),
    .A2(\V1/V1/V2/V3/w1 ),
    .ZN(\V1/V1/V2/V3/w4 ));
 XOR2_X2 \V1/V1/V2/V3/HA1/_1_  (.A(\V1/V1/V2/V3/w2 ),
    .B(\V1/V1/V2/V3/w1 ),
    .Z(\V1/V1/V2/v3 [1]));
 AND2_X1 \V1/V1/V2/V3/HA2/_0_  (.A1(\V1/V1/V2/V3/w4 ),
    .A2(\V1/V1/V2/V3/w3 ),
    .ZN(\V1/V1/V2/v3 [3]));
 XOR2_X2 \V1/V1/V2/V3/HA2/_1_  (.A(\V1/V1/V2/V3/w4 ),
    .B(\V1/V1/V2/V3/w3 ),
    .Z(\V1/V1/V2/v3 [2]));
 AND2_X1 \V1/V1/V2/V3/_0_  (.A1(A[4]),
    .A2(B[2]),
    .ZN(\V1/V1/V2/v3 [0]));
 AND2_X1 \V1/V1/V2/V3/_1_  (.A1(A[4]),
    .A2(B[3]),
    .ZN(\V1/V1/V2/V3/w1 ));
 AND2_X1 \V1/V1/V2/V3/_2_  (.A1(B[2]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V3/w2 ));
 AND2_X1 \V1/V1/V2/V3/_3_  (.A1(B[3]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V3/w3 ));
 AND2_X1 \V1/V1/V2/V4/HA1/_0_  (.A1(\V1/V1/V2/V4/w2 ),
    .A2(\V1/V1/V2/V4/w1 ),
    .ZN(\V1/V1/V2/V4/w4 ));
 XOR2_X2 \V1/V1/V2/V4/HA1/_1_  (.A(\V1/V1/V2/V4/w2 ),
    .B(\V1/V1/V2/V4/w1 ),
    .Z(\V1/V1/V2/v4 [1]));
 AND2_X1 \V1/V1/V2/V4/HA2/_0_  (.A1(\V1/V1/V2/V4/w4 ),
    .A2(\V1/V1/V2/V4/w3 ),
    .ZN(\V1/V1/V2/v4 [3]));
 XOR2_X2 \V1/V1/V2/V4/HA2/_1_  (.A(\V1/V1/V2/V4/w4 ),
    .B(\V1/V1/V2/V4/w3 ),
    .Z(\V1/V1/V2/v4 [2]));
 AND2_X1 \V1/V1/V2/V4/_0_  (.A1(A[6]),
    .A2(B[2]),
    .ZN(\V1/V1/V2/v4 [0]));
 AND2_X1 \V1/V1/V2/V4/_1_  (.A1(A[6]),
    .A2(B[3]),
    .ZN(\V1/V1/V2/V4/w1 ));
 AND2_X1 \V1/V1/V2/V4/_2_  (.A1(B[2]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V4/w2 ));
 AND2_X1 \V1/V1/V2/V4/_3_  (.A1(B[3]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V4/w3 ));
 OR2_X1 \V1/V1/V2/_0_  (.A1(\V1/V1/V2/c1 ),
    .A2(\V1/V1/V2/c2 ),
    .ZN(\V1/V1/V2/c3 ));
 AND2_X1 \V1/V1/V3/A1/M1/M1/_0_  (.A1(\V1/V1/V3/v2 [0]),
    .A2(\V1/V1/V3/v3 [0]),
    .ZN(\V1/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M1/M1/_1_  (.A(\V1/V1/V3/v2 [0]),
    .B(\V1/V1/V3/v3 [0]),
    .Z(\V1/V1/V3/A1/M1/s1 ));
 AND2_X1 \V1/V1/V3/A1/M1/M2/_0_  (.A1(\V1/V1/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M1/M2/_1_  (.A(\V1/V1/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/V3/s1 [0]));
 OR2_X1 \V1/V1/V3/A1/M1/_0_  (.A1(\V1/V1/V3/A1/M1/c1 ),
    .A2(\V1/V1/V3/A1/M1/c2 ),
    .ZN(\V1/V1/V3/A1/c1 ));
 AND2_X1 \V1/V1/V3/A1/M2/M1/_0_  (.A1(\V1/V1/V3/v2 [1]),
    .A2(\V1/V1/V3/v3 [1]),
    .ZN(\V1/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M2/M1/_1_  (.A(\V1/V1/V3/v2 [1]),
    .B(\V1/V1/V3/v3 [1]),
    .Z(\V1/V1/V3/A1/M2/s1 ));
 AND2_X1 \V1/V1/V3/A1/M2/M2/_0_  (.A1(\V1/V1/V3/A1/M2/s1 ),
    .A2(\V1/V1/V3/A1/c1 ),
    .ZN(\V1/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M2/M2/_1_  (.A(\V1/V1/V3/A1/M2/s1 ),
    .B(\V1/V1/V3/A1/c1 ),
    .Z(\V1/V1/V3/s1 [1]));
 OR2_X1 \V1/V1/V3/A1/M2/_0_  (.A1(\V1/V1/V3/A1/M2/c1 ),
    .A2(\V1/V1/V3/A1/M2/c2 ),
    .ZN(\V1/V1/V3/A1/c2 ));
 AND2_X1 \V1/V1/V3/A1/M3/M1/_0_  (.A1(\V1/V1/V3/v2 [2]),
    .A2(\V1/V1/V3/v3 [2]),
    .ZN(\V1/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M3/M1/_1_  (.A(\V1/V1/V3/v2 [2]),
    .B(\V1/V1/V3/v3 [2]),
    .Z(\V1/V1/V3/A1/M3/s1 ));
 AND2_X1 \V1/V1/V3/A1/M3/M2/_0_  (.A1(\V1/V1/V3/A1/M3/s1 ),
    .A2(\V1/V1/V3/A1/c2 ),
    .ZN(\V1/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M3/M2/_1_  (.A(\V1/V1/V3/A1/M3/s1 ),
    .B(\V1/V1/V3/A1/c2 ),
    .Z(\V1/V1/V3/s1 [2]));
 OR2_X1 \V1/V1/V3/A1/M3/_0_  (.A1(\V1/V1/V3/A1/M3/c1 ),
    .A2(\V1/V1/V3/A1/M3/c2 ),
    .ZN(\V1/V1/V3/A1/c3 ));
 AND2_X1 \V1/V1/V3/A1/M4/M1/_0_  (.A1(\V1/V1/V3/v2 [3]),
    .A2(\V1/V1/V3/v3 [3]),
    .ZN(\V1/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M4/M1/_1_  (.A(\V1/V1/V3/v2 [3]),
    .B(\V1/V1/V3/v3 [3]),
    .Z(\V1/V1/V3/A1/M4/s1 ));
 AND2_X1 \V1/V1/V3/A1/M4/M2/_0_  (.A1(\V1/V1/V3/A1/M4/s1 ),
    .A2(\V1/V1/V3/A1/c3 ),
    .ZN(\V1/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M4/M2/_1_  (.A(\V1/V1/V3/A1/M4/s1 ),
    .B(\V1/V1/V3/A1/c3 ),
    .Z(\V1/V1/V3/s1 [3]));
 OR2_X1 \V1/V1/V3/A1/M4/_0_  (.A1(\V1/V1/V3/A1/M4/c1 ),
    .A2(\V1/V1/V3/A1/M4/c2 ),
    .ZN(\V1/V1/V3/c1 ));
 AND2_X1 \V1/V1/V3/A2/M1/M1/_0_  (.A1(\V1/V1/V3/s1 [0]),
    .A2(\V1/V1/V3/v1 [2]),
    .ZN(\V1/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M1/M1/_1_  (.A(\V1/V1/V3/s1 [0]),
    .B(\V1/V1/V3/v1 [2]),
    .Z(\V1/V1/V3/A2/M1/s1 ));
 AND2_X1 \V1/V1/V3/A2/M1/M2/_0_  (.A1(\V1/V1/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M1/M2/_1_  (.A(\V1/V1/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v3 [2]));
 OR2_X1 \V1/V1/V3/A2/M1/_0_  (.A1(\V1/V1/V3/A2/M1/c1 ),
    .A2(\V1/V1/V3/A2/M1/c2 ),
    .ZN(\V1/V1/V3/A2/c1 ));
 AND2_X1 \V1/V1/V3/A2/M2/M1/_0_  (.A1(\V1/V1/V3/s1 [1]),
    .A2(\V1/V1/V3/v1 [3]),
    .ZN(\V1/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M2/M1/_1_  (.A(\V1/V1/V3/s1 [1]),
    .B(\V1/V1/V3/v1 [3]),
    .Z(\V1/V1/V3/A2/M2/s1 ));
 AND2_X1 \V1/V1/V3/A2/M2/M2/_0_  (.A1(\V1/V1/V3/A2/M2/s1 ),
    .A2(\V1/V1/V3/A2/c1 ),
    .ZN(\V1/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M2/M2/_1_  (.A(\V1/V1/V3/A2/M2/s1 ),
    .B(\V1/V1/V3/A2/c1 ),
    .Z(\V1/V1/v3 [3]));
 OR2_X1 \V1/V1/V3/A2/M2/_0_  (.A1(\V1/V1/V3/A2/M2/c1 ),
    .A2(\V1/V1/V3/A2/M2/c2 ),
    .ZN(\V1/V1/V3/A2/c2 ));
 AND2_X1 \V1/V1/V3/A2/M3/M1/_0_  (.A1(\V1/V1/V3/s1 [2]),
    .A2(ground),
    .ZN(\V1/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M3/M1/_1_  (.A(\V1/V1/V3/s1 [2]),
    .B(ground),
    .Z(\V1/V1/V3/A2/M3/s1 ));
 AND2_X1 \V1/V1/V3/A2/M3/M2/_0_  (.A1(\V1/V1/V3/A2/M3/s1 ),
    .A2(\V1/V1/V3/A2/c2 ),
    .ZN(\V1/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M3/M2/_1_  (.A(\V1/V1/V3/A2/M3/s1 ),
    .B(\V1/V1/V3/A2/c2 ),
    .Z(\V1/V1/V3/s2 [2]));
 OR2_X1 \V1/V1/V3/A2/M3/_0_  (.A1(\V1/V1/V3/A2/M3/c1 ),
    .A2(\V1/V1/V3/A2/M3/c2 ),
    .ZN(\V1/V1/V3/A2/c3 ));
 AND2_X1 \V1/V1/V3/A2/M4/M1/_0_  (.A1(\V1/V1/V3/s1 [3]),
    .A2(ground),
    .ZN(\V1/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M4/M1/_1_  (.A(\V1/V1/V3/s1 [3]),
    .B(ground),
    .Z(\V1/V1/V3/A2/M4/s1 ));
 AND2_X1 \V1/V1/V3/A2/M4/M2/_0_  (.A1(\V1/V1/V3/A2/M4/s1 ),
    .A2(\V1/V1/V3/A2/c3 ),
    .ZN(\V1/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M4/M2/_1_  (.A(\V1/V1/V3/A2/M4/s1 ),
    .B(\V1/V1/V3/A2/c3 ),
    .Z(\V1/V1/V3/s2 [3]));
 OR2_X1 \V1/V1/V3/A2/M4/_0_  (.A1(\V1/V1/V3/A2/M4/c1 ),
    .A2(\V1/V1/V3/A2/M4/c2 ),
    .ZN(\V1/V1/V3/c2 ));
 AND2_X1 \V1/V1/V3/A3/M1/M1/_0_  (.A1(\V1/V1/V3/v4 [0]),
    .A2(\V1/V1/V3/s2 [2]),
    .ZN(\V1/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M1/M1/_1_  (.A(\V1/V1/V3/v4 [0]),
    .B(\V1/V1/V3/s2 [2]),
    .Z(\V1/V1/V3/A3/M1/s1 ));
 AND2_X1 \V1/V1/V3/A3/M1/M2/_0_  (.A1(\V1/V1/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M1/M2/_1_  (.A(\V1/V1/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v3 [4]));
 OR2_X1 \V1/V1/V3/A3/M1/_0_  (.A1(\V1/V1/V3/A3/M1/c1 ),
    .A2(\V1/V1/V3/A3/M1/c2 ),
    .ZN(\V1/V1/V3/A3/c1 ));
 AND2_X1 \V1/V1/V3/A3/M2/M1/_0_  (.A1(\V1/V1/V3/v4 [1]),
    .A2(\V1/V1/V3/s2 [3]),
    .ZN(\V1/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M2/M1/_1_  (.A(\V1/V1/V3/v4 [1]),
    .B(\V1/V1/V3/s2 [3]),
    .Z(\V1/V1/V3/A3/M2/s1 ));
 AND2_X1 \V1/V1/V3/A3/M2/M2/_0_  (.A1(\V1/V1/V3/A3/M2/s1 ),
    .A2(\V1/V1/V3/A3/c1 ),
    .ZN(\V1/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M2/M2/_1_  (.A(\V1/V1/V3/A3/M2/s1 ),
    .B(\V1/V1/V3/A3/c1 ),
    .Z(\V1/V1/v3 [5]));
 OR2_X1 \V1/V1/V3/A3/M2/_0_  (.A1(\V1/V1/V3/A3/M2/c1 ),
    .A2(\V1/V1/V3/A3/M2/c2 ),
    .ZN(\V1/V1/V3/A3/c2 ));
 AND2_X1 \V1/V1/V3/A3/M3/M1/_0_  (.A1(\V1/V1/V3/v4 [2]),
    .A2(\V1/V1/V3/c3 ),
    .ZN(\V1/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M3/M1/_1_  (.A(\V1/V1/V3/v4 [2]),
    .B(\V1/V1/V3/c3 ),
    .Z(\V1/V1/V3/A3/M3/s1 ));
 AND2_X1 \V1/V1/V3/A3/M3/M2/_0_  (.A1(\V1/V1/V3/A3/M3/s1 ),
    .A2(\V1/V1/V3/A3/c2 ),
    .ZN(\V1/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M3/M2/_1_  (.A(\V1/V1/V3/A3/M3/s1 ),
    .B(\V1/V1/V3/A3/c2 ),
    .Z(\V1/V1/v3 [6]));
 OR2_X1 \V1/V1/V3/A3/M3/_0_  (.A1(\V1/V1/V3/A3/M3/c1 ),
    .A2(\V1/V1/V3/A3/M3/c2 ),
    .ZN(\V1/V1/V3/A3/c3 ));
 AND2_X1 \V1/V1/V3/A3/M4/M1/_0_  (.A1(\V1/V1/V3/v4 [3]),
    .A2(ground),
    .ZN(\V1/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M4/M1/_1_  (.A(\V1/V1/V3/v4 [3]),
    .B(ground),
    .Z(\V1/V1/V3/A3/M4/s1 ));
 AND2_X1 \V1/V1/V3/A3/M4/M2/_0_  (.A1(\V1/V1/V3/A3/M4/s1 ),
    .A2(\V1/V1/V3/A3/c3 ),
    .ZN(\V1/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M4/M2/_1_  (.A(\V1/V1/V3/A3/M4/s1 ),
    .B(\V1/V1/V3/A3/c3 ),
    .Z(\V1/V1/v3 [7]));
 OR2_X1 \V1/V1/V3/A3/M4/_0_  (.A1(\V1/V1/V3/A3/M4/c1 ),
    .A2(\V1/V1/V3/A3/M4/c2 ),
    .ZN(\V1/V1/V3/overflow ));
 AND2_X1 \V1/V1/V3/V1/HA1/_0_  (.A1(\V1/V1/V3/V1/w2 ),
    .A2(\V1/V1/V3/V1/w1 ),
    .ZN(\V1/V1/V3/V1/w4 ));
 XOR2_X2 \V1/V1/V3/V1/HA1/_1_  (.A(\V1/V1/V3/V1/w2 ),
    .B(\V1/V1/V3/V1/w1 ),
    .Z(\V1/V1/v3 [1]));
 AND2_X1 \V1/V1/V3/V1/HA2/_0_  (.A1(\V1/V1/V3/V1/w4 ),
    .A2(\V1/V1/V3/V1/w3 ),
    .ZN(\V1/V1/V3/v1 [3]));
 XOR2_X2 \V1/V1/V3/V1/HA2/_1_  (.A(\V1/V1/V3/V1/w4 ),
    .B(\V1/V1/V3/V1/w3 ),
    .Z(\V1/V1/V3/v1 [2]));
 AND2_X1 \V1/V1/V3/V1/_0_  (.A1(A[0]),
    .A2(B[4]),
    .ZN(\V1/V1/v3 [0]));
 AND2_X1 \V1/V1/V3/V1/_1_  (.A1(A[0]),
    .A2(B[5]),
    .ZN(\V1/V1/V3/V1/w1 ));
 AND2_X1 \V1/V1/V3/V1/_2_  (.A1(B[4]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V1/w2 ));
 AND2_X1 \V1/V1/V3/V1/_3_  (.A1(B[5]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V1/w3 ));
 AND2_X1 \V1/V1/V3/V2/HA1/_0_  (.A1(\V1/V1/V3/V2/w2 ),
    .A2(\V1/V1/V3/V2/w1 ),
    .ZN(\V1/V1/V3/V2/w4 ));
 XOR2_X2 \V1/V1/V3/V2/HA1/_1_  (.A(\V1/V1/V3/V2/w2 ),
    .B(\V1/V1/V3/V2/w1 ),
    .Z(\V1/V1/V3/v2 [1]));
 AND2_X1 \V1/V1/V3/V2/HA2/_0_  (.A1(\V1/V1/V3/V2/w4 ),
    .A2(\V1/V1/V3/V2/w3 ),
    .ZN(\V1/V1/V3/v2 [3]));
 XOR2_X2 \V1/V1/V3/V2/HA2/_1_  (.A(\V1/V1/V3/V2/w4 ),
    .B(\V1/V1/V3/V2/w3 ),
    .Z(\V1/V1/V3/v2 [2]));
 AND2_X1 \V1/V1/V3/V2/_0_  (.A1(A[2]),
    .A2(B[4]),
    .ZN(\V1/V1/V3/v2 [0]));
 AND2_X1 \V1/V1/V3/V2/_1_  (.A1(A[2]),
    .A2(B[5]),
    .ZN(\V1/V1/V3/V2/w1 ));
 AND2_X1 \V1/V1/V3/V2/_2_  (.A1(B[4]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V2/w2 ));
 AND2_X1 \V1/V1/V3/V2/_3_  (.A1(B[5]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V2/w3 ));
 AND2_X1 \V1/V1/V3/V3/HA1/_0_  (.A1(\V1/V1/V3/V3/w2 ),
    .A2(\V1/V1/V3/V3/w1 ),
    .ZN(\V1/V1/V3/V3/w4 ));
 XOR2_X2 \V1/V1/V3/V3/HA1/_1_  (.A(\V1/V1/V3/V3/w2 ),
    .B(\V1/V1/V3/V3/w1 ),
    .Z(\V1/V1/V3/v3 [1]));
 AND2_X1 \V1/V1/V3/V3/HA2/_0_  (.A1(\V1/V1/V3/V3/w4 ),
    .A2(\V1/V1/V3/V3/w3 ),
    .ZN(\V1/V1/V3/v3 [3]));
 XOR2_X2 \V1/V1/V3/V3/HA2/_1_  (.A(\V1/V1/V3/V3/w4 ),
    .B(\V1/V1/V3/V3/w3 ),
    .Z(\V1/V1/V3/v3 [2]));
 AND2_X1 \V1/V1/V3/V3/_0_  (.A1(A[0]),
    .A2(B[6]),
    .ZN(\V1/V1/V3/v3 [0]));
 AND2_X1 \V1/V1/V3/V3/_1_  (.A1(A[0]),
    .A2(B[7]),
    .ZN(\V1/V1/V3/V3/w1 ));
 AND2_X1 \V1/V1/V3/V3/_2_  (.A1(B[6]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V3/w2 ));
 AND2_X1 \V1/V1/V3/V3/_3_  (.A1(B[7]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V3/w3 ));
 AND2_X1 \V1/V1/V3/V4/HA1/_0_  (.A1(\V1/V1/V3/V4/w2 ),
    .A2(\V1/V1/V3/V4/w1 ),
    .ZN(\V1/V1/V3/V4/w4 ));
 XOR2_X2 \V1/V1/V3/V4/HA1/_1_  (.A(\V1/V1/V3/V4/w2 ),
    .B(\V1/V1/V3/V4/w1 ),
    .Z(\V1/V1/V3/v4 [1]));
 AND2_X1 \V1/V1/V3/V4/HA2/_0_  (.A1(\V1/V1/V3/V4/w4 ),
    .A2(\V1/V1/V3/V4/w3 ),
    .ZN(\V1/V1/V3/v4 [3]));
 XOR2_X2 \V1/V1/V3/V4/HA2/_1_  (.A(\V1/V1/V3/V4/w4 ),
    .B(\V1/V1/V3/V4/w3 ),
    .Z(\V1/V1/V3/v4 [2]));
 AND2_X1 \V1/V1/V3/V4/_0_  (.A1(A[2]),
    .A2(B[6]),
    .ZN(\V1/V1/V3/v4 [0]));
 AND2_X1 \V1/V1/V3/V4/_1_  (.A1(A[2]),
    .A2(B[7]),
    .ZN(\V1/V1/V3/V4/w1 ));
 AND2_X1 \V1/V1/V3/V4/_2_  (.A1(B[6]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V4/w2 ));
 AND2_X1 \V1/V1/V3/V4/_3_  (.A1(B[7]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V4/w3 ));
 OR2_X1 \V1/V1/V3/_0_  (.A1(\V1/V1/V3/c1 ),
    .A2(\V1/V1/V3/c2 ),
    .ZN(\V1/V1/V3/c3 ));
 AND2_X1 \V1/V1/V4/A1/M1/M1/_0_  (.A1(\V1/V1/V4/v2 [0]),
    .A2(\V1/V1/V4/v3 [0]),
    .ZN(\V1/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M1/M1/_1_  (.A(\V1/V1/V4/v2 [0]),
    .B(\V1/V1/V4/v3 [0]),
    .Z(\V1/V1/V4/A1/M1/s1 ));
 AND2_X1 \V1/V1/V4/A1/M1/M2/_0_  (.A1(\V1/V1/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M1/M2/_1_  (.A(\V1/V1/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/V4/s1 [0]));
 OR2_X1 \V1/V1/V4/A1/M1/_0_  (.A1(\V1/V1/V4/A1/M1/c1 ),
    .A2(\V1/V1/V4/A1/M1/c2 ),
    .ZN(\V1/V1/V4/A1/c1 ));
 AND2_X1 \V1/V1/V4/A1/M2/M1/_0_  (.A1(\V1/V1/V4/v2 [1]),
    .A2(\V1/V1/V4/v3 [1]),
    .ZN(\V1/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M2/M1/_1_  (.A(\V1/V1/V4/v2 [1]),
    .B(\V1/V1/V4/v3 [1]),
    .Z(\V1/V1/V4/A1/M2/s1 ));
 AND2_X1 \V1/V1/V4/A1/M2/M2/_0_  (.A1(\V1/V1/V4/A1/M2/s1 ),
    .A2(\V1/V1/V4/A1/c1 ),
    .ZN(\V1/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M2/M2/_1_  (.A(\V1/V1/V4/A1/M2/s1 ),
    .B(\V1/V1/V4/A1/c1 ),
    .Z(\V1/V1/V4/s1 [1]));
 OR2_X1 \V1/V1/V4/A1/M2/_0_  (.A1(\V1/V1/V4/A1/M2/c1 ),
    .A2(\V1/V1/V4/A1/M2/c2 ),
    .ZN(\V1/V1/V4/A1/c2 ));
 AND2_X1 \V1/V1/V4/A1/M3/M1/_0_  (.A1(\V1/V1/V4/v2 [2]),
    .A2(\V1/V1/V4/v3 [2]),
    .ZN(\V1/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M3/M1/_1_  (.A(\V1/V1/V4/v2 [2]),
    .B(\V1/V1/V4/v3 [2]),
    .Z(\V1/V1/V4/A1/M3/s1 ));
 AND2_X1 \V1/V1/V4/A1/M3/M2/_0_  (.A1(\V1/V1/V4/A1/M3/s1 ),
    .A2(\V1/V1/V4/A1/c2 ),
    .ZN(\V1/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M3/M2/_1_  (.A(\V1/V1/V4/A1/M3/s1 ),
    .B(\V1/V1/V4/A1/c2 ),
    .Z(\V1/V1/V4/s1 [2]));
 OR2_X1 \V1/V1/V4/A1/M3/_0_  (.A1(\V1/V1/V4/A1/M3/c1 ),
    .A2(\V1/V1/V4/A1/M3/c2 ),
    .ZN(\V1/V1/V4/A1/c3 ));
 AND2_X1 \V1/V1/V4/A1/M4/M1/_0_  (.A1(\V1/V1/V4/v2 [3]),
    .A2(\V1/V1/V4/v3 [3]),
    .ZN(\V1/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M4/M1/_1_  (.A(\V1/V1/V4/v2 [3]),
    .B(\V1/V1/V4/v3 [3]),
    .Z(\V1/V1/V4/A1/M4/s1 ));
 AND2_X1 \V1/V1/V4/A1/M4/M2/_0_  (.A1(\V1/V1/V4/A1/M4/s1 ),
    .A2(\V1/V1/V4/A1/c3 ),
    .ZN(\V1/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M4/M2/_1_  (.A(\V1/V1/V4/A1/M4/s1 ),
    .B(\V1/V1/V4/A1/c3 ),
    .Z(\V1/V1/V4/s1 [3]));
 OR2_X1 \V1/V1/V4/A1/M4/_0_  (.A1(\V1/V1/V4/A1/M4/c1 ),
    .A2(\V1/V1/V4/A1/M4/c2 ),
    .ZN(\V1/V1/V4/c1 ));
 AND2_X1 \V1/V1/V4/A2/M1/M1/_0_  (.A1(\V1/V1/V4/s1 [0]),
    .A2(\V1/V1/V4/v1 [2]),
    .ZN(\V1/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M1/M1/_1_  (.A(\V1/V1/V4/s1 [0]),
    .B(\V1/V1/V4/v1 [2]),
    .Z(\V1/V1/V4/A2/M1/s1 ));
 AND2_X1 \V1/V1/V4/A2/M1/M2/_0_  (.A1(\V1/V1/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M1/M2/_1_  (.A(\V1/V1/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v4 [2]));
 OR2_X1 \V1/V1/V4/A2/M1/_0_  (.A1(\V1/V1/V4/A2/M1/c1 ),
    .A2(\V1/V1/V4/A2/M1/c2 ),
    .ZN(\V1/V1/V4/A2/c1 ));
 AND2_X1 \V1/V1/V4/A2/M2/M1/_0_  (.A1(\V1/V1/V4/s1 [1]),
    .A2(\V1/V1/V4/v1 [3]),
    .ZN(\V1/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M2/M1/_1_  (.A(\V1/V1/V4/s1 [1]),
    .B(\V1/V1/V4/v1 [3]),
    .Z(\V1/V1/V4/A2/M2/s1 ));
 AND2_X1 \V1/V1/V4/A2/M2/M2/_0_  (.A1(\V1/V1/V4/A2/M2/s1 ),
    .A2(\V1/V1/V4/A2/c1 ),
    .ZN(\V1/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M2/M2/_1_  (.A(\V1/V1/V4/A2/M2/s1 ),
    .B(\V1/V1/V4/A2/c1 ),
    .Z(\V1/V1/v4 [3]));
 OR2_X1 \V1/V1/V4/A2/M2/_0_  (.A1(\V1/V1/V4/A2/M2/c1 ),
    .A2(\V1/V1/V4/A2/M2/c2 ),
    .ZN(\V1/V1/V4/A2/c2 ));
 AND2_X1 \V1/V1/V4/A2/M3/M1/_0_  (.A1(\V1/V1/V4/s1 [2]),
    .A2(ground),
    .ZN(\V1/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M3/M1/_1_  (.A(\V1/V1/V4/s1 [2]),
    .B(ground),
    .Z(\V1/V1/V4/A2/M3/s1 ));
 AND2_X1 \V1/V1/V4/A2/M3/M2/_0_  (.A1(\V1/V1/V4/A2/M3/s1 ),
    .A2(\V1/V1/V4/A2/c2 ),
    .ZN(\V1/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M3/M2/_1_  (.A(\V1/V1/V4/A2/M3/s1 ),
    .B(\V1/V1/V4/A2/c2 ),
    .Z(\V1/V1/V4/s2 [2]));
 OR2_X1 \V1/V1/V4/A2/M3/_0_  (.A1(\V1/V1/V4/A2/M3/c1 ),
    .A2(\V1/V1/V4/A2/M3/c2 ),
    .ZN(\V1/V1/V4/A2/c3 ));
 AND2_X1 \V1/V1/V4/A2/M4/M1/_0_  (.A1(\V1/V1/V4/s1 [3]),
    .A2(ground),
    .ZN(\V1/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M4/M1/_1_  (.A(\V1/V1/V4/s1 [3]),
    .B(ground),
    .Z(\V1/V1/V4/A2/M4/s1 ));
 AND2_X1 \V1/V1/V4/A2/M4/M2/_0_  (.A1(\V1/V1/V4/A2/M4/s1 ),
    .A2(\V1/V1/V4/A2/c3 ),
    .ZN(\V1/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M4/M2/_1_  (.A(\V1/V1/V4/A2/M4/s1 ),
    .B(\V1/V1/V4/A2/c3 ),
    .Z(\V1/V1/V4/s2 [3]));
 OR2_X1 \V1/V1/V4/A2/M4/_0_  (.A1(\V1/V1/V4/A2/M4/c1 ),
    .A2(\V1/V1/V4/A2/M4/c2 ),
    .ZN(\V1/V1/V4/c2 ));
 AND2_X1 \V1/V1/V4/A3/M1/M1/_0_  (.A1(\V1/V1/V4/v4 [0]),
    .A2(\V1/V1/V4/s2 [2]),
    .ZN(\V1/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M1/M1/_1_  (.A(\V1/V1/V4/v4 [0]),
    .B(\V1/V1/V4/s2 [2]),
    .Z(\V1/V1/V4/A3/M1/s1 ));
 AND2_X1 \V1/V1/V4/A3/M1/M2/_0_  (.A1(\V1/V1/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M1/M2/_1_  (.A(\V1/V1/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V1/v4 [4]));
 OR2_X1 \V1/V1/V4/A3/M1/_0_  (.A1(\V1/V1/V4/A3/M1/c1 ),
    .A2(\V1/V1/V4/A3/M1/c2 ),
    .ZN(\V1/V1/V4/A3/c1 ));
 AND2_X1 \V1/V1/V4/A3/M2/M1/_0_  (.A1(\V1/V1/V4/v4 [1]),
    .A2(\V1/V1/V4/s2 [3]),
    .ZN(\V1/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M2/M1/_1_  (.A(\V1/V1/V4/v4 [1]),
    .B(\V1/V1/V4/s2 [3]),
    .Z(\V1/V1/V4/A3/M2/s1 ));
 AND2_X1 \V1/V1/V4/A3/M2/M2/_0_  (.A1(\V1/V1/V4/A3/M2/s1 ),
    .A2(\V1/V1/V4/A3/c1 ),
    .ZN(\V1/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M2/M2/_1_  (.A(\V1/V1/V4/A3/M2/s1 ),
    .B(\V1/V1/V4/A3/c1 ),
    .Z(\V1/V1/v4 [5]));
 OR2_X1 \V1/V1/V4/A3/M2/_0_  (.A1(\V1/V1/V4/A3/M2/c1 ),
    .A2(\V1/V1/V4/A3/M2/c2 ),
    .ZN(\V1/V1/V4/A3/c2 ));
 AND2_X1 \V1/V1/V4/A3/M3/M1/_0_  (.A1(\V1/V1/V4/v4 [2]),
    .A2(\V1/V1/V4/c3 ),
    .ZN(\V1/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M3/M1/_1_  (.A(\V1/V1/V4/v4 [2]),
    .B(\V1/V1/V4/c3 ),
    .Z(\V1/V1/V4/A3/M3/s1 ));
 AND2_X1 \V1/V1/V4/A3/M3/M2/_0_  (.A1(\V1/V1/V4/A3/M3/s1 ),
    .A2(\V1/V1/V4/A3/c2 ),
    .ZN(\V1/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M3/M2/_1_  (.A(\V1/V1/V4/A3/M3/s1 ),
    .B(\V1/V1/V4/A3/c2 ),
    .Z(\V1/V1/v4 [6]));
 OR2_X1 \V1/V1/V4/A3/M3/_0_  (.A1(\V1/V1/V4/A3/M3/c1 ),
    .A2(\V1/V1/V4/A3/M3/c2 ),
    .ZN(\V1/V1/V4/A3/c3 ));
 AND2_X1 \V1/V1/V4/A3/M4/M1/_0_  (.A1(\V1/V1/V4/v4 [3]),
    .A2(ground),
    .ZN(\V1/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M4/M1/_1_  (.A(\V1/V1/V4/v4 [3]),
    .B(ground),
    .Z(\V1/V1/V4/A3/M4/s1 ));
 AND2_X1 \V1/V1/V4/A3/M4/M2/_0_  (.A1(\V1/V1/V4/A3/M4/s1 ),
    .A2(\V1/V1/V4/A3/c3 ),
    .ZN(\V1/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M4/M2/_1_  (.A(\V1/V1/V4/A3/M4/s1 ),
    .B(\V1/V1/V4/A3/c3 ),
    .Z(\V1/V1/v4 [7]));
 OR2_X1 \V1/V1/V4/A3/M4/_0_  (.A1(\V1/V1/V4/A3/M4/c1 ),
    .A2(\V1/V1/V4/A3/M4/c2 ),
    .ZN(\V1/V1/V4/overflow ));
 AND2_X1 \V1/V1/V4/V1/HA1/_0_  (.A1(\V1/V1/V4/V1/w2 ),
    .A2(\V1/V1/V4/V1/w1 ),
    .ZN(\V1/V1/V4/V1/w4 ));
 XOR2_X2 \V1/V1/V4/V1/HA1/_1_  (.A(\V1/V1/V4/V1/w2 ),
    .B(\V1/V1/V4/V1/w1 ),
    .Z(\V1/V1/v4 [1]));
 AND2_X1 \V1/V1/V4/V1/HA2/_0_  (.A1(\V1/V1/V4/V1/w4 ),
    .A2(\V1/V1/V4/V1/w3 ),
    .ZN(\V1/V1/V4/v1 [3]));
 XOR2_X2 \V1/V1/V4/V1/HA2/_1_  (.A(\V1/V1/V4/V1/w4 ),
    .B(\V1/V1/V4/V1/w3 ),
    .Z(\V1/V1/V4/v1 [2]));
 AND2_X1 \V1/V1/V4/V1/_0_  (.A1(A[4]),
    .A2(B[4]),
    .ZN(\V1/V1/v4 [0]));
 AND2_X1 \V1/V1/V4/V1/_1_  (.A1(A[4]),
    .A2(B[5]),
    .ZN(\V1/V1/V4/V1/w1 ));
 AND2_X1 \V1/V1/V4/V1/_2_  (.A1(B[4]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V1/w2 ));
 AND2_X1 \V1/V1/V4/V1/_3_  (.A1(B[5]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V1/w3 ));
 AND2_X1 \V1/V1/V4/V2/HA1/_0_  (.A1(\V1/V1/V4/V2/w2 ),
    .A2(\V1/V1/V4/V2/w1 ),
    .ZN(\V1/V1/V4/V2/w4 ));
 XOR2_X2 \V1/V1/V4/V2/HA1/_1_  (.A(\V1/V1/V4/V2/w2 ),
    .B(\V1/V1/V4/V2/w1 ),
    .Z(\V1/V1/V4/v2 [1]));
 AND2_X1 \V1/V1/V4/V2/HA2/_0_  (.A1(\V1/V1/V4/V2/w4 ),
    .A2(\V1/V1/V4/V2/w3 ),
    .ZN(\V1/V1/V4/v2 [3]));
 XOR2_X2 \V1/V1/V4/V2/HA2/_1_  (.A(\V1/V1/V4/V2/w4 ),
    .B(\V1/V1/V4/V2/w3 ),
    .Z(\V1/V1/V4/v2 [2]));
 AND2_X1 \V1/V1/V4/V2/_0_  (.A1(A[6]),
    .A2(B[4]),
    .ZN(\V1/V1/V4/v2 [0]));
 AND2_X1 \V1/V1/V4/V2/_1_  (.A1(A[6]),
    .A2(B[5]),
    .ZN(\V1/V1/V4/V2/w1 ));
 AND2_X1 \V1/V1/V4/V2/_2_  (.A1(B[4]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V2/w2 ));
 AND2_X1 \V1/V1/V4/V2/_3_  (.A1(B[5]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V2/w3 ));
 AND2_X1 \V1/V1/V4/V3/HA1/_0_  (.A1(\V1/V1/V4/V3/w2 ),
    .A2(\V1/V1/V4/V3/w1 ),
    .ZN(\V1/V1/V4/V3/w4 ));
 XOR2_X2 \V1/V1/V4/V3/HA1/_1_  (.A(\V1/V1/V4/V3/w2 ),
    .B(\V1/V1/V4/V3/w1 ),
    .Z(\V1/V1/V4/v3 [1]));
 AND2_X1 \V1/V1/V4/V3/HA2/_0_  (.A1(\V1/V1/V4/V3/w4 ),
    .A2(\V1/V1/V4/V3/w3 ),
    .ZN(\V1/V1/V4/v3 [3]));
 XOR2_X2 \V1/V1/V4/V3/HA2/_1_  (.A(\V1/V1/V4/V3/w4 ),
    .B(\V1/V1/V4/V3/w3 ),
    .Z(\V1/V1/V4/v3 [2]));
 AND2_X1 \V1/V1/V4/V3/_0_  (.A1(A[4]),
    .A2(B[6]),
    .ZN(\V1/V1/V4/v3 [0]));
 AND2_X1 \V1/V1/V4/V3/_1_  (.A1(A[4]),
    .A2(B[7]),
    .ZN(\V1/V1/V4/V3/w1 ));
 AND2_X1 \V1/V1/V4/V3/_2_  (.A1(B[6]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V3/w2 ));
 AND2_X1 \V1/V1/V4/V3/_3_  (.A1(B[7]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V3/w3 ));
 AND2_X1 \V1/V1/V4/V4/HA1/_0_  (.A1(\V1/V1/V4/V4/w2 ),
    .A2(\V1/V1/V4/V4/w1 ),
    .ZN(\V1/V1/V4/V4/w4 ));
 XOR2_X2 \V1/V1/V4/V4/HA1/_1_  (.A(\V1/V1/V4/V4/w2 ),
    .B(\V1/V1/V4/V4/w1 ),
    .Z(\V1/V1/V4/v4 [1]));
 AND2_X1 \V1/V1/V4/V4/HA2/_0_  (.A1(\V1/V1/V4/V4/w4 ),
    .A2(\V1/V1/V4/V4/w3 ),
    .ZN(\V1/V1/V4/v4 [3]));
 XOR2_X2 \V1/V1/V4/V4/HA2/_1_  (.A(\V1/V1/V4/V4/w4 ),
    .B(\V1/V1/V4/V4/w3 ),
    .Z(\V1/V1/V4/v4 [2]));
 AND2_X1 \V1/V1/V4/V4/_0_  (.A1(A[6]),
    .A2(B[6]),
    .ZN(\V1/V1/V4/v4 [0]));
 AND2_X1 \V1/V1/V4/V4/_1_  (.A1(A[6]),
    .A2(B[7]),
    .ZN(\V1/V1/V4/V4/w1 ));
 AND2_X1 \V1/V1/V4/V4/_2_  (.A1(B[6]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V4/w2 ));
 AND2_X1 \V1/V1/V4/V4/_3_  (.A1(B[7]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V4/w3 ));
 OR2_X1 \V1/V1/V4/_0_  (.A1(\V1/V1/V4/c1 ),
    .A2(\V1/V1/V4/c2 ),
    .ZN(\V1/V1/V4/c3 ));
 OR2_X1 \V1/V1/_0_  (.A1(\V1/V1/c1 ),
    .A2(\V1/V1/c2 ),
    .ZN(\V1/V1/c3 ));
 AND2_X1 \V1/V2/A1/A1/M1/M1/_0_  (.A1(\V1/V2/v2 [0]),
    .A2(\V1/V2/v3 [0]),
    .ZN(\V1/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M1/M1/_1_  (.A(\V1/V2/v2 [0]),
    .B(\V1/V2/v3 [0]),
    .Z(\V1/V2/A1/A1/M1/s1 ));
 AND2_X1 \V1/V2/A1/A1/M1/M2/_0_  (.A1(\V1/V2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M1/M2/_1_  (.A(\V1/V2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/s1 [0]));
 OR2_X1 \V1/V2/A1/A1/M1/_0_  (.A1(\V1/V2/A1/A1/M1/c1 ),
    .A2(\V1/V2/A1/A1/M1/c2 ),
    .ZN(\V1/V2/A1/A1/c1 ));
 AND2_X1 \V1/V2/A1/A1/M2/M1/_0_  (.A1(\V1/V2/v2 [1]),
    .A2(\V1/V2/v3 [1]),
    .ZN(\V1/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M2/M1/_1_  (.A(\V1/V2/v2 [1]),
    .B(\V1/V2/v3 [1]),
    .Z(\V1/V2/A1/A1/M2/s1 ));
 AND2_X1 \V1/V2/A1/A1/M2/M2/_0_  (.A1(\V1/V2/A1/A1/M2/s1 ),
    .A2(\V1/V2/A1/A1/c1 ),
    .ZN(\V1/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M2/M2/_1_  (.A(\V1/V2/A1/A1/M2/s1 ),
    .B(\V1/V2/A1/A1/c1 ),
    .Z(\V1/V2/s1 [1]));
 OR2_X1 \V1/V2/A1/A1/M2/_0_  (.A1(\V1/V2/A1/A1/M2/c1 ),
    .A2(\V1/V2/A1/A1/M2/c2 ),
    .ZN(\V1/V2/A1/A1/c2 ));
 AND2_X1 \V1/V2/A1/A1/M3/M1/_0_  (.A1(\V1/V2/v2 [2]),
    .A2(\V1/V2/v3 [2]),
    .ZN(\V1/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M3/M1/_1_  (.A(\V1/V2/v2 [2]),
    .B(\V1/V2/v3 [2]),
    .Z(\V1/V2/A1/A1/M3/s1 ));
 AND2_X1 \V1/V2/A1/A1/M3/M2/_0_  (.A1(\V1/V2/A1/A1/M3/s1 ),
    .A2(\V1/V2/A1/A1/c2 ),
    .ZN(\V1/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M3/M2/_1_  (.A(\V1/V2/A1/A1/M3/s1 ),
    .B(\V1/V2/A1/A1/c2 ),
    .Z(\V1/V2/s1 [2]));
 OR2_X1 \V1/V2/A1/A1/M3/_0_  (.A1(\V1/V2/A1/A1/M3/c1 ),
    .A2(\V1/V2/A1/A1/M3/c2 ),
    .ZN(\V1/V2/A1/A1/c3 ));
 AND2_X1 \V1/V2/A1/A1/M4/M1/_0_  (.A1(\V1/V2/v2 [3]),
    .A2(\V1/V2/v3 [3]),
    .ZN(\V1/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M4/M1/_1_  (.A(\V1/V2/v2 [3]),
    .B(\V1/V2/v3 [3]),
    .Z(\V1/V2/A1/A1/M4/s1 ));
 AND2_X1 \V1/V2/A1/A1/M4/M2/_0_  (.A1(\V1/V2/A1/A1/M4/s1 ),
    .A2(\V1/V2/A1/A1/c3 ),
    .ZN(\V1/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M4/M2/_1_  (.A(\V1/V2/A1/A1/M4/s1 ),
    .B(\V1/V2/A1/A1/c3 ),
    .Z(\V1/V2/s1 [3]));
 OR2_X1 \V1/V2/A1/A1/M4/_0_  (.A1(\V1/V2/A1/A1/M4/c1 ),
    .A2(\V1/V2/A1/A1/M4/c2 ),
    .ZN(\V1/V2/A1/c1 ));
 AND2_X1 \V1/V2/A1/A2/M1/M1/_0_  (.A1(\V1/V2/v2 [4]),
    .A2(\V1/V2/v3 [4]),
    .ZN(\V1/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M1/M1/_1_  (.A(\V1/V2/v2 [4]),
    .B(\V1/V2/v3 [4]),
    .Z(\V1/V2/A1/A2/M1/s1 ));
 AND2_X1 \V1/V2/A1/A2/M1/M2/_0_  (.A1(\V1/V2/A1/A2/M1/s1 ),
    .A2(\V1/V2/A1/c1 ),
    .ZN(\V1/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M1/M2/_1_  (.A(\V1/V2/A1/A2/M1/s1 ),
    .B(\V1/V2/A1/c1 ),
    .Z(\V1/V2/s1 [4]));
 OR2_X1 \V1/V2/A1/A2/M1/_0_  (.A1(\V1/V2/A1/A2/M1/c1 ),
    .A2(\V1/V2/A1/A2/M1/c2 ),
    .ZN(\V1/V2/A1/A2/c1 ));
 AND2_X1 \V1/V2/A1/A2/M2/M1/_0_  (.A1(\V1/V2/v2 [5]),
    .A2(\V1/V2/v3 [5]),
    .ZN(\V1/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M2/M1/_1_  (.A(\V1/V2/v2 [5]),
    .B(\V1/V2/v3 [5]),
    .Z(\V1/V2/A1/A2/M2/s1 ));
 AND2_X1 \V1/V2/A1/A2/M2/M2/_0_  (.A1(\V1/V2/A1/A2/M2/s1 ),
    .A2(\V1/V2/A1/A2/c1 ),
    .ZN(\V1/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M2/M2/_1_  (.A(\V1/V2/A1/A2/M2/s1 ),
    .B(\V1/V2/A1/A2/c1 ),
    .Z(\V1/V2/s1 [5]));
 OR2_X1 \V1/V2/A1/A2/M2/_0_  (.A1(\V1/V2/A1/A2/M2/c1 ),
    .A2(\V1/V2/A1/A2/M2/c2 ),
    .ZN(\V1/V2/A1/A2/c2 ));
 AND2_X1 \V1/V2/A1/A2/M3/M1/_0_  (.A1(\V1/V2/v2 [6]),
    .A2(\V1/V2/v3 [6]),
    .ZN(\V1/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M3/M1/_1_  (.A(\V1/V2/v2 [6]),
    .B(\V1/V2/v3 [6]),
    .Z(\V1/V2/A1/A2/M3/s1 ));
 AND2_X1 \V1/V2/A1/A2/M3/M2/_0_  (.A1(\V1/V2/A1/A2/M3/s1 ),
    .A2(\V1/V2/A1/A2/c2 ),
    .ZN(\V1/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M3/M2/_1_  (.A(\V1/V2/A1/A2/M3/s1 ),
    .B(\V1/V2/A1/A2/c2 ),
    .Z(\V1/V2/s1 [6]));
 OR2_X1 \V1/V2/A1/A2/M3/_0_  (.A1(\V1/V2/A1/A2/M3/c1 ),
    .A2(\V1/V2/A1/A2/M3/c2 ),
    .ZN(\V1/V2/A1/A2/c3 ));
 AND2_X1 \V1/V2/A1/A2/M4/M1/_0_  (.A1(\V1/V2/v2 [7]),
    .A2(\V1/V2/v3 [7]),
    .ZN(\V1/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M4/M1/_1_  (.A(\V1/V2/v2 [7]),
    .B(\V1/V2/v3 [7]),
    .Z(\V1/V2/A1/A2/M4/s1 ));
 AND2_X1 \V1/V2/A1/A2/M4/M2/_0_  (.A1(\V1/V2/A1/A2/M4/s1 ),
    .A2(\V1/V2/A1/A2/c3 ),
    .ZN(\V1/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M4/M2/_1_  (.A(\V1/V2/A1/A2/M4/s1 ),
    .B(\V1/V2/A1/A2/c3 ),
    .Z(\V1/V2/s1 [7]));
 OR2_X1 \V1/V2/A1/A2/M4/_0_  (.A1(\V1/V2/A1/A2/M4/c1 ),
    .A2(\V1/V2/A1/A2/M4/c2 ),
    .ZN(\V1/V2/c1 ));
 AND2_X1 \V1/V2/A2/A1/M1/M1/_0_  (.A1(\V1/V2/s1 [0]),
    .A2(\V1/V2/v1 [4]),
    .ZN(\V1/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M1/M1/_1_  (.A(\V1/V2/s1 [0]),
    .B(\V1/V2/v1 [4]),
    .Z(\V1/V2/A2/A1/M1/s1 ));
 AND2_X1 \V1/V2/A2/A1/M1/M2/_0_  (.A1(\V1/V2/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M1/M2/_1_  (.A(\V1/V2/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v2 [4]));
 OR2_X1 \V1/V2/A2/A1/M1/_0_  (.A1(\V1/V2/A2/A1/M1/c1 ),
    .A2(\V1/V2/A2/A1/M1/c2 ),
    .ZN(\V1/V2/A2/A1/c1 ));
 AND2_X1 \V1/V2/A2/A1/M2/M1/_0_  (.A1(\V1/V2/s1 [1]),
    .A2(\V1/V2/v1 [5]),
    .ZN(\V1/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M2/M1/_1_  (.A(\V1/V2/s1 [1]),
    .B(\V1/V2/v1 [5]),
    .Z(\V1/V2/A2/A1/M2/s1 ));
 AND2_X1 \V1/V2/A2/A1/M2/M2/_0_  (.A1(\V1/V2/A2/A1/M2/s1 ),
    .A2(\V1/V2/A2/A1/c1 ),
    .ZN(\V1/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M2/M2/_1_  (.A(\V1/V2/A2/A1/M2/s1 ),
    .B(\V1/V2/A2/A1/c1 ),
    .Z(\V1/v2 [5]));
 OR2_X1 \V1/V2/A2/A1/M2/_0_  (.A1(\V1/V2/A2/A1/M2/c1 ),
    .A2(\V1/V2/A2/A1/M2/c2 ),
    .ZN(\V1/V2/A2/A1/c2 ));
 AND2_X1 \V1/V2/A2/A1/M3/M1/_0_  (.A1(\V1/V2/s1 [2]),
    .A2(\V1/V2/v1 [6]),
    .ZN(\V1/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M3/M1/_1_  (.A(\V1/V2/s1 [2]),
    .B(\V1/V2/v1 [6]),
    .Z(\V1/V2/A2/A1/M3/s1 ));
 AND2_X1 \V1/V2/A2/A1/M3/M2/_0_  (.A1(\V1/V2/A2/A1/M3/s1 ),
    .A2(\V1/V2/A2/A1/c2 ),
    .ZN(\V1/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M3/M2/_1_  (.A(\V1/V2/A2/A1/M3/s1 ),
    .B(\V1/V2/A2/A1/c2 ),
    .Z(\V1/v2 [6]));
 OR2_X1 \V1/V2/A2/A1/M3/_0_  (.A1(\V1/V2/A2/A1/M3/c1 ),
    .A2(\V1/V2/A2/A1/M3/c2 ),
    .ZN(\V1/V2/A2/A1/c3 ));
 AND2_X1 \V1/V2/A2/A1/M4/M1/_0_  (.A1(\V1/V2/s1 [3]),
    .A2(\V1/V2/v1 [7]),
    .ZN(\V1/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M4/M1/_1_  (.A(\V1/V2/s1 [3]),
    .B(\V1/V2/v1 [7]),
    .Z(\V1/V2/A2/A1/M4/s1 ));
 AND2_X1 \V1/V2/A2/A1/M4/M2/_0_  (.A1(\V1/V2/A2/A1/M4/s1 ),
    .A2(\V1/V2/A2/A1/c3 ),
    .ZN(\V1/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M4/M2/_1_  (.A(\V1/V2/A2/A1/M4/s1 ),
    .B(\V1/V2/A2/A1/c3 ),
    .Z(\V1/v2 [7]));
 OR2_X1 \V1/V2/A2/A1/M4/_0_  (.A1(\V1/V2/A2/A1/M4/c1 ),
    .A2(\V1/V2/A2/A1/M4/c2 ),
    .ZN(\V1/V2/A2/c1 ));
 AND2_X1 \V1/V2/A2/A2/M1/M1/_0_  (.A1(\V1/V2/s1 [4]),
    .A2(ground),
    .ZN(\V1/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M1/M1/_1_  (.A(\V1/V2/s1 [4]),
    .B(ground),
    .Z(\V1/V2/A2/A2/M1/s1 ));
 AND2_X1 \V1/V2/A2/A2/M1/M2/_0_  (.A1(\V1/V2/A2/A2/M1/s1 ),
    .A2(\V1/V2/A2/c1 ),
    .ZN(\V1/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M1/M2/_1_  (.A(\V1/V2/A2/A2/M1/s1 ),
    .B(\V1/V2/A2/c1 ),
    .Z(\V1/V2/s2 [4]));
 OR2_X1 \V1/V2/A2/A2/M1/_0_  (.A1(\V1/V2/A2/A2/M1/c1 ),
    .A2(\V1/V2/A2/A2/M1/c2 ),
    .ZN(\V1/V2/A2/A2/c1 ));
 AND2_X1 \V1/V2/A2/A2/M2/M1/_0_  (.A1(\V1/V2/s1 [5]),
    .A2(ground),
    .ZN(\V1/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M2/M1/_1_  (.A(\V1/V2/s1 [5]),
    .B(ground),
    .Z(\V1/V2/A2/A2/M2/s1 ));
 AND2_X1 \V1/V2/A2/A2/M2/M2/_0_  (.A1(\V1/V2/A2/A2/M2/s1 ),
    .A2(\V1/V2/A2/A2/c1 ),
    .ZN(\V1/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M2/M2/_1_  (.A(\V1/V2/A2/A2/M2/s1 ),
    .B(\V1/V2/A2/A2/c1 ),
    .Z(\V1/V2/s2 [5]));
 OR2_X1 \V1/V2/A2/A2/M2/_0_  (.A1(\V1/V2/A2/A2/M2/c1 ),
    .A2(\V1/V2/A2/A2/M2/c2 ),
    .ZN(\V1/V2/A2/A2/c2 ));
 AND2_X1 \V1/V2/A2/A2/M3/M1/_0_  (.A1(\V1/V2/s1 [6]),
    .A2(ground),
    .ZN(\V1/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M3/M1/_1_  (.A(\V1/V2/s1 [6]),
    .B(ground),
    .Z(\V1/V2/A2/A2/M3/s1 ));
 AND2_X1 \V1/V2/A2/A2/M3/M2/_0_  (.A1(\V1/V2/A2/A2/M3/s1 ),
    .A2(\V1/V2/A2/A2/c2 ),
    .ZN(\V1/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M3/M2/_1_  (.A(\V1/V2/A2/A2/M3/s1 ),
    .B(\V1/V2/A2/A2/c2 ),
    .Z(\V1/V2/s2 [6]));
 OR2_X1 \V1/V2/A2/A2/M3/_0_  (.A1(\V1/V2/A2/A2/M3/c1 ),
    .A2(\V1/V2/A2/A2/M3/c2 ),
    .ZN(\V1/V2/A2/A2/c3 ));
 AND2_X1 \V1/V2/A2/A2/M4/M1/_0_  (.A1(\V1/V2/s1 [7]),
    .A2(ground),
    .ZN(\V1/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M4/M1/_1_  (.A(\V1/V2/s1 [7]),
    .B(ground),
    .Z(\V1/V2/A2/A2/M4/s1 ));
 AND2_X1 \V1/V2/A2/A2/M4/M2/_0_  (.A1(\V1/V2/A2/A2/M4/s1 ),
    .A2(\V1/V2/A2/A2/c3 ),
    .ZN(\V1/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M4/M2/_1_  (.A(\V1/V2/A2/A2/M4/s1 ),
    .B(\V1/V2/A2/A2/c3 ),
    .Z(\V1/V2/s2 [7]));
 OR2_X1 \V1/V2/A2/A2/M4/_0_  (.A1(\V1/V2/A2/A2/M4/c1 ),
    .A2(\V1/V2/A2/A2/M4/c2 ),
    .ZN(\V1/V2/c2 ));
 AND2_X1 \V1/V2/A3/A1/M1/M1/_0_  (.A1(\V1/V2/v4 [0]),
    .A2(\V1/V2/s2 [4]),
    .ZN(\V1/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M1/M1/_1_  (.A(\V1/V2/v4 [0]),
    .B(\V1/V2/s2 [4]),
    .Z(\V1/V2/A3/A1/M1/s1 ));
 AND2_X1 \V1/V2/A3/A1/M1/M2/_0_  (.A1(\V1/V2/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M1/M2/_1_  (.A(\V1/V2/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v2 [8]));
 OR2_X1 \V1/V2/A3/A1/M1/_0_  (.A1(\V1/V2/A3/A1/M1/c1 ),
    .A2(\V1/V2/A3/A1/M1/c2 ),
    .ZN(\V1/V2/A3/A1/c1 ));
 AND2_X1 \V1/V2/A3/A1/M2/M1/_0_  (.A1(\V1/V2/v4 [1]),
    .A2(\V1/V2/s2 [5]),
    .ZN(\V1/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M2/M1/_1_  (.A(\V1/V2/v4 [1]),
    .B(\V1/V2/s2 [5]),
    .Z(\V1/V2/A3/A1/M2/s1 ));
 AND2_X1 \V1/V2/A3/A1/M2/M2/_0_  (.A1(\V1/V2/A3/A1/M2/s1 ),
    .A2(\V1/V2/A3/A1/c1 ),
    .ZN(\V1/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M2/M2/_1_  (.A(\V1/V2/A3/A1/M2/s1 ),
    .B(\V1/V2/A3/A1/c1 ),
    .Z(\V1/v2 [9]));
 OR2_X1 \V1/V2/A3/A1/M2/_0_  (.A1(\V1/V2/A3/A1/M2/c1 ),
    .A2(\V1/V2/A3/A1/M2/c2 ),
    .ZN(\V1/V2/A3/A1/c2 ));
 AND2_X1 \V1/V2/A3/A1/M3/M1/_0_  (.A1(\V1/V2/v4 [2]),
    .A2(\V1/V2/s2 [6]),
    .ZN(\V1/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M3/M1/_1_  (.A(\V1/V2/v4 [2]),
    .B(\V1/V2/s2 [6]),
    .Z(\V1/V2/A3/A1/M3/s1 ));
 AND2_X1 \V1/V2/A3/A1/M3/M2/_0_  (.A1(\V1/V2/A3/A1/M3/s1 ),
    .A2(\V1/V2/A3/A1/c2 ),
    .ZN(\V1/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M3/M2/_1_  (.A(\V1/V2/A3/A1/M3/s1 ),
    .B(\V1/V2/A3/A1/c2 ),
    .Z(\V1/v2 [10]));
 OR2_X1 \V1/V2/A3/A1/M3/_0_  (.A1(\V1/V2/A3/A1/M3/c1 ),
    .A2(\V1/V2/A3/A1/M3/c2 ),
    .ZN(\V1/V2/A3/A1/c3 ));
 AND2_X1 \V1/V2/A3/A1/M4/M1/_0_  (.A1(\V1/V2/v4 [3]),
    .A2(\V1/V2/s2 [7]),
    .ZN(\V1/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M4/M1/_1_  (.A(\V1/V2/v4 [3]),
    .B(\V1/V2/s2 [7]),
    .Z(\V1/V2/A3/A1/M4/s1 ));
 AND2_X1 \V1/V2/A3/A1/M4/M2/_0_  (.A1(\V1/V2/A3/A1/M4/s1 ),
    .A2(\V1/V2/A3/A1/c3 ),
    .ZN(\V1/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M4/M2/_1_  (.A(\V1/V2/A3/A1/M4/s1 ),
    .B(\V1/V2/A3/A1/c3 ),
    .Z(\V1/v2 [11]));
 OR2_X1 \V1/V2/A3/A1/M4/_0_  (.A1(\V1/V2/A3/A1/M4/c1 ),
    .A2(\V1/V2/A3/A1/M4/c2 ),
    .ZN(\V1/V2/A3/c1 ));
 AND2_X1 \V1/V2/A3/A2/M1/M1/_0_  (.A1(\V1/V2/v4 [4]),
    .A2(\V1/V2/c3 ),
    .ZN(\V1/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M1/M1/_1_  (.A(\V1/V2/v4 [4]),
    .B(\V1/V2/c3 ),
    .Z(\V1/V2/A3/A2/M1/s1 ));
 AND2_X1 \V1/V2/A3/A2/M1/M2/_0_  (.A1(\V1/V2/A3/A2/M1/s1 ),
    .A2(\V1/V2/A3/c1 ),
    .ZN(\V1/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M1/M2/_1_  (.A(\V1/V2/A3/A2/M1/s1 ),
    .B(\V1/V2/A3/c1 ),
    .Z(\V1/v2 [12]));
 OR2_X1 \V1/V2/A3/A2/M1/_0_  (.A1(\V1/V2/A3/A2/M1/c1 ),
    .A2(\V1/V2/A3/A2/M1/c2 ),
    .ZN(\V1/V2/A3/A2/c1 ));
 AND2_X1 \V1/V2/A3/A2/M2/M1/_0_  (.A1(\V1/V2/v4 [5]),
    .A2(ground),
    .ZN(\V1/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M2/M1/_1_  (.A(\V1/V2/v4 [5]),
    .B(ground),
    .Z(\V1/V2/A3/A2/M2/s1 ));
 AND2_X1 \V1/V2/A3/A2/M2/M2/_0_  (.A1(\V1/V2/A3/A2/M2/s1 ),
    .A2(\V1/V2/A3/A2/c1 ),
    .ZN(\V1/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M2/M2/_1_  (.A(\V1/V2/A3/A2/M2/s1 ),
    .B(\V1/V2/A3/A2/c1 ),
    .Z(\V1/v2 [13]));
 OR2_X1 \V1/V2/A3/A2/M2/_0_  (.A1(\V1/V2/A3/A2/M2/c1 ),
    .A2(\V1/V2/A3/A2/M2/c2 ),
    .ZN(\V1/V2/A3/A2/c2 ));
 AND2_X1 \V1/V2/A3/A2/M3/M1/_0_  (.A1(\V1/V2/v4 [6]),
    .A2(ground),
    .ZN(\V1/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M3/M1/_1_  (.A(\V1/V2/v4 [6]),
    .B(ground),
    .Z(\V1/V2/A3/A2/M3/s1 ));
 AND2_X1 \V1/V2/A3/A2/M3/M2/_0_  (.A1(\V1/V2/A3/A2/M3/s1 ),
    .A2(\V1/V2/A3/A2/c2 ),
    .ZN(\V1/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M3/M2/_1_  (.A(\V1/V2/A3/A2/M3/s1 ),
    .B(\V1/V2/A3/A2/c2 ),
    .Z(\V1/v2 [14]));
 OR2_X1 \V1/V2/A3/A2/M3/_0_  (.A1(\V1/V2/A3/A2/M3/c1 ),
    .A2(\V1/V2/A3/A2/M3/c2 ),
    .ZN(\V1/V2/A3/A2/c3 ));
 AND2_X1 \V1/V2/A3/A2/M4/M1/_0_  (.A1(\V1/V2/v4 [7]),
    .A2(ground),
    .ZN(\V1/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M4/M1/_1_  (.A(\V1/V2/v4 [7]),
    .B(ground),
    .Z(\V1/V2/A3/A2/M4/s1 ));
 AND2_X1 \V1/V2/A3/A2/M4/M2/_0_  (.A1(\V1/V2/A3/A2/M4/s1 ),
    .A2(\V1/V2/A3/A2/c3 ),
    .ZN(\V1/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M4/M2/_1_  (.A(\V1/V2/A3/A2/M4/s1 ),
    .B(\V1/V2/A3/A2/c3 ),
    .Z(\V1/v2 [15]));
 OR2_X1 \V1/V2/A3/A2/M4/_0_  (.A1(\V1/V2/A3/A2/M4/c1 ),
    .A2(\V1/V2/A3/A2/M4/c2 ),
    .ZN(\V1/V2/overflow ));
 AND2_X1 \V1/V2/V1/A1/M1/M1/_0_  (.A1(\V1/V2/V1/v2 [0]),
    .A2(\V1/V2/V1/v3 [0]),
    .ZN(\V1/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M1/M1/_1_  (.A(\V1/V2/V1/v2 [0]),
    .B(\V1/V2/V1/v3 [0]),
    .Z(\V1/V2/V1/A1/M1/s1 ));
 AND2_X1 \V1/V2/V1/A1/M1/M2/_0_  (.A1(\V1/V2/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M1/M2/_1_  (.A(\V1/V2/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/V1/s1 [0]));
 OR2_X1 \V1/V2/V1/A1/M1/_0_  (.A1(\V1/V2/V1/A1/M1/c1 ),
    .A2(\V1/V2/V1/A1/M1/c2 ),
    .ZN(\V1/V2/V1/A1/c1 ));
 AND2_X1 \V1/V2/V1/A1/M2/M1/_0_  (.A1(\V1/V2/V1/v2 [1]),
    .A2(\V1/V2/V1/v3 [1]),
    .ZN(\V1/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M2/M1/_1_  (.A(\V1/V2/V1/v2 [1]),
    .B(\V1/V2/V1/v3 [1]),
    .Z(\V1/V2/V1/A1/M2/s1 ));
 AND2_X1 \V1/V2/V1/A1/M2/M2/_0_  (.A1(\V1/V2/V1/A1/M2/s1 ),
    .A2(\V1/V2/V1/A1/c1 ),
    .ZN(\V1/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M2/M2/_1_  (.A(\V1/V2/V1/A1/M2/s1 ),
    .B(\V1/V2/V1/A1/c1 ),
    .Z(\V1/V2/V1/s1 [1]));
 OR2_X1 \V1/V2/V1/A1/M2/_0_  (.A1(\V1/V2/V1/A1/M2/c1 ),
    .A2(\V1/V2/V1/A1/M2/c2 ),
    .ZN(\V1/V2/V1/A1/c2 ));
 AND2_X1 \V1/V2/V1/A1/M3/M1/_0_  (.A1(\V1/V2/V1/v2 [2]),
    .A2(\V1/V2/V1/v3 [2]),
    .ZN(\V1/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M3/M1/_1_  (.A(\V1/V2/V1/v2 [2]),
    .B(\V1/V2/V1/v3 [2]),
    .Z(\V1/V2/V1/A1/M3/s1 ));
 AND2_X1 \V1/V2/V1/A1/M3/M2/_0_  (.A1(\V1/V2/V1/A1/M3/s1 ),
    .A2(\V1/V2/V1/A1/c2 ),
    .ZN(\V1/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M3/M2/_1_  (.A(\V1/V2/V1/A1/M3/s1 ),
    .B(\V1/V2/V1/A1/c2 ),
    .Z(\V1/V2/V1/s1 [2]));
 OR2_X1 \V1/V2/V1/A1/M3/_0_  (.A1(\V1/V2/V1/A1/M3/c1 ),
    .A2(\V1/V2/V1/A1/M3/c2 ),
    .ZN(\V1/V2/V1/A1/c3 ));
 AND2_X1 \V1/V2/V1/A1/M4/M1/_0_  (.A1(\V1/V2/V1/v2 [3]),
    .A2(\V1/V2/V1/v3 [3]),
    .ZN(\V1/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M4/M1/_1_  (.A(\V1/V2/V1/v2 [3]),
    .B(\V1/V2/V1/v3 [3]),
    .Z(\V1/V2/V1/A1/M4/s1 ));
 AND2_X1 \V1/V2/V1/A1/M4/M2/_0_  (.A1(\V1/V2/V1/A1/M4/s1 ),
    .A2(\V1/V2/V1/A1/c3 ),
    .ZN(\V1/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M4/M2/_1_  (.A(\V1/V2/V1/A1/M4/s1 ),
    .B(\V1/V2/V1/A1/c3 ),
    .Z(\V1/V2/V1/s1 [3]));
 OR2_X1 \V1/V2/V1/A1/M4/_0_  (.A1(\V1/V2/V1/A1/M4/c1 ),
    .A2(\V1/V2/V1/A1/M4/c2 ),
    .ZN(\V1/V2/V1/c1 ));
 AND2_X1 \V1/V2/V1/A2/M1/M1/_0_  (.A1(\V1/V2/V1/s1 [0]),
    .A2(\V1/V2/V1/v1 [2]),
    .ZN(\V1/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M1/M1/_1_  (.A(\V1/V2/V1/s1 [0]),
    .B(\V1/V2/V1/v1 [2]),
    .Z(\V1/V2/V1/A2/M1/s1 ));
 AND2_X1 \V1/V2/V1/A2/M1/M2/_0_  (.A1(\V1/V2/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M1/M2/_1_  (.A(\V1/V2/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/v2 [2]));
 OR2_X1 \V1/V2/V1/A2/M1/_0_  (.A1(\V1/V2/V1/A2/M1/c1 ),
    .A2(\V1/V2/V1/A2/M1/c2 ),
    .ZN(\V1/V2/V1/A2/c1 ));
 AND2_X1 \V1/V2/V1/A2/M2/M1/_0_  (.A1(\V1/V2/V1/s1 [1]),
    .A2(\V1/V2/V1/v1 [3]),
    .ZN(\V1/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M2/M1/_1_  (.A(\V1/V2/V1/s1 [1]),
    .B(\V1/V2/V1/v1 [3]),
    .Z(\V1/V2/V1/A2/M2/s1 ));
 AND2_X1 \V1/V2/V1/A2/M2/M2/_0_  (.A1(\V1/V2/V1/A2/M2/s1 ),
    .A2(\V1/V2/V1/A2/c1 ),
    .ZN(\V1/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M2/M2/_1_  (.A(\V1/V2/V1/A2/M2/s1 ),
    .B(\V1/V2/V1/A2/c1 ),
    .Z(\V1/v2 [3]));
 OR2_X1 \V1/V2/V1/A2/M2/_0_  (.A1(\V1/V2/V1/A2/M2/c1 ),
    .A2(\V1/V2/V1/A2/M2/c2 ),
    .ZN(\V1/V2/V1/A2/c2 ));
 AND2_X1 \V1/V2/V1/A2/M3/M1/_0_  (.A1(\V1/V2/V1/s1 [2]),
    .A2(ground),
    .ZN(\V1/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M3/M1/_1_  (.A(\V1/V2/V1/s1 [2]),
    .B(ground),
    .Z(\V1/V2/V1/A2/M3/s1 ));
 AND2_X1 \V1/V2/V1/A2/M3/M2/_0_  (.A1(\V1/V2/V1/A2/M3/s1 ),
    .A2(\V1/V2/V1/A2/c2 ),
    .ZN(\V1/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M3/M2/_1_  (.A(\V1/V2/V1/A2/M3/s1 ),
    .B(\V1/V2/V1/A2/c2 ),
    .Z(\V1/V2/V1/s2 [2]));
 OR2_X1 \V1/V2/V1/A2/M3/_0_  (.A1(\V1/V2/V1/A2/M3/c1 ),
    .A2(\V1/V2/V1/A2/M3/c2 ),
    .ZN(\V1/V2/V1/A2/c3 ));
 AND2_X1 \V1/V2/V1/A2/M4/M1/_0_  (.A1(\V1/V2/V1/s1 [3]),
    .A2(ground),
    .ZN(\V1/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M4/M1/_1_  (.A(\V1/V2/V1/s1 [3]),
    .B(ground),
    .Z(\V1/V2/V1/A2/M4/s1 ));
 AND2_X1 \V1/V2/V1/A2/M4/M2/_0_  (.A1(\V1/V2/V1/A2/M4/s1 ),
    .A2(\V1/V2/V1/A2/c3 ),
    .ZN(\V1/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M4/M2/_1_  (.A(\V1/V2/V1/A2/M4/s1 ),
    .B(\V1/V2/V1/A2/c3 ),
    .Z(\V1/V2/V1/s2 [3]));
 OR2_X1 \V1/V2/V1/A2/M4/_0_  (.A1(\V1/V2/V1/A2/M4/c1 ),
    .A2(\V1/V2/V1/A2/M4/c2 ),
    .ZN(\V1/V2/V1/c2 ));
 AND2_X1 \V1/V2/V1/A3/M1/M1/_0_  (.A1(\V1/V2/V1/v4 [0]),
    .A2(\V1/V2/V1/s2 [2]),
    .ZN(\V1/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M1/M1/_1_  (.A(\V1/V2/V1/v4 [0]),
    .B(\V1/V2/V1/s2 [2]),
    .Z(\V1/V2/V1/A3/M1/s1 ));
 AND2_X1 \V1/V2/V1/A3/M1/M2/_0_  (.A1(\V1/V2/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M1/M2/_1_  (.A(\V1/V2/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v1 [4]));
 OR2_X1 \V1/V2/V1/A3/M1/_0_  (.A1(\V1/V2/V1/A3/M1/c1 ),
    .A2(\V1/V2/V1/A3/M1/c2 ),
    .ZN(\V1/V2/V1/A3/c1 ));
 AND2_X1 \V1/V2/V1/A3/M2/M1/_0_  (.A1(\V1/V2/V1/v4 [1]),
    .A2(\V1/V2/V1/s2 [3]),
    .ZN(\V1/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M2/M1/_1_  (.A(\V1/V2/V1/v4 [1]),
    .B(\V1/V2/V1/s2 [3]),
    .Z(\V1/V2/V1/A3/M2/s1 ));
 AND2_X1 \V1/V2/V1/A3/M2/M2/_0_  (.A1(\V1/V2/V1/A3/M2/s1 ),
    .A2(\V1/V2/V1/A3/c1 ),
    .ZN(\V1/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M2/M2/_1_  (.A(\V1/V2/V1/A3/M2/s1 ),
    .B(\V1/V2/V1/A3/c1 ),
    .Z(\V1/V2/v1 [5]));
 OR2_X1 \V1/V2/V1/A3/M2/_0_  (.A1(\V1/V2/V1/A3/M2/c1 ),
    .A2(\V1/V2/V1/A3/M2/c2 ),
    .ZN(\V1/V2/V1/A3/c2 ));
 AND2_X1 \V1/V2/V1/A3/M3/M1/_0_  (.A1(\V1/V2/V1/v4 [2]),
    .A2(\V1/V2/V1/c3 ),
    .ZN(\V1/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M3/M1/_1_  (.A(\V1/V2/V1/v4 [2]),
    .B(\V1/V2/V1/c3 ),
    .Z(\V1/V2/V1/A3/M3/s1 ));
 AND2_X1 \V1/V2/V1/A3/M3/M2/_0_  (.A1(\V1/V2/V1/A3/M3/s1 ),
    .A2(\V1/V2/V1/A3/c2 ),
    .ZN(\V1/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M3/M2/_1_  (.A(\V1/V2/V1/A3/M3/s1 ),
    .B(\V1/V2/V1/A3/c2 ),
    .Z(\V1/V2/v1 [6]));
 OR2_X1 \V1/V2/V1/A3/M3/_0_  (.A1(\V1/V2/V1/A3/M3/c1 ),
    .A2(\V1/V2/V1/A3/M3/c2 ),
    .ZN(\V1/V2/V1/A3/c3 ));
 AND2_X1 \V1/V2/V1/A3/M4/M1/_0_  (.A1(\V1/V2/V1/v4 [3]),
    .A2(ground),
    .ZN(\V1/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M4/M1/_1_  (.A(\V1/V2/V1/v4 [3]),
    .B(ground),
    .Z(\V1/V2/V1/A3/M4/s1 ));
 AND2_X1 \V1/V2/V1/A3/M4/M2/_0_  (.A1(\V1/V2/V1/A3/M4/s1 ),
    .A2(\V1/V2/V1/A3/c3 ),
    .ZN(\V1/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M4/M2/_1_  (.A(\V1/V2/V1/A3/M4/s1 ),
    .B(\V1/V2/V1/A3/c3 ),
    .Z(\V1/V2/v1 [7]));
 OR2_X1 \V1/V2/V1/A3/M4/_0_  (.A1(\V1/V2/V1/A3/M4/c1 ),
    .A2(\V1/V2/V1/A3/M4/c2 ),
    .ZN(\V1/V2/V1/overflow ));
 AND2_X1 \V1/V2/V1/V1/HA1/_0_  (.A1(\V1/V2/V1/V1/w2 ),
    .A2(\V1/V2/V1/V1/w1 ),
    .ZN(\V1/V2/V1/V1/w4 ));
 XOR2_X2 \V1/V2/V1/V1/HA1/_1_  (.A(\V1/V2/V1/V1/w2 ),
    .B(\V1/V2/V1/V1/w1 ),
    .Z(\V1/v2 [1]));
 AND2_X1 \V1/V2/V1/V1/HA2/_0_  (.A1(\V1/V2/V1/V1/w4 ),
    .A2(\V1/V2/V1/V1/w3 ),
    .ZN(\V1/V2/V1/v1 [3]));
 XOR2_X2 \V1/V2/V1/V1/HA2/_1_  (.A(\V1/V2/V1/V1/w4 ),
    .B(\V1/V2/V1/V1/w3 ),
    .Z(\V1/V2/V1/v1 [2]));
 AND2_X1 \V1/V2/V1/V1/_0_  (.A1(A[8]),
    .A2(B[0]),
    .ZN(\V1/v2 [0]));
 AND2_X1 \V1/V2/V1/V1/_1_  (.A1(A[8]),
    .A2(B[1]),
    .ZN(\V1/V2/V1/V1/w1 ));
 AND2_X1 \V1/V2/V1/V1/_2_  (.A1(B[0]),
    .A2(A[9]),
    .ZN(\V1/V2/V1/V1/w2 ));
 AND2_X1 \V1/V2/V1/V1/_3_  (.A1(B[1]),
    .A2(A[9]),
    .ZN(\V1/V2/V1/V1/w3 ));
 AND2_X1 \V1/V2/V1/V2/HA1/_0_  (.A1(\V1/V2/V1/V2/w2 ),
    .A2(\V1/V2/V1/V2/w1 ),
    .ZN(\V1/V2/V1/V2/w4 ));
 XOR2_X2 \V1/V2/V1/V2/HA1/_1_  (.A(\V1/V2/V1/V2/w2 ),
    .B(\V1/V2/V1/V2/w1 ),
    .Z(\V1/V2/V1/v2 [1]));
 AND2_X1 \V1/V2/V1/V2/HA2/_0_  (.A1(\V1/V2/V1/V2/w4 ),
    .A2(\V1/V2/V1/V2/w3 ),
    .ZN(\V1/V2/V1/v2 [3]));
 XOR2_X2 \V1/V2/V1/V2/HA2/_1_  (.A(\V1/V2/V1/V2/w4 ),
    .B(\V1/V2/V1/V2/w3 ),
    .Z(\V1/V2/V1/v2 [2]));
 AND2_X1 \V1/V2/V1/V2/_0_  (.A1(A[10]),
    .A2(B[0]),
    .ZN(\V1/V2/V1/v2 [0]));
 AND2_X1 \V1/V2/V1/V2/_1_  (.A1(A[10]),
    .A2(B[1]),
    .ZN(\V1/V2/V1/V2/w1 ));
 AND2_X1 \V1/V2/V1/V2/_2_  (.A1(B[0]),
    .A2(A[11]),
    .ZN(\V1/V2/V1/V2/w2 ));
 AND2_X1 \V1/V2/V1/V2/_3_  (.A1(B[1]),
    .A2(A[11]),
    .ZN(\V1/V2/V1/V2/w3 ));
 AND2_X1 \V1/V2/V1/V3/HA1/_0_  (.A1(\V1/V2/V1/V3/w2 ),
    .A2(\V1/V2/V1/V3/w1 ),
    .ZN(\V1/V2/V1/V3/w4 ));
 XOR2_X2 \V1/V2/V1/V3/HA1/_1_  (.A(\V1/V2/V1/V3/w2 ),
    .B(\V1/V2/V1/V3/w1 ),
    .Z(\V1/V2/V1/v3 [1]));
 AND2_X1 \V1/V2/V1/V3/HA2/_0_  (.A1(\V1/V2/V1/V3/w4 ),
    .A2(\V1/V2/V1/V3/w3 ),
    .ZN(\V1/V2/V1/v3 [3]));
 XOR2_X2 \V1/V2/V1/V3/HA2/_1_  (.A(\V1/V2/V1/V3/w4 ),
    .B(\V1/V2/V1/V3/w3 ),
    .Z(\V1/V2/V1/v3 [2]));
 AND2_X1 \V1/V2/V1/V3/_0_  (.A1(A[8]),
    .A2(B[2]),
    .ZN(\V1/V2/V1/v3 [0]));
 AND2_X1 \V1/V2/V1/V3/_1_  (.A1(A[8]),
    .A2(B[3]),
    .ZN(\V1/V2/V1/V3/w1 ));
 AND2_X1 \V1/V2/V1/V3/_2_  (.A1(B[2]),
    .A2(A[9]),
    .ZN(\V1/V2/V1/V3/w2 ));
 AND2_X1 \V1/V2/V1/V3/_3_  (.A1(B[3]),
    .A2(A[9]),
    .ZN(\V1/V2/V1/V3/w3 ));
 AND2_X1 \V1/V2/V1/V4/HA1/_0_  (.A1(\V1/V2/V1/V4/w2 ),
    .A2(\V1/V2/V1/V4/w1 ),
    .ZN(\V1/V2/V1/V4/w4 ));
 XOR2_X2 \V1/V2/V1/V4/HA1/_1_  (.A(\V1/V2/V1/V4/w2 ),
    .B(\V1/V2/V1/V4/w1 ),
    .Z(\V1/V2/V1/v4 [1]));
 AND2_X1 \V1/V2/V1/V4/HA2/_0_  (.A1(\V1/V2/V1/V4/w4 ),
    .A2(\V1/V2/V1/V4/w3 ),
    .ZN(\V1/V2/V1/v4 [3]));
 XOR2_X2 \V1/V2/V1/V4/HA2/_1_  (.A(\V1/V2/V1/V4/w4 ),
    .B(\V1/V2/V1/V4/w3 ),
    .Z(\V1/V2/V1/v4 [2]));
 AND2_X1 \V1/V2/V1/V4/_0_  (.A1(A[10]),
    .A2(B[2]),
    .ZN(\V1/V2/V1/v4 [0]));
 AND2_X1 \V1/V2/V1/V4/_1_  (.A1(A[10]),
    .A2(B[3]),
    .ZN(\V1/V2/V1/V4/w1 ));
 AND2_X1 \V1/V2/V1/V4/_2_  (.A1(B[2]),
    .A2(A[11]),
    .ZN(\V1/V2/V1/V4/w2 ));
 AND2_X1 \V1/V2/V1/V4/_3_  (.A1(B[3]),
    .A2(A[11]),
    .ZN(\V1/V2/V1/V4/w3 ));
 OR2_X2 \V1/V2/V1/_0_  (.A1(\V1/V2/V1/c1 ),
    .A2(\V1/V2/V1/c2 ),
    .ZN(\V1/V2/V1/c3 ));
 AND2_X1 \V1/V2/V2/A1/M1/M1/_0_  (.A1(\V1/V2/V2/v2 [0]),
    .A2(\V1/V2/V2/v3 [0]),
    .ZN(\V1/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M1/M1/_1_  (.A(\V1/V2/V2/v2 [0]),
    .B(\V1/V2/V2/v3 [0]),
    .Z(\V1/V2/V2/A1/M1/s1 ));
 AND2_X1 \V1/V2/V2/A1/M1/M2/_0_  (.A1(\V1/V2/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M1/M2/_1_  (.A(\V1/V2/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/V2/s1 [0]));
 OR2_X1 \V1/V2/V2/A1/M1/_0_  (.A1(\V1/V2/V2/A1/M1/c1 ),
    .A2(\V1/V2/V2/A1/M1/c2 ),
    .ZN(\V1/V2/V2/A1/c1 ));
 AND2_X1 \V1/V2/V2/A1/M2/M1/_0_  (.A1(\V1/V2/V2/v2 [1]),
    .A2(\V1/V2/V2/v3 [1]),
    .ZN(\V1/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M2/M1/_1_  (.A(\V1/V2/V2/v2 [1]),
    .B(\V1/V2/V2/v3 [1]),
    .Z(\V1/V2/V2/A1/M2/s1 ));
 AND2_X1 \V1/V2/V2/A1/M2/M2/_0_  (.A1(\V1/V2/V2/A1/M2/s1 ),
    .A2(\V1/V2/V2/A1/c1 ),
    .ZN(\V1/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M2/M2/_1_  (.A(\V1/V2/V2/A1/M2/s1 ),
    .B(\V1/V2/V2/A1/c1 ),
    .Z(\V1/V2/V2/s1 [1]));
 OR2_X1 \V1/V2/V2/A1/M2/_0_  (.A1(\V1/V2/V2/A1/M2/c1 ),
    .A2(\V1/V2/V2/A1/M2/c2 ),
    .ZN(\V1/V2/V2/A1/c2 ));
 AND2_X1 \V1/V2/V2/A1/M3/M1/_0_  (.A1(\V1/V2/V2/v2 [2]),
    .A2(\V1/V2/V2/v3 [2]),
    .ZN(\V1/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M3/M1/_1_  (.A(\V1/V2/V2/v2 [2]),
    .B(\V1/V2/V2/v3 [2]),
    .Z(\V1/V2/V2/A1/M3/s1 ));
 AND2_X1 \V1/V2/V2/A1/M3/M2/_0_  (.A1(\V1/V2/V2/A1/M3/s1 ),
    .A2(\V1/V2/V2/A1/c2 ),
    .ZN(\V1/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M3/M2/_1_  (.A(\V1/V2/V2/A1/M3/s1 ),
    .B(\V1/V2/V2/A1/c2 ),
    .Z(\V1/V2/V2/s1 [2]));
 OR2_X1 \V1/V2/V2/A1/M3/_0_  (.A1(\V1/V2/V2/A1/M3/c1 ),
    .A2(\V1/V2/V2/A1/M3/c2 ),
    .ZN(\V1/V2/V2/A1/c3 ));
 AND2_X1 \V1/V2/V2/A1/M4/M1/_0_  (.A1(\V1/V2/V2/v2 [3]),
    .A2(\V1/V2/V2/v3 [3]),
    .ZN(\V1/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M4/M1/_1_  (.A(\V1/V2/V2/v2 [3]),
    .B(\V1/V2/V2/v3 [3]),
    .Z(\V1/V2/V2/A1/M4/s1 ));
 AND2_X1 \V1/V2/V2/A1/M4/M2/_0_  (.A1(\V1/V2/V2/A1/M4/s1 ),
    .A2(\V1/V2/V2/A1/c3 ),
    .ZN(\V1/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M4/M2/_1_  (.A(\V1/V2/V2/A1/M4/s1 ),
    .B(\V1/V2/V2/A1/c3 ),
    .Z(\V1/V2/V2/s1 [3]));
 OR2_X1 \V1/V2/V2/A1/M4/_0_  (.A1(\V1/V2/V2/A1/M4/c1 ),
    .A2(\V1/V2/V2/A1/M4/c2 ),
    .ZN(\V1/V2/V2/c1 ));
 AND2_X1 \V1/V2/V2/A2/M1/M1/_0_  (.A1(\V1/V2/V2/s1 [0]),
    .A2(\V1/V2/V2/v1 [2]),
    .ZN(\V1/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M1/M1/_1_  (.A(\V1/V2/V2/s1 [0]),
    .B(\V1/V2/V2/v1 [2]),
    .Z(\V1/V2/V2/A2/M1/s1 ));
 AND2_X1 \V1/V2/V2/A2/M1/M2/_0_  (.A1(\V1/V2/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M1/M2/_1_  (.A(\V1/V2/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v2 [2]));
 OR2_X1 \V1/V2/V2/A2/M1/_0_  (.A1(\V1/V2/V2/A2/M1/c1 ),
    .A2(\V1/V2/V2/A2/M1/c2 ),
    .ZN(\V1/V2/V2/A2/c1 ));
 AND2_X1 \V1/V2/V2/A2/M2/M1/_0_  (.A1(\V1/V2/V2/s1 [1]),
    .A2(\V1/V2/V2/v1 [3]),
    .ZN(\V1/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M2/M1/_1_  (.A(\V1/V2/V2/s1 [1]),
    .B(\V1/V2/V2/v1 [3]),
    .Z(\V1/V2/V2/A2/M2/s1 ));
 AND2_X1 \V1/V2/V2/A2/M2/M2/_0_  (.A1(\V1/V2/V2/A2/M2/s1 ),
    .A2(\V1/V2/V2/A2/c1 ),
    .ZN(\V1/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M2/M2/_1_  (.A(\V1/V2/V2/A2/M2/s1 ),
    .B(\V1/V2/V2/A2/c1 ),
    .Z(\V1/V2/v2 [3]));
 OR2_X1 \V1/V2/V2/A2/M2/_0_  (.A1(\V1/V2/V2/A2/M2/c1 ),
    .A2(\V1/V2/V2/A2/M2/c2 ),
    .ZN(\V1/V2/V2/A2/c2 ));
 AND2_X1 \V1/V2/V2/A2/M3/M1/_0_  (.A1(\V1/V2/V2/s1 [2]),
    .A2(ground),
    .ZN(\V1/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M3/M1/_1_  (.A(\V1/V2/V2/s1 [2]),
    .B(ground),
    .Z(\V1/V2/V2/A2/M3/s1 ));
 AND2_X1 \V1/V2/V2/A2/M3/M2/_0_  (.A1(\V1/V2/V2/A2/M3/s1 ),
    .A2(\V1/V2/V2/A2/c2 ),
    .ZN(\V1/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M3/M2/_1_  (.A(\V1/V2/V2/A2/M3/s1 ),
    .B(\V1/V2/V2/A2/c2 ),
    .Z(\V1/V2/V2/s2 [2]));
 OR2_X1 \V1/V2/V2/A2/M3/_0_  (.A1(\V1/V2/V2/A2/M3/c1 ),
    .A2(\V1/V2/V2/A2/M3/c2 ),
    .ZN(\V1/V2/V2/A2/c3 ));
 AND2_X1 \V1/V2/V2/A2/M4/M1/_0_  (.A1(\V1/V2/V2/s1 [3]),
    .A2(ground),
    .ZN(\V1/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M4/M1/_1_  (.A(\V1/V2/V2/s1 [3]),
    .B(ground),
    .Z(\V1/V2/V2/A2/M4/s1 ));
 AND2_X1 \V1/V2/V2/A2/M4/M2/_0_  (.A1(\V1/V2/V2/A2/M4/s1 ),
    .A2(\V1/V2/V2/A2/c3 ),
    .ZN(\V1/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M4/M2/_1_  (.A(\V1/V2/V2/A2/M4/s1 ),
    .B(\V1/V2/V2/A2/c3 ),
    .Z(\V1/V2/V2/s2 [3]));
 OR2_X1 \V1/V2/V2/A2/M4/_0_  (.A1(\V1/V2/V2/A2/M4/c1 ),
    .A2(\V1/V2/V2/A2/M4/c2 ),
    .ZN(\V1/V2/V2/c2 ));
 AND2_X1 \V1/V2/V2/A3/M1/M1/_0_  (.A1(\V1/V2/V2/v4 [0]),
    .A2(\V1/V2/V2/s2 [2]),
    .ZN(\V1/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M1/M1/_1_  (.A(\V1/V2/V2/v4 [0]),
    .B(\V1/V2/V2/s2 [2]),
    .Z(\V1/V2/V2/A3/M1/s1 ));
 AND2_X1 \V1/V2/V2/A3/M1/M2/_0_  (.A1(\V1/V2/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M1/M2/_1_  (.A(\V1/V2/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v2 [4]));
 OR2_X1 \V1/V2/V2/A3/M1/_0_  (.A1(\V1/V2/V2/A3/M1/c1 ),
    .A2(\V1/V2/V2/A3/M1/c2 ),
    .ZN(\V1/V2/V2/A3/c1 ));
 AND2_X1 \V1/V2/V2/A3/M2/M1/_0_  (.A1(\V1/V2/V2/v4 [1]),
    .A2(\V1/V2/V2/s2 [3]),
    .ZN(\V1/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M2/M1/_1_  (.A(\V1/V2/V2/v4 [1]),
    .B(\V1/V2/V2/s2 [3]),
    .Z(\V1/V2/V2/A3/M2/s1 ));
 AND2_X1 \V1/V2/V2/A3/M2/M2/_0_  (.A1(\V1/V2/V2/A3/M2/s1 ),
    .A2(\V1/V2/V2/A3/c1 ),
    .ZN(\V1/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M2/M2/_1_  (.A(\V1/V2/V2/A3/M2/s1 ),
    .B(\V1/V2/V2/A3/c1 ),
    .Z(\V1/V2/v2 [5]));
 OR2_X1 \V1/V2/V2/A3/M2/_0_  (.A1(\V1/V2/V2/A3/M2/c1 ),
    .A2(\V1/V2/V2/A3/M2/c2 ),
    .ZN(\V1/V2/V2/A3/c2 ));
 AND2_X1 \V1/V2/V2/A3/M3/M1/_0_  (.A1(\V1/V2/V2/v4 [2]),
    .A2(\V1/V2/V2/c3 ),
    .ZN(\V1/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M3/M1/_1_  (.A(\V1/V2/V2/v4 [2]),
    .B(\V1/V2/V2/c3 ),
    .Z(\V1/V2/V2/A3/M3/s1 ));
 AND2_X1 \V1/V2/V2/A3/M3/M2/_0_  (.A1(\V1/V2/V2/A3/M3/s1 ),
    .A2(\V1/V2/V2/A3/c2 ),
    .ZN(\V1/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M3/M2/_1_  (.A(\V1/V2/V2/A3/M3/s1 ),
    .B(\V1/V2/V2/A3/c2 ),
    .Z(\V1/V2/v2 [6]));
 OR2_X1 \V1/V2/V2/A3/M3/_0_  (.A1(\V1/V2/V2/A3/M3/c1 ),
    .A2(\V1/V2/V2/A3/M3/c2 ),
    .ZN(\V1/V2/V2/A3/c3 ));
 AND2_X1 \V1/V2/V2/A3/M4/M1/_0_  (.A1(\V1/V2/V2/v4 [3]),
    .A2(ground),
    .ZN(\V1/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M4/M1/_1_  (.A(\V1/V2/V2/v4 [3]),
    .B(ground),
    .Z(\V1/V2/V2/A3/M4/s1 ));
 AND2_X1 \V1/V2/V2/A3/M4/M2/_0_  (.A1(\V1/V2/V2/A3/M4/s1 ),
    .A2(\V1/V2/V2/A3/c3 ),
    .ZN(\V1/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M4/M2/_1_  (.A(\V1/V2/V2/A3/M4/s1 ),
    .B(\V1/V2/V2/A3/c3 ),
    .Z(\V1/V2/v2 [7]));
 OR2_X1 \V1/V2/V2/A3/M4/_0_  (.A1(\V1/V2/V2/A3/M4/c1 ),
    .A2(\V1/V2/V2/A3/M4/c2 ),
    .ZN(\V1/V2/V2/overflow ));
 AND2_X1 \V1/V2/V2/V1/HA1/_0_  (.A1(\V1/V2/V2/V1/w2 ),
    .A2(\V1/V2/V2/V1/w1 ),
    .ZN(\V1/V2/V2/V1/w4 ));
 XOR2_X2 \V1/V2/V2/V1/HA1/_1_  (.A(\V1/V2/V2/V1/w2 ),
    .B(\V1/V2/V2/V1/w1 ),
    .Z(\V1/V2/v2 [1]));
 AND2_X1 \V1/V2/V2/V1/HA2/_0_  (.A1(\V1/V2/V2/V1/w4 ),
    .A2(\V1/V2/V2/V1/w3 ),
    .ZN(\V1/V2/V2/v1 [3]));
 XOR2_X2 \V1/V2/V2/V1/HA2/_1_  (.A(\V1/V2/V2/V1/w4 ),
    .B(\V1/V2/V2/V1/w3 ),
    .Z(\V1/V2/V2/v1 [2]));
 AND2_X1 \V1/V2/V2/V1/_0_  (.A1(A[12]),
    .A2(B[0]),
    .ZN(\V1/V2/v2 [0]));
 AND2_X1 \V1/V2/V2/V1/_1_  (.A1(A[12]),
    .A2(B[1]),
    .ZN(\V1/V2/V2/V1/w1 ));
 AND2_X1 \V1/V2/V2/V1/_2_  (.A1(B[0]),
    .A2(A[13]),
    .ZN(\V1/V2/V2/V1/w2 ));
 AND2_X1 \V1/V2/V2/V1/_3_  (.A1(B[1]),
    .A2(A[13]),
    .ZN(\V1/V2/V2/V1/w3 ));
 AND2_X1 \V1/V2/V2/V2/HA1/_0_  (.A1(\V1/V2/V2/V2/w2 ),
    .A2(\V1/V2/V2/V2/w1 ),
    .ZN(\V1/V2/V2/V2/w4 ));
 XOR2_X2 \V1/V2/V2/V2/HA1/_1_  (.A(\V1/V2/V2/V2/w2 ),
    .B(\V1/V2/V2/V2/w1 ),
    .Z(\V1/V2/V2/v2 [1]));
 AND2_X1 \V1/V2/V2/V2/HA2/_0_  (.A1(\V1/V2/V2/V2/w4 ),
    .A2(\V1/V2/V2/V2/w3 ),
    .ZN(\V1/V2/V2/v2 [3]));
 XOR2_X2 \V1/V2/V2/V2/HA2/_1_  (.A(\V1/V2/V2/V2/w4 ),
    .B(\V1/V2/V2/V2/w3 ),
    .Z(\V1/V2/V2/v2 [2]));
 AND2_X1 \V1/V2/V2/V2/_0_  (.A1(A[14]),
    .A2(B[0]),
    .ZN(\V1/V2/V2/v2 [0]));
 AND2_X1 \V1/V2/V2/V2/_1_  (.A1(A[14]),
    .A2(B[1]),
    .ZN(\V1/V2/V2/V2/w1 ));
 AND2_X1 \V1/V2/V2/V2/_2_  (.A1(B[0]),
    .A2(A[15]),
    .ZN(\V1/V2/V2/V2/w2 ));
 AND2_X1 \V1/V2/V2/V2/_3_  (.A1(B[1]),
    .A2(A[15]),
    .ZN(\V1/V2/V2/V2/w3 ));
 AND2_X1 \V1/V2/V2/V3/HA1/_0_  (.A1(\V1/V2/V2/V3/w2 ),
    .A2(\V1/V2/V2/V3/w1 ),
    .ZN(\V1/V2/V2/V3/w4 ));
 XOR2_X2 \V1/V2/V2/V3/HA1/_1_  (.A(\V1/V2/V2/V3/w2 ),
    .B(\V1/V2/V2/V3/w1 ),
    .Z(\V1/V2/V2/v3 [1]));
 AND2_X1 \V1/V2/V2/V3/HA2/_0_  (.A1(\V1/V2/V2/V3/w4 ),
    .A2(\V1/V2/V2/V3/w3 ),
    .ZN(\V1/V2/V2/v3 [3]));
 XOR2_X2 \V1/V2/V2/V3/HA2/_1_  (.A(\V1/V2/V2/V3/w4 ),
    .B(\V1/V2/V2/V3/w3 ),
    .Z(\V1/V2/V2/v3 [2]));
 AND2_X1 \V1/V2/V2/V3/_0_  (.A1(A[12]),
    .A2(B[2]),
    .ZN(\V1/V2/V2/v3 [0]));
 AND2_X1 \V1/V2/V2/V3/_1_  (.A1(A[12]),
    .A2(B[3]),
    .ZN(\V1/V2/V2/V3/w1 ));
 AND2_X1 \V1/V2/V2/V3/_2_  (.A1(B[2]),
    .A2(A[13]),
    .ZN(\V1/V2/V2/V3/w2 ));
 AND2_X1 \V1/V2/V2/V3/_3_  (.A1(B[3]),
    .A2(A[13]),
    .ZN(\V1/V2/V2/V3/w3 ));
 AND2_X1 \V1/V2/V2/V4/HA1/_0_  (.A1(\V1/V2/V2/V4/w2 ),
    .A2(\V1/V2/V2/V4/w1 ),
    .ZN(\V1/V2/V2/V4/w4 ));
 XOR2_X2 \V1/V2/V2/V4/HA1/_1_  (.A(\V1/V2/V2/V4/w2 ),
    .B(\V1/V2/V2/V4/w1 ),
    .Z(\V1/V2/V2/v4 [1]));
 AND2_X1 \V1/V2/V2/V4/HA2/_0_  (.A1(\V1/V2/V2/V4/w4 ),
    .A2(\V1/V2/V2/V4/w3 ),
    .ZN(\V1/V2/V2/v4 [3]));
 XOR2_X2 \V1/V2/V2/V4/HA2/_1_  (.A(\V1/V2/V2/V4/w4 ),
    .B(\V1/V2/V2/V4/w3 ),
    .Z(\V1/V2/V2/v4 [2]));
 AND2_X1 \V1/V2/V2/V4/_0_  (.A1(A[14]),
    .A2(B[2]),
    .ZN(\V1/V2/V2/v4 [0]));
 AND2_X1 \V1/V2/V2/V4/_1_  (.A1(A[14]),
    .A2(B[3]),
    .ZN(\V1/V2/V2/V4/w1 ));
 AND2_X1 \V1/V2/V2/V4/_2_  (.A1(B[2]),
    .A2(A[15]),
    .ZN(\V1/V2/V2/V4/w2 ));
 AND2_X1 \V1/V2/V2/V4/_3_  (.A1(B[3]),
    .A2(A[15]),
    .ZN(\V1/V2/V2/V4/w3 ));
 OR2_X1 \V1/V2/V2/_0_  (.A1(\V1/V2/V2/c1 ),
    .A2(\V1/V2/V2/c2 ),
    .ZN(\V1/V2/V2/c3 ));
 AND2_X1 \V1/V2/V3/A1/M1/M1/_0_  (.A1(\V1/V2/V3/v2 [0]),
    .A2(\V1/V2/V3/v3 [0]),
    .ZN(\V1/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M1/M1/_1_  (.A(\V1/V2/V3/v2 [0]),
    .B(\V1/V2/V3/v3 [0]),
    .Z(\V1/V2/V3/A1/M1/s1 ));
 AND2_X1 \V1/V2/V3/A1/M1/M2/_0_  (.A1(\V1/V2/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M1/M2/_1_  (.A(\V1/V2/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/V3/s1 [0]));
 OR2_X1 \V1/V2/V3/A1/M1/_0_  (.A1(\V1/V2/V3/A1/M1/c1 ),
    .A2(\V1/V2/V3/A1/M1/c2 ),
    .ZN(\V1/V2/V3/A1/c1 ));
 AND2_X1 \V1/V2/V3/A1/M2/M1/_0_  (.A1(\V1/V2/V3/v2 [1]),
    .A2(\V1/V2/V3/v3 [1]),
    .ZN(\V1/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M2/M1/_1_  (.A(\V1/V2/V3/v2 [1]),
    .B(\V1/V2/V3/v3 [1]),
    .Z(\V1/V2/V3/A1/M2/s1 ));
 AND2_X1 \V1/V2/V3/A1/M2/M2/_0_  (.A1(\V1/V2/V3/A1/M2/s1 ),
    .A2(\V1/V2/V3/A1/c1 ),
    .ZN(\V1/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M2/M2/_1_  (.A(\V1/V2/V3/A1/M2/s1 ),
    .B(\V1/V2/V3/A1/c1 ),
    .Z(\V1/V2/V3/s1 [1]));
 OR2_X1 \V1/V2/V3/A1/M2/_0_  (.A1(\V1/V2/V3/A1/M2/c1 ),
    .A2(\V1/V2/V3/A1/M2/c2 ),
    .ZN(\V1/V2/V3/A1/c2 ));
 AND2_X1 \V1/V2/V3/A1/M3/M1/_0_  (.A1(\V1/V2/V3/v2 [2]),
    .A2(\V1/V2/V3/v3 [2]),
    .ZN(\V1/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M3/M1/_1_  (.A(\V1/V2/V3/v2 [2]),
    .B(\V1/V2/V3/v3 [2]),
    .Z(\V1/V2/V3/A1/M3/s1 ));
 AND2_X1 \V1/V2/V3/A1/M3/M2/_0_  (.A1(\V1/V2/V3/A1/M3/s1 ),
    .A2(\V1/V2/V3/A1/c2 ),
    .ZN(\V1/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M3/M2/_1_  (.A(\V1/V2/V3/A1/M3/s1 ),
    .B(\V1/V2/V3/A1/c2 ),
    .Z(\V1/V2/V3/s1 [2]));
 OR2_X1 \V1/V2/V3/A1/M3/_0_  (.A1(\V1/V2/V3/A1/M3/c1 ),
    .A2(\V1/V2/V3/A1/M3/c2 ),
    .ZN(\V1/V2/V3/A1/c3 ));
 AND2_X1 \V1/V2/V3/A1/M4/M1/_0_  (.A1(\V1/V2/V3/v2 [3]),
    .A2(\V1/V2/V3/v3 [3]),
    .ZN(\V1/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M4/M1/_1_  (.A(\V1/V2/V3/v2 [3]),
    .B(\V1/V2/V3/v3 [3]),
    .Z(\V1/V2/V3/A1/M4/s1 ));
 AND2_X1 \V1/V2/V3/A1/M4/M2/_0_  (.A1(\V1/V2/V3/A1/M4/s1 ),
    .A2(\V1/V2/V3/A1/c3 ),
    .ZN(\V1/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M4/M2/_1_  (.A(\V1/V2/V3/A1/M4/s1 ),
    .B(\V1/V2/V3/A1/c3 ),
    .Z(\V1/V2/V3/s1 [3]));
 OR2_X1 \V1/V2/V3/A1/M4/_0_  (.A1(\V1/V2/V3/A1/M4/c1 ),
    .A2(\V1/V2/V3/A1/M4/c2 ),
    .ZN(\V1/V2/V3/c1 ));
 AND2_X1 \V1/V2/V3/A2/M1/M1/_0_  (.A1(\V1/V2/V3/s1 [0]),
    .A2(\V1/V2/V3/v1 [2]),
    .ZN(\V1/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M1/M1/_1_  (.A(\V1/V2/V3/s1 [0]),
    .B(\V1/V2/V3/v1 [2]),
    .Z(\V1/V2/V3/A2/M1/s1 ));
 AND2_X1 \V1/V2/V3/A2/M1/M2/_0_  (.A1(\V1/V2/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M1/M2/_1_  (.A(\V1/V2/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v3 [2]));
 OR2_X1 \V1/V2/V3/A2/M1/_0_  (.A1(\V1/V2/V3/A2/M1/c1 ),
    .A2(\V1/V2/V3/A2/M1/c2 ),
    .ZN(\V1/V2/V3/A2/c1 ));
 AND2_X1 \V1/V2/V3/A2/M2/M1/_0_  (.A1(\V1/V2/V3/s1 [1]),
    .A2(\V1/V2/V3/v1 [3]),
    .ZN(\V1/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M2/M1/_1_  (.A(\V1/V2/V3/s1 [1]),
    .B(\V1/V2/V3/v1 [3]),
    .Z(\V1/V2/V3/A2/M2/s1 ));
 AND2_X1 \V1/V2/V3/A2/M2/M2/_0_  (.A1(\V1/V2/V3/A2/M2/s1 ),
    .A2(\V1/V2/V3/A2/c1 ),
    .ZN(\V1/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M2/M2/_1_  (.A(\V1/V2/V3/A2/M2/s1 ),
    .B(\V1/V2/V3/A2/c1 ),
    .Z(\V1/V2/v3 [3]));
 OR2_X1 \V1/V2/V3/A2/M2/_0_  (.A1(\V1/V2/V3/A2/M2/c1 ),
    .A2(\V1/V2/V3/A2/M2/c2 ),
    .ZN(\V1/V2/V3/A2/c2 ));
 AND2_X1 \V1/V2/V3/A2/M3/M1/_0_  (.A1(\V1/V2/V3/s1 [2]),
    .A2(ground),
    .ZN(\V1/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M3/M1/_1_  (.A(\V1/V2/V3/s1 [2]),
    .B(ground),
    .Z(\V1/V2/V3/A2/M3/s1 ));
 AND2_X1 \V1/V2/V3/A2/M3/M2/_0_  (.A1(\V1/V2/V3/A2/M3/s1 ),
    .A2(\V1/V2/V3/A2/c2 ),
    .ZN(\V1/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M3/M2/_1_  (.A(\V1/V2/V3/A2/M3/s1 ),
    .B(\V1/V2/V3/A2/c2 ),
    .Z(\V1/V2/V3/s2 [2]));
 OR2_X1 \V1/V2/V3/A2/M3/_0_  (.A1(\V1/V2/V3/A2/M3/c1 ),
    .A2(\V1/V2/V3/A2/M3/c2 ),
    .ZN(\V1/V2/V3/A2/c3 ));
 AND2_X1 \V1/V2/V3/A2/M4/M1/_0_  (.A1(\V1/V2/V3/s1 [3]),
    .A2(ground),
    .ZN(\V1/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M4/M1/_1_  (.A(\V1/V2/V3/s1 [3]),
    .B(ground),
    .Z(\V1/V2/V3/A2/M4/s1 ));
 AND2_X1 \V1/V2/V3/A2/M4/M2/_0_  (.A1(\V1/V2/V3/A2/M4/s1 ),
    .A2(\V1/V2/V3/A2/c3 ),
    .ZN(\V1/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M4/M2/_1_  (.A(\V1/V2/V3/A2/M4/s1 ),
    .B(\V1/V2/V3/A2/c3 ),
    .Z(\V1/V2/V3/s2 [3]));
 OR2_X1 \V1/V2/V3/A2/M4/_0_  (.A1(\V1/V2/V3/A2/M4/c1 ),
    .A2(\V1/V2/V3/A2/M4/c2 ),
    .ZN(\V1/V2/V3/c2 ));
 AND2_X1 \V1/V2/V3/A3/M1/M1/_0_  (.A1(\V1/V2/V3/v4 [0]),
    .A2(\V1/V2/V3/s2 [2]),
    .ZN(\V1/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M1/M1/_1_  (.A(\V1/V2/V3/v4 [0]),
    .B(\V1/V2/V3/s2 [2]),
    .Z(\V1/V2/V3/A3/M1/s1 ));
 AND2_X1 \V1/V2/V3/A3/M1/M2/_0_  (.A1(\V1/V2/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M1/M2/_1_  (.A(\V1/V2/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v3 [4]));
 OR2_X1 \V1/V2/V3/A3/M1/_0_  (.A1(\V1/V2/V3/A3/M1/c1 ),
    .A2(\V1/V2/V3/A3/M1/c2 ),
    .ZN(\V1/V2/V3/A3/c1 ));
 AND2_X1 \V1/V2/V3/A3/M2/M1/_0_  (.A1(\V1/V2/V3/v4 [1]),
    .A2(\V1/V2/V3/s2 [3]),
    .ZN(\V1/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M2/M1/_1_  (.A(\V1/V2/V3/v4 [1]),
    .B(\V1/V2/V3/s2 [3]),
    .Z(\V1/V2/V3/A3/M2/s1 ));
 AND2_X1 \V1/V2/V3/A3/M2/M2/_0_  (.A1(\V1/V2/V3/A3/M2/s1 ),
    .A2(\V1/V2/V3/A3/c1 ),
    .ZN(\V1/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M2/M2/_1_  (.A(\V1/V2/V3/A3/M2/s1 ),
    .B(\V1/V2/V3/A3/c1 ),
    .Z(\V1/V2/v3 [5]));
 OR2_X1 \V1/V2/V3/A3/M2/_0_  (.A1(\V1/V2/V3/A3/M2/c1 ),
    .A2(\V1/V2/V3/A3/M2/c2 ),
    .ZN(\V1/V2/V3/A3/c2 ));
 AND2_X1 \V1/V2/V3/A3/M3/M1/_0_  (.A1(\V1/V2/V3/v4 [2]),
    .A2(\V1/V2/V3/c3 ),
    .ZN(\V1/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M3/M1/_1_  (.A(\V1/V2/V3/v4 [2]),
    .B(\V1/V2/V3/c3 ),
    .Z(\V1/V2/V3/A3/M3/s1 ));
 AND2_X1 \V1/V2/V3/A3/M3/M2/_0_  (.A1(\V1/V2/V3/A3/M3/s1 ),
    .A2(\V1/V2/V3/A3/c2 ),
    .ZN(\V1/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M3/M2/_1_  (.A(\V1/V2/V3/A3/M3/s1 ),
    .B(\V1/V2/V3/A3/c2 ),
    .Z(\V1/V2/v3 [6]));
 OR2_X1 \V1/V2/V3/A3/M3/_0_  (.A1(\V1/V2/V3/A3/M3/c1 ),
    .A2(\V1/V2/V3/A3/M3/c2 ),
    .ZN(\V1/V2/V3/A3/c3 ));
 AND2_X1 \V1/V2/V3/A3/M4/M1/_0_  (.A1(\V1/V2/V3/v4 [3]),
    .A2(ground),
    .ZN(\V1/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M4/M1/_1_  (.A(\V1/V2/V3/v4 [3]),
    .B(ground),
    .Z(\V1/V2/V3/A3/M4/s1 ));
 AND2_X1 \V1/V2/V3/A3/M4/M2/_0_  (.A1(\V1/V2/V3/A3/M4/s1 ),
    .A2(\V1/V2/V3/A3/c3 ),
    .ZN(\V1/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M4/M2/_1_  (.A(\V1/V2/V3/A3/M4/s1 ),
    .B(\V1/V2/V3/A3/c3 ),
    .Z(\V1/V2/v3 [7]));
 OR2_X1 \V1/V2/V3/A3/M4/_0_  (.A1(\V1/V2/V3/A3/M4/c1 ),
    .A2(\V1/V2/V3/A3/M4/c2 ),
    .ZN(\V1/V2/V3/overflow ));
 AND2_X1 \V1/V2/V3/V1/HA1/_0_  (.A1(\V1/V2/V3/V1/w2 ),
    .A2(\V1/V2/V3/V1/w1 ),
    .ZN(\V1/V2/V3/V1/w4 ));
 XOR2_X2 \V1/V2/V3/V1/HA1/_1_  (.A(\V1/V2/V3/V1/w2 ),
    .B(\V1/V2/V3/V1/w1 ),
    .Z(\V1/V2/v3 [1]));
 AND2_X1 \V1/V2/V3/V1/HA2/_0_  (.A1(\V1/V2/V3/V1/w4 ),
    .A2(\V1/V2/V3/V1/w3 ),
    .ZN(\V1/V2/V3/v1 [3]));
 XOR2_X2 \V1/V2/V3/V1/HA2/_1_  (.A(\V1/V2/V3/V1/w4 ),
    .B(\V1/V2/V3/V1/w3 ),
    .Z(\V1/V2/V3/v1 [2]));
 AND2_X1 \V1/V2/V3/V1/_0_  (.A1(A[8]),
    .A2(B[4]),
    .ZN(\V1/V2/v3 [0]));
 AND2_X1 \V1/V2/V3/V1/_1_  (.A1(A[8]),
    .A2(B[5]),
    .ZN(\V1/V2/V3/V1/w1 ));
 AND2_X1 \V1/V2/V3/V1/_2_  (.A1(B[4]),
    .A2(A[9]),
    .ZN(\V1/V2/V3/V1/w2 ));
 AND2_X1 \V1/V2/V3/V1/_3_  (.A1(B[5]),
    .A2(A[9]),
    .ZN(\V1/V2/V3/V1/w3 ));
 AND2_X1 \V1/V2/V3/V2/HA1/_0_  (.A1(\V1/V2/V3/V2/w2 ),
    .A2(\V1/V2/V3/V2/w1 ),
    .ZN(\V1/V2/V3/V2/w4 ));
 XOR2_X2 \V1/V2/V3/V2/HA1/_1_  (.A(\V1/V2/V3/V2/w2 ),
    .B(\V1/V2/V3/V2/w1 ),
    .Z(\V1/V2/V3/v2 [1]));
 AND2_X1 \V1/V2/V3/V2/HA2/_0_  (.A1(\V1/V2/V3/V2/w4 ),
    .A2(\V1/V2/V3/V2/w3 ),
    .ZN(\V1/V2/V3/v2 [3]));
 XOR2_X2 \V1/V2/V3/V2/HA2/_1_  (.A(\V1/V2/V3/V2/w4 ),
    .B(\V1/V2/V3/V2/w3 ),
    .Z(\V1/V2/V3/v2 [2]));
 AND2_X1 \V1/V2/V3/V2/_0_  (.A1(A[10]),
    .A2(B[4]),
    .ZN(\V1/V2/V3/v2 [0]));
 AND2_X1 \V1/V2/V3/V2/_1_  (.A1(A[10]),
    .A2(B[5]),
    .ZN(\V1/V2/V3/V2/w1 ));
 AND2_X1 \V1/V2/V3/V2/_2_  (.A1(B[4]),
    .A2(A[11]),
    .ZN(\V1/V2/V3/V2/w2 ));
 AND2_X1 \V1/V2/V3/V2/_3_  (.A1(B[5]),
    .A2(A[11]),
    .ZN(\V1/V2/V3/V2/w3 ));
 AND2_X1 \V1/V2/V3/V3/HA1/_0_  (.A1(\V1/V2/V3/V3/w2 ),
    .A2(\V1/V2/V3/V3/w1 ),
    .ZN(\V1/V2/V3/V3/w4 ));
 XOR2_X2 \V1/V2/V3/V3/HA1/_1_  (.A(\V1/V2/V3/V3/w2 ),
    .B(\V1/V2/V3/V3/w1 ),
    .Z(\V1/V2/V3/v3 [1]));
 AND2_X1 \V1/V2/V3/V3/HA2/_0_  (.A1(\V1/V2/V3/V3/w4 ),
    .A2(\V1/V2/V3/V3/w3 ),
    .ZN(\V1/V2/V3/v3 [3]));
 XOR2_X2 \V1/V2/V3/V3/HA2/_1_  (.A(\V1/V2/V3/V3/w4 ),
    .B(\V1/V2/V3/V3/w3 ),
    .Z(\V1/V2/V3/v3 [2]));
 AND2_X1 \V1/V2/V3/V3/_0_  (.A1(A[8]),
    .A2(B[6]),
    .ZN(\V1/V2/V3/v3 [0]));
 AND2_X1 \V1/V2/V3/V3/_1_  (.A1(A[8]),
    .A2(B[7]),
    .ZN(\V1/V2/V3/V3/w1 ));
 AND2_X1 \V1/V2/V3/V3/_2_  (.A1(B[6]),
    .A2(A[9]),
    .ZN(\V1/V2/V3/V3/w2 ));
 AND2_X1 \V1/V2/V3/V3/_3_  (.A1(B[7]),
    .A2(A[9]),
    .ZN(\V1/V2/V3/V3/w3 ));
 AND2_X1 \V1/V2/V3/V4/HA1/_0_  (.A1(\V1/V2/V3/V4/w2 ),
    .A2(\V1/V2/V3/V4/w1 ),
    .ZN(\V1/V2/V3/V4/w4 ));
 XOR2_X2 \V1/V2/V3/V4/HA1/_1_  (.A(\V1/V2/V3/V4/w2 ),
    .B(\V1/V2/V3/V4/w1 ),
    .Z(\V1/V2/V3/v4 [1]));
 AND2_X1 \V1/V2/V3/V4/HA2/_0_  (.A1(\V1/V2/V3/V4/w4 ),
    .A2(\V1/V2/V3/V4/w3 ),
    .ZN(\V1/V2/V3/v4 [3]));
 XOR2_X2 \V1/V2/V3/V4/HA2/_1_  (.A(\V1/V2/V3/V4/w4 ),
    .B(\V1/V2/V3/V4/w3 ),
    .Z(\V1/V2/V3/v4 [2]));
 AND2_X1 \V1/V2/V3/V4/_0_  (.A1(A[10]),
    .A2(B[6]),
    .ZN(\V1/V2/V3/v4 [0]));
 AND2_X1 \V1/V2/V3/V4/_1_  (.A1(A[10]),
    .A2(B[7]),
    .ZN(\V1/V2/V3/V4/w1 ));
 AND2_X1 \V1/V2/V3/V4/_2_  (.A1(B[6]),
    .A2(A[11]),
    .ZN(\V1/V2/V3/V4/w2 ));
 AND2_X1 \V1/V2/V3/V4/_3_  (.A1(B[7]),
    .A2(A[11]),
    .ZN(\V1/V2/V3/V4/w3 ));
 OR2_X1 \V1/V2/V3/_0_  (.A1(\V1/V2/V3/c1 ),
    .A2(\V1/V2/V3/c2 ),
    .ZN(\V1/V2/V3/c3 ));
 AND2_X1 \V1/V2/V4/A1/M1/M1/_0_  (.A1(\V1/V2/V4/v2 [0]),
    .A2(\V1/V2/V4/v3 [0]),
    .ZN(\V1/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M1/M1/_1_  (.A(\V1/V2/V4/v2 [0]),
    .B(\V1/V2/V4/v3 [0]),
    .Z(\V1/V2/V4/A1/M1/s1 ));
 AND2_X1 \V1/V2/V4/A1/M1/M2/_0_  (.A1(\V1/V2/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M1/M2/_1_  (.A(\V1/V2/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/V4/s1 [0]));
 OR2_X1 \V1/V2/V4/A1/M1/_0_  (.A1(\V1/V2/V4/A1/M1/c1 ),
    .A2(\V1/V2/V4/A1/M1/c2 ),
    .ZN(\V1/V2/V4/A1/c1 ));
 AND2_X1 \V1/V2/V4/A1/M2/M1/_0_  (.A1(\V1/V2/V4/v2 [1]),
    .A2(\V1/V2/V4/v3 [1]),
    .ZN(\V1/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M2/M1/_1_  (.A(\V1/V2/V4/v2 [1]),
    .B(\V1/V2/V4/v3 [1]),
    .Z(\V1/V2/V4/A1/M2/s1 ));
 AND2_X1 \V1/V2/V4/A1/M2/M2/_0_  (.A1(\V1/V2/V4/A1/M2/s1 ),
    .A2(\V1/V2/V4/A1/c1 ),
    .ZN(\V1/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M2/M2/_1_  (.A(\V1/V2/V4/A1/M2/s1 ),
    .B(\V1/V2/V4/A1/c1 ),
    .Z(\V1/V2/V4/s1 [1]));
 OR2_X1 \V1/V2/V4/A1/M2/_0_  (.A1(\V1/V2/V4/A1/M2/c1 ),
    .A2(\V1/V2/V4/A1/M2/c2 ),
    .ZN(\V1/V2/V4/A1/c2 ));
 AND2_X1 \V1/V2/V4/A1/M3/M1/_0_  (.A1(\V1/V2/V4/v2 [2]),
    .A2(\V1/V2/V4/v3 [2]),
    .ZN(\V1/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M3/M1/_1_  (.A(\V1/V2/V4/v2 [2]),
    .B(\V1/V2/V4/v3 [2]),
    .Z(\V1/V2/V4/A1/M3/s1 ));
 AND2_X1 \V1/V2/V4/A1/M3/M2/_0_  (.A1(\V1/V2/V4/A1/M3/s1 ),
    .A2(\V1/V2/V4/A1/c2 ),
    .ZN(\V1/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M3/M2/_1_  (.A(\V1/V2/V4/A1/M3/s1 ),
    .B(\V1/V2/V4/A1/c2 ),
    .Z(\V1/V2/V4/s1 [2]));
 OR2_X1 \V1/V2/V4/A1/M3/_0_  (.A1(\V1/V2/V4/A1/M3/c1 ),
    .A2(\V1/V2/V4/A1/M3/c2 ),
    .ZN(\V1/V2/V4/A1/c3 ));
 AND2_X1 \V1/V2/V4/A1/M4/M1/_0_  (.A1(\V1/V2/V4/v2 [3]),
    .A2(\V1/V2/V4/v3 [3]),
    .ZN(\V1/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M4/M1/_1_  (.A(\V1/V2/V4/v2 [3]),
    .B(\V1/V2/V4/v3 [3]),
    .Z(\V1/V2/V4/A1/M4/s1 ));
 AND2_X1 \V1/V2/V4/A1/M4/M2/_0_  (.A1(\V1/V2/V4/A1/M4/s1 ),
    .A2(\V1/V2/V4/A1/c3 ),
    .ZN(\V1/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M4/M2/_1_  (.A(\V1/V2/V4/A1/M4/s1 ),
    .B(\V1/V2/V4/A1/c3 ),
    .Z(\V1/V2/V4/s1 [3]));
 OR2_X1 \V1/V2/V4/A1/M4/_0_  (.A1(\V1/V2/V4/A1/M4/c1 ),
    .A2(\V1/V2/V4/A1/M4/c2 ),
    .ZN(\V1/V2/V4/c1 ));
 AND2_X1 \V1/V2/V4/A2/M1/M1/_0_  (.A1(\V1/V2/V4/s1 [0]),
    .A2(\V1/V2/V4/v1 [2]),
    .ZN(\V1/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M1/M1/_1_  (.A(\V1/V2/V4/s1 [0]),
    .B(\V1/V2/V4/v1 [2]),
    .Z(\V1/V2/V4/A2/M1/s1 ));
 AND2_X1 \V1/V2/V4/A2/M1/M2/_0_  (.A1(\V1/V2/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M1/M2/_1_  (.A(\V1/V2/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v4 [2]));
 OR2_X1 \V1/V2/V4/A2/M1/_0_  (.A1(\V1/V2/V4/A2/M1/c1 ),
    .A2(\V1/V2/V4/A2/M1/c2 ),
    .ZN(\V1/V2/V4/A2/c1 ));
 AND2_X1 \V1/V2/V4/A2/M2/M1/_0_  (.A1(\V1/V2/V4/s1 [1]),
    .A2(\V1/V2/V4/v1 [3]),
    .ZN(\V1/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M2/M1/_1_  (.A(\V1/V2/V4/s1 [1]),
    .B(\V1/V2/V4/v1 [3]),
    .Z(\V1/V2/V4/A2/M2/s1 ));
 AND2_X1 \V1/V2/V4/A2/M2/M2/_0_  (.A1(\V1/V2/V4/A2/M2/s1 ),
    .A2(\V1/V2/V4/A2/c1 ),
    .ZN(\V1/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M2/M2/_1_  (.A(\V1/V2/V4/A2/M2/s1 ),
    .B(\V1/V2/V4/A2/c1 ),
    .Z(\V1/V2/v4 [3]));
 OR2_X1 \V1/V2/V4/A2/M2/_0_  (.A1(\V1/V2/V4/A2/M2/c1 ),
    .A2(\V1/V2/V4/A2/M2/c2 ),
    .ZN(\V1/V2/V4/A2/c2 ));
 AND2_X1 \V1/V2/V4/A2/M3/M1/_0_  (.A1(\V1/V2/V4/s1 [2]),
    .A2(ground),
    .ZN(\V1/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M3/M1/_1_  (.A(\V1/V2/V4/s1 [2]),
    .B(ground),
    .Z(\V1/V2/V4/A2/M3/s1 ));
 AND2_X1 \V1/V2/V4/A2/M3/M2/_0_  (.A1(\V1/V2/V4/A2/M3/s1 ),
    .A2(\V1/V2/V4/A2/c2 ),
    .ZN(\V1/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M3/M2/_1_  (.A(\V1/V2/V4/A2/M3/s1 ),
    .B(\V1/V2/V4/A2/c2 ),
    .Z(\V1/V2/V4/s2 [2]));
 OR2_X1 \V1/V2/V4/A2/M3/_0_  (.A1(\V1/V2/V4/A2/M3/c1 ),
    .A2(\V1/V2/V4/A2/M3/c2 ),
    .ZN(\V1/V2/V4/A2/c3 ));
 AND2_X1 \V1/V2/V4/A2/M4/M1/_0_  (.A1(\V1/V2/V4/s1 [3]),
    .A2(ground),
    .ZN(\V1/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M4/M1/_1_  (.A(\V1/V2/V4/s1 [3]),
    .B(ground),
    .Z(\V1/V2/V4/A2/M4/s1 ));
 AND2_X1 \V1/V2/V4/A2/M4/M2/_0_  (.A1(\V1/V2/V4/A2/M4/s1 ),
    .A2(\V1/V2/V4/A2/c3 ),
    .ZN(\V1/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M4/M2/_1_  (.A(\V1/V2/V4/A2/M4/s1 ),
    .B(\V1/V2/V4/A2/c3 ),
    .Z(\V1/V2/V4/s2 [3]));
 OR2_X1 \V1/V2/V4/A2/M4/_0_  (.A1(\V1/V2/V4/A2/M4/c1 ),
    .A2(\V1/V2/V4/A2/M4/c2 ),
    .ZN(\V1/V2/V4/c2 ));
 AND2_X1 \V1/V2/V4/A3/M1/M1/_0_  (.A1(\V1/V2/V4/v4 [0]),
    .A2(\V1/V2/V4/s2 [2]),
    .ZN(\V1/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M1/M1/_1_  (.A(\V1/V2/V4/v4 [0]),
    .B(\V1/V2/V4/s2 [2]),
    .Z(\V1/V2/V4/A3/M1/s1 ));
 AND2_X1 \V1/V2/V4/A3/M1/M2/_0_  (.A1(\V1/V2/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M1/M2/_1_  (.A(\V1/V2/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V2/v4 [4]));
 OR2_X1 \V1/V2/V4/A3/M1/_0_  (.A1(\V1/V2/V4/A3/M1/c1 ),
    .A2(\V1/V2/V4/A3/M1/c2 ),
    .ZN(\V1/V2/V4/A3/c1 ));
 AND2_X1 \V1/V2/V4/A3/M2/M1/_0_  (.A1(\V1/V2/V4/v4 [1]),
    .A2(\V1/V2/V4/s2 [3]),
    .ZN(\V1/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M2/M1/_1_  (.A(\V1/V2/V4/v4 [1]),
    .B(\V1/V2/V4/s2 [3]),
    .Z(\V1/V2/V4/A3/M2/s1 ));
 AND2_X1 \V1/V2/V4/A3/M2/M2/_0_  (.A1(\V1/V2/V4/A3/M2/s1 ),
    .A2(\V1/V2/V4/A3/c1 ),
    .ZN(\V1/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M2/M2/_1_  (.A(\V1/V2/V4/A3/M2/s1 ),
    .B(\V1/V2/V4/A3/c1 ),
    .Z(\V1/V2/v4 [5]));
 OR2_X1 \V1/V2/V4/A3/M2/_0_  (.A1(\V1/V2/V4/A3/M2/c1 ),
    .A2(\V1/V2/V4/A3/M2/c2 ),
    .ZN(\V1/V2/V4/A3/c2 ));
 AND2_X1 \V1/V2/V4/A3/M3/M1/_0_  (.A1(\V1/V2/V4/v4 [2]),
    .A2(\V1/V2/V4/c3 ),
    .ZN(\V1/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M3/M1/_1_  (.A(\V1/V2/V4/v4 [2]),
    .B(\V1/V2/V4/c3 ),
    .Z(\V1/V2/V4/A3/M3/s1 ));
 AND2_X1 \V1/V2/V4/A3/M3/M2/_0_  (.A1(\V1/V2/V4/A3/M3/s1 ),
    .A2(\V1/V2/V4/A3/c2 ),
    .ZN(\V1/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M3/M2/_1_  (.A(\V1/V2/V4/A3/M3/s1 ),
    .B(\V1/V2/V4/A3/c2 ),
    .Z(\V1/V2/v4 [6]));
 OR2_X1 \V1/V2/V4/A3/M3/_0_  (.A1(\V1/V2/V4/A3/M3/c1 ),
    .A2(\V1/V2/V4/A3/M3/c2 ),
    .ZN(\V1/V2/V4/A3/c3 ));
 AND2_X1 \V1/V2/V4/A3/M4/M1/_0_  (.A1(\V1/V2/V4/v4 [3]),
    .A2(ground),
    .ZN(\V1/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M4/M1/_1_  (.A(\V1/V2/V4/v4 [3]),
    .B(ground),
    .Z(\V1/V2/V4/A3/M4/s1 ));
 AND2_X1 \V1/V2/V4/A3/M4/M2/_0_  (.A1(\V1/V2/V4/A3/M4/s1 ),
    .A2(\V1/V2/V4/A3/c3 ),
    .ZN(\V1/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M4/M2/_1_  (.A(\V1/V2/V4/A3/M4/s1 ),
    .B(\V1/V2/V4/A3/c3 ),
    .Z(\V1/V2/v4 [7]));
 OR2_X1 \V1/V2/V4/A3/M4/_0_  (.A1(\V1/V2/V4/A3/M4/c1 ),
    .A2(\V1/V2/V4/A3/M4/c2 ),
    .ZN(\V1/V2/V4/overflow ));
 AND2_X1 \V1/V2/V4/V1/HA1/_0_  (.A1(\V1/V2/V4/V1/w2 ),
    .A2(\V1/V2/V4/V1/w1 ),
    .ZN(\V1/V2/V4/V1/w4 ));
 XOR2_X2 \V1/V2/V4/V1/HA1/_1_  (.A(\V1/V2/V4/V1/w2 ),
    .B(\V1/V2/V4/V1/w1 ),
    .Z(\V1/V2/v4 [1]));
 AND2_X1 \V1/V2/V4/V1/HA2/_0_  (.A1(\V1/V2/V4/V1/w4 ),
    .A2(\V1/V2/V4/V1/w3 ),
    .ZN(\V1/V2/V4/v1 [3]));
 XOR2_X2 \V1/V2/V4/V1/HA2/_1_  (.A(\V1/V2/V4/V1/w4 ),
    .B(\V1/V2/V4/V1/w3 ),
    .Z(\V1/V2/V4/v1 [2]));
 AND2_X1 \V1/V2/V4/V1/_0_  (.A1(A[12]),
    .A2(B[4]),
    .ZN(\V1/V2/v4 [0]));
 AND2_X1 \V1/V2/V4/V1/_1_  (.A1(A[12]),
    .A2(B[5]),
    .ZN(\V1/V2/V4/V1/w1 ));
 AND2_X1 \V1/V2/V4/V1/_2_  (.A1(B[4]),
    .A2(A[13]),
    .ZN(\V1/V2/V4/V1/w2 ));
 AND2_X1 \V1/V2/V4/V1/_3_  (.A1(B[5]),
    .A2(A[13]),
    .ZN(\V1/V2/V4/V1/w3 ));
 AND2_X1 \V1/V2/V4/V2/HA1/_0_  (.A1(\V1/V2/V4/V2/w2 ),
    .A2(\V1/V2/V4/V2/w1 ),
    .ZN(\V1/V2/V4/V2/w4 ));
 XOR2_X2 \V1/V2/V4/V2/HA1/_1_  (.A(\V1/V2/V4/V2/w2 ),
    .B(\V1/V2/V4/V2/w1 ),
    .Z(\V1/V2/V4/v2 [1]));
 AND2_X1 \V1/V2/V4/V2/HA2/_0_  (.A1(\V1/V2/V4/V2/w4 ),
    .A2(\V1/V2/V4/V2/w3 ),
    .ZN(\V1/V2/V4/v2 [3]));
 XOR2_X2 \V1/V2/V4/V2/HA2/_1_  (.A(\V1/V2/V4/V2/w4 ),
    .B(\V1/V2/V4/V2/w3 ),
    .Z(\V1/V2/V4/v2 [2]));
 AND2_X1 \V1/V2/V4/V2/_0_  (.A1(A[14]),
    .A2(B[4]),
    .ZN(\V1/V2/V4/v2 [0]));
 AND2_X1 \V1/V2/V4/V2/_1_  (.A1(A[14]),
    .A2(B[5]),
    .ZN(\V1/V2/V4/V2/w1 ));
 AND2_X1 \V1/V2/V4/V2/_2_  (.A1(B[4]),
    .A2(A[15]),
    .ZN(\V1/V2/V4/V2/w2 ));
 AND2_X1 \V1/V2/V4/V2/_3_  (.A1(B[5]),
    .A2(A[15]),
    .ZN(\V1/V2/V4/V2/w3 ));
 AND2_X1 \V1/V2/V4/V3/HA1/_0_  (.A1(\V1/V2/V4/V3/w2 ),
    .A2(\V1/V2/V4/V3/w1 ),
    .ZN(\V1/V2/V4/V3/w4 ));
 XOR2_X2 \V1/V2/V4/V3/HA1/_1_  (.A(\V1/V2/V4/V3/w2 ),
    .B(\V1/V2/V4/V3/w1 ),
    .Z(\V1/V2/V4/v3 [1]));
 AND2_X1 \V1/V2/V4/V3/HA2/_0_  (.A1(\V1/V2/V4/V3/w4 ),
    .A2(\V1/V2/V4/V3/w3 ),
    .ZN(\V1/V2/V4/v3 [3]));
 XOR2_X2 \V1/V2/V4/V3/HA2/_1_  (.A(\V1/V2/V4/V3/w4 ),
    .B(\V1/V2/V4/V3/w3 ),
    .Z(\V1/V2/V4/v3 [2]));
 AND2_X1 \V1/V2/V4/V3/_0_  (.A1(A[12]),
    .A2(B[6]),
    .ZN(\V1/V2/V4/v3 [0]));
 AND2_X1 \V1/V2/V4/V3/_1_  (.A1(A[12]),
    .A2(B[7]),
    .ZN(\V1/V2/V4/V3/w1 ));
 AND2_X1 \V1/V2/V4/V3/_2_  (.A1(B[6]),
    .A2(A[13]),
    .ZN(\V1/V2/V4/V3/w2 ));
 AND2_X1 \V1/V2/V4/V3/_3_  (.A1(B[7]),
    .A2(A[13]),
    .ZN(\V1/V2/V4/V3/w3 ));
 AND2_X1 \V1/V2/V4/V4/HA1/_0_  (.A1(\V1/V2/V4/V4/w2 ),
    .A2(\V1/V2/V4/V4/w1 ),
    .ZN(\V1/V2/V4/V4/w4 ));
 XOR2_X2 \V1/V2/V4/V4/HA1/_1_  (.A(\V1/V2/V4/V4/w2 ),
    .B(\V1/V2/V4/V4/w1 ),
    .Z(\V1/V2/V4/v4 [1]));
 AND2_X1 \V1/V2/V4/V4/HA2/_0_  (.A1(\V1/V2/V4/V4/w4 ),
    .A2(\V1/V2/V4/V4/w3 ),
    .ZN(\V1/V2/V4/v4 [3]));
 XOR2_X2 \V1/V2/V4/V4/HA2/_1_  (.A(\V1/V2/V4/V4/w4 ),
    .B(\V1/V2/V4/V4/w3 ),
    .Z(\V1/V2/V4/v4 [2]));
 AND2_X1 \V1/V2/V4/V4/_0_  (.A1(A[14]),
    .A2(B[6]),
    .ZN(\V1/V2/V4/v4 [0]));
 AND2_X1 \V1/V2/V4/V4/_1_  (.A1(A[14]),
    .A2(B[7]),
    .ZN(\V1/V2/V4/V4/w1 ));
 AND2_X1 \V1/V2/V4/V4/_2_  (.A1(B[6]),
    .A2(A[15]),
    .ZN(\V1/V2/V4/V4/w2 ));
 AND2_X1 \V1/V2/V4/V4/_3_  (.A1(B[7]),
    .A2(A[15]),
    .ZN(\V1/V2/V4/V4/w3 ));
 OR2_X1 \V1/V2/V4/_0_  (.A1(\V1/V2/V4/c1 ),
    .A2(\V1/V2/V4/c2 ),
    .ZN(\V1/V2/V4/c3 ));
 OR2_X1 \V1/V2/_0_  (.A1(\V1/V2/c1 ),
    .A2(\V1/V2/c2 ),
    .ZN(\V1/V2/c3 ));
 AND2_X1 \V1/V3/A1/A1/M1/M1/_0_  (.A1(\V1/V3/v2 [0]),
    .A2(\V1/V3/v3 [0]),
    .ZN(\V1/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M1/M1/_1_  (.A(\V1/V3/v2 [0]),
    .B(\V1/V3/v3 [0]),
    .Z(\V1/V3/A1/A1/M1/s1 ));
 AND2_X1 \V1/V3/A1/A1/M1/M2/_0_  (.A1(\V1/V3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M1/M2/_1_  (.A(\V1/V3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/s1 [0]));
 OR2_X1 \V1/V3/A1/A1/M1/_0_  (.A1(\V1/V3/A1/A1/M1/c1 ),
    .A2(\V1/V3/A1/A1/M1/c2 ),
    .ZN(\V1/V3/A1/A1/c1 ));
 AND2_X1 \V1/V3/A1/A1/M2/M1/_0_  (.A1(\V1/V3/v2 [1]),
    .A2(\V1/V3/v3 [1]),
    .ZN(\V1/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M2/M1/_1_  (.A(\V1/V3/v2 [1]),
    .B(\V1/V3/v3 [1]),
    .Z(\V1/V3/A1/A1/M2/s1 ));
 AND2_X1 \V1/V3/A1/A1/M2/M2/_0_  (.A1(\V1/V3/A1/A1/M2/s1 ),
    .A2(\V1/V3/A1/A1/c1 ),
    .ZN(\V1/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M2/M2/_1_  (.A(\V1/V3/A1/A1/M2/s1 ),
    .B(\V1/V3/A1/A1/c1 ),
    .Z(\V1/V3/s1 [1]));
 OR2_X1 \V1/V3/A1/A1/M2/_0_  (.A1(\V1/V3/A1/A1/M2/c1 ),
    .A2(\V1/V3/A1/A1/M2/c2 ),
    .ZN(\V1/V3/A1/A1/c2 ));
 AND2_X1 \V1/V3/A1/A1/M3/M1/_0_  (.A1(\V1/V3/v2 [2]),
    .A2(\V1/V3/v3 [2]),
    .ZN(\V1/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M3/M1/_1_  (.A(\V1/V3/v2 [2]),
    .B(\V1/V3/v3 [2]),
    .Z(\V1/V3/A1/A1/M3/s1 ));
 AND2_X1 \V1/V3/A1/A1/M3/M2/_0_  (.A1(\V1/V3/A1/A1/M3/s1 ),
    .A2(\V1/V3/A1/A1/c2 ),
    .ZN(\V1/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M3/M2/_1_  (.A(\V1/V3/A1/A1/M3/s1 ),
    .B(\V1/V3/A1/A1/c2 ),
    .Z(\V1/V3/s1 [2]));
 OR2_X1 \V1/V3/A1/A1/M3/_0_  (.A1(\V1/V3/A1/A1/M3/c1 ),
    .A2(\V1/V3/A1/A1/M3/c2 ),
    .ZN(\V1/V3/A1/A1/c3 ));
 AND2_X1 \V1/V3/A1/A1/M4/M1/_0_  (.A1(\V1/V3/v2 [3]),
    .A2(\V1/V3/v3 [3]),
    .ZN(\V1/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M4/M1/_1_  (.A(\V1/V3/v2 [3]),
    .B(\V1/V3/v3 [3]),
    .Z(\V1/V3/A1/A1/M4/s1 ));
 AND2_X1 \V1/V3/A1/A1/M4/M2/_0_  (.A1(\V1/V3/A1/A1/M4/s1 ),
    .A2(\V1/V3/A1/A1/c3 ),
    .ZN(\V1/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M4/M2/_1_  (.A(\V1/V3/A1/A1/M4/s1 ),
    .B(\V1/V3/A1/A1/c3 ),
    .Z(\V1/V3/s1 [3]));
 OR2_X1 \V1/V3/A1/A1/M4/_0_  (.A1(\V1/V3/A1/A1/M4/c1 ),
    .A2(\V1/V3/A1/A1/M4/c2 ),
    .ZN(\V1/V3/A1/c1 ));
 AND2_X1 \V1/V3/A1/A2/M1/M1/_0_  (.A1(\V1/V3/v2 [4]),
    .A2(\V1/V3/v3 [4]),
    .ZN(\V1/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M1/M1/_1_  (.A(\V1/V3/v2 [4]),
    .B(\V1/V3/v3 [4]),
    .Z(\V1/V3/A1/A2/M1/s1 ));
 AND2_X1 \V1/V3/A1/A2/M1/M2/_0_  (.A1(\V1/V3/A1/A2/M1/s1 ),
    .A2(\V1/V3/A1/c1 ),
    .ZN(\V1/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M1/M2/_1_  (.A(\V1/V3/A1/A2/M1/s1 ),
    .B(\V1/V3/A1/c1 ),
    .Z(\V1/V3/s1 [4]));
 OR2_X1 \V1/V3/A1/A2/M1/_0_  (.A1(\V1/V3/A1/A2/M1/c1 ),
    .A2(\V1/V3/A1/A2/M1/c2 ),
    .ZN(\V1/V3/A1/A2/c1 ));
 AND2_X1 \V1/V3/A1/A2/M2/M1/_0_  (.A1(\V1/V3/v2 [5]),
    .A2(\V1/V3/v3 [5]),
    .ZN(\V1/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M2/M1/_1_  (.A(\V1/V3/v2 [5]),
    .B(\V1/V3/v3 [5]),
    .Z(\V1/V3/A1/A2/M2/s1 ));
 AND2_X1 \V1/V3/A1/A2/M2/M2/_0_  (.A1(\V1/V3/A1/A2/M2/s1 ),
    .A2(\V1/V3/A1/A2/c1 ),
    .ZN(\V1/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M2/M2/_1_  (.A(\V1/V3/A1/A2/M2/s1 ),
    .B(\V1/V3/A1/A2/c1 ),
    .Z(\V1/V3/s1 [5]));
 OR2_X1 \V1/V3/A1/A2/M2/_0_  (.A1(\V1/V3/A1/A2/M2/c1 ),
    .A2(\V1/V3/A1/A2/M2/c2 ),
    .ZN(\V1/V3/A1/A2/c2 ));
 AND2_X1 \V1/V3/A1/A2/M3/M1/_0_  (.A1(\V1/V3/v2 [6]),
    .A2(\V1/V3/v3 [6]),
    .ZN(\V1/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M3/M1/_1_  (.A(\V1/V3/v2 [6]),
    .B(\V1/V3/v3 [6]),
    .Z(\V1/V3/A1/A2/M3/s1 ));
 AND2_X1 \V1/V3/A1/A2/M3/M2/_0_  (.A1(\V1/V3/A1/A2/M3/s1 ),
    .A2(\V1/V3/A1/A2/c2 ),
    .ZN(\V1/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M3/M2/_1_  (.A(\V1/V3/A1/A2/M3/s1 ),
    .B(\V1/V3/A1/A2/c2 ),
    .Z(\V1/V3/s1 [6]));
 OR2_X1 \V1/V3/A1/A2/M3/_0_  (.A1(\V1/V3/A1/A2/M3/c1 ),
    .A2(\V1/V3/A1/A2/M3/c2 ),
    .ZN(\V1/V3/A1/A2/c3 ));
 AND2_X1 \V1/V3/A1/A2/M4/M1/_0_  (.A1(\V1/V3/v2 [7]),
    .A2(\V1/V3/v3 [7]),
    .ZN(\V1/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M4/M1/_1_  (.A(\V1/V3/v2 [7]),
    .B(\V1/V3/v3 [7]),
    .Z(\V1/V3/A1/A2/M4/s1 ));
 AND2_X1 \V1/V3/A1/A2/M4/M2/_0_  (.A1(\V1/V3/A1/A2/M4/s1 ),
    .A2(\V1/V3/A1/A2/c3 ),
    .ZN(\V1/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M4/M2/_1_  (.A(\V1/V3/A1/A2/M4/s1 ),
    .B(\V1/V3/A1/A2/c3 ),
    .Z(\V1/V3/s1 [7]));
 OR2_X1 \V1/V3/A1/A2/M4/_0_  (.A1(\V1/V3/A1/A2/M4/c1 ),
    .A2(\V1/V3/A1/A2/M4/c2 ),
    .ZN(\V1/V3/c1 ));
 AND2_X1 \V1/V3/A2/A1/M1/M1/_0_  (.A1(\V1/V3/s1 [0]),
    .A2(\V1/V3/v1 [4]),
    .ZN(\V1/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M1/M1/_1_  (.A(\V1/V3/s1 [0]),
    .B(\V1/V3/v1 [4]),
    .Z(\V1/V3/A2/A1/M1/s1 ));
 AND2_X1 \V1/V3/A2/A1/M1/M2/_0_  (.A1(\V1/V3/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M1/M2/_1_  (.A(\V1/V3/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v3 [4]));
 OR2_X1 \V1/V3/A2/A1/M1/_0_  (.A1(\V1/V3/A2/A1/M1/c1 ),
    .A2(\V1/V3/A2/A1/M1/c2 ),
    .ZN(\V1/V3/A2/A1/c1 ));
 AND2_X1 \V1/V3/A2/A1/M2/M1/_0_  (.A1(\V1/V3/s1 [1]),
    .A2(\V1/V3/v1 [5]),
    .ZN(\V1/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M2/M1/_1_  (.A(\V1/V3/s1 [1]),
    .B(\V1/V3/v1 [5]),
    .Z(\V1/V3/A2/A1/M2/s1 ));
 AND2_X1 \V1/V3/A2/A1/M2/M2/_0_  (.A1(\V1/V3/A2/A1/M2/s1 ),
    .A2(\V1/V3/A2/A1/c1 ),
    .ZN(\V1/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M2/M2/_1_  (.A(\V1/V3/A2/A1/M2/s1 ),
    .B(\V1/V3/A2/A1/c1 ),
    .Z(\V1/v3 [5]));
 OR2_X1 \V1/V3/A2/A1/M2/_0_  (.A1(\V1/V3/A2/A1/M2/c1 ),
    .A2(\V1/V3/A2/A1/M2/c2 ),
    .ZN(\V1/V3/A2/A1/c2 ));
 AND2_X1 \V1/V3/A2/A1/M3/M1/_0_  (.A1(\V1/V3/s1 [2]),
    .A2(\V1/V3/v1 [6]),
    .ZN(\V1/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M3/M1/_1_  (.A(\V1/V3/s1 [2]),
    .B(\V1/V3/v1 [6]),
    .Z(\V1/V3/A2/A1/M3/s1 ));
 AND2_X1 \V1/V3/A2/A1/M3/M2/_0_  (.A1(\V1/V3/A2/A1/M3/s1 ),
    .A2(\V1/V3/A2/A1/c2 ),
    .ZN(\V1/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M3/M2/_1_  (.A(\V1/V3/A2/A1/M3/s1 ),
    .B(\V1/V3/A2/A1/c2 ),
    .Z(\V1/v3 [6]));
 OR2_X1 \V1/V3/A2/A1/M3/_0_  (.A1(\V1/V3/A2/A1/M3/c1 ),
    .A2(\V1/V3/A2/A1/M3/c2 ),
    .ZN(\V1/V3/A2/A1/c3 ));
 AND2_X1 \V1/V3/A2/A1/M4/M1/_0_  (.A1(\V1/V3/s1 [3]),
    .A2(\V1/V3/v1 [7]),
    .ZN(\V1/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M4/M1/_1_  (.A(\V1/V3/s1 [3]),
    .B(\V1/V3/v1 [7]),
    .Z(\V1/V3/A2/A1/M4/s1 ));
 AND2_X1 \V1/V3/A2/A1/M4/M2/_0_  (.A1(\V1/V3/A2/A1/M4/s1 ),
    .A2(\V1/V3/A2/A1/c3 ),
    .ZN(\V1/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M4/M2/_1_  (.A(\V1/V3/A2/A1/M4/s1 ),
    .B(\V1/V3/A2/A1/c3 ),
    .Z(\V1/v3 [7]));
 OR2_X1 \V1/V3/A2/A1/M4/_0_  (.A1(\V1/V3/A2/A1/M4/c1 ),
    .A2(\V1/V3/A2/A1/M4/c2 ),
    .ZN(\V1/V3/A2/c1 ));
 AND2_X1 \V1/V3/A2/A2/M1/M1/_0_  (.A1(\V1/V3/s1 [4]),
    .A2(ground),
    .ZN(\V1/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M1/M1/_1_  (.A(\V1/V3/s1 [4]),
    .B(ground),
    .Z(\V1/V3/A2/A2/M1/s1 ));
 AND2_X1 \V1/V3/A2/A2/M1/M2/_0_  (.A1(\V1/V3/A2/A2/M1/s1 ),
    .A2(\V1/V3/A2/c1 ),
    .ZN(\V1/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M1/M2/_1_  (.A(\V1/V3/A2/A2/M1/s1 ),
    .B(\V1/V3/A2/c1 ),
    .Z(\V1/V3/s2 [4]));
 OR2_X1 \V1/V3/A2/A2/M1/_0_  (.A1(\V1/V3/A2/A2/M1/c1 ),
    .A2(\V1/V3/A2/A2/M1/c2 ),
    .ZN(\V1/V3/A2/A2/c1 ));
 AND2_X1 \V1/V3/A2/A2/M2/M1/_0_  (.A1(\V1/V3/s1 [5]),
    .A2(ground),
    .ZN(\V1/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M2/M1/_1_  (.A(\V1/V3/s1 [5]),
    .B(ground),
    .Z(\V1/V3/A2/A2/M2/s1 ));
 AND2_X1 \V1/V3/A2/A2/M2/M2/_0_  (.A1(\V1/V3/A2/A2/M2/s1 ),
    .A2(\V1/V3/A2/A2/c1 ),
    .ZN(\V1/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M2/M2/_1_  (.A(\V1/V3/A2/A2/M2/s1 ),
    .B(\V1/V3/A2/A2/c1 ),
    .Z(\V1/V3/s2 [5]));
 OR2_X1 \V1/V3/A2/A2/M2/_0_  (.A1(\V1/V3/A2/A2/M2/c1 ),
    .A2(\V1/V3/A2/A2/M2/c2 ),
    .ZN(\V1/V3/A2/A2/c2 ));
 AND2_X1 \V1/V3/A2/A2/M3/M1/_0_  (.A1(\V1/V3/s1 [6]),
    .A2(ground),
    .ZN(\V1/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M3/M1/_1_  (.A(\V1/V3/s1 [6]),
    .B(ground),
    .Z(\V1/V3/A2/A2/M3/s1 ));
 AND2_X1 \V1/V3/A2/A2/M3/M2/_0_  (.A1(\V1/V3/A2/A2/M3/s1 ),
    .A2(\V1/V3/A2/A2/c2 ),
    .ZN(\V1/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M3/M2/_1_  (.A(\V1/V3/A2/A2/M3/s1 ),
    .B(\V1/V3/A2/A2/c2 ),
    .Z(\V1/V3/s2 [6]));
 OR2_X1 \V1/V3/A2/A2/M3/_0_  (.A1(\V1/V3/A2/A2/M3/c1 ),
    .A2(\V1/V3/A2/A2/M3/c2 ),
    .ZN(\V1/V3/A2/A2/c3 ));
 AND2_X1 \V1/V3/A2/A2/M4/M1/_0_  (.A1(\V1/V3/s1 [7]),
    .A2(ground),
    .ZN(\V1/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M4/M1/_1_  (.A(\V1/V3/s1 [7]),
    .B(ground),
    .Z(\V1/V3/A2/A2/M4/s1 ));
 AND2_X1 \V1/V3/A2/A2/M4/M2/_0_  (.A1(\V1/V3/A2/A2/M4/s1 ),
    .A2(\V1/V3/A2/A2/c3 ),
    .ZN(\V1/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M4/M2/_1_  (.A(\V1/V3/A2/A2/M4/s1 ),
    .B(\V1/V3/A2/A2/c3 ),
    .Z(\V1/V3/s2 [7]));
 OR2_X1 \V1/V3/A2/A2/M4/_0_  (.A1(\V1/V3/A2/A2/M4/c1 ),
    .A2(\V1/V3/A2/A2/M4/c2 ),
    .ZN(\V1/V3/c2 ));
 AND2_X1 \V1/V3/A3/A1/M1/M1/_0_  (.A1(\V1/V3/v4 [0]),
    .A2(\V1/V3/s2 [4]),
    .ZN(\V1/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M1/M1/_1_  (.A(\V1/V3/v4 [0]),
    .B(\V1/V3/s2 [4]),
    .Z(\V1/V3/A3/A1/M1/s1 ));
 AND2_X1 \V1/V3/A3/A1/M1/M2/_0_  (.A1(\V1/V3/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M1/M2/_1_  (.A(\V1/V3/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v3 [8]));
 OR2_X1 \V1/V3/A3/A1/M1/_0_  (.A1(\V1/V3/A3/A1/M1/c1 ),
    .A2(\V1/V3/A3/A1/M1/c2 ),
    .ZN(\V1/V3/A3/A1/c1 ));
 AND2_X1 \V1/V3/A3/A1/M2/M1/_0_  (.A1(\V1/V3/v4 [1]),
    .A2(\V1/V3/s2 [5]),
    .ZN(\V1/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M2/M1/_1_  (.A(\V1/V3/v4 [1]),
    .B(\V1/V3/s2 [5]),
    .Z(\V1/V3/A3/A1/M2/s1 ));
 AND2_X1 \V1/V3/A3/A1/M2/M2/_0_  (.A1(\V1/V3/A3/A1/M2/s1 ),
    .A2(\V1/V3/A3/A1/c1 ),
    .ZN(\V1/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M2/M2/_1_  (.A(\V1/V3/A3/A1/M2/s1 ),
    .B(\V1/V3/A3/A1/c1 ),
    .Z(\V1/v3 [9]));
 OR2_X1 \V1/V3/A3/A1/M2/_0_  (.A1(\V1/V3/A3/A1/M2/c1 ),
    .A2(\V1/V3/A3/A1/M2/c2 ),
    .ZN(\V1/V3/A3/A1/c2 ));
 AND2_X1 \V1/V3/A3/A1/M3/M1/_0_  (.A1(\V1/V3/v4 [2]),
    .A2(\V1/V3/s2 [6]),
    .ZN(\V1/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M3/M1/_1_  (.A(\V1/V3/v4 [2]),
    .B(\V1/V3/s2 [6]),
    .Z(\V1/V3/A3/A1/M3/s1 ));
 AND2_X1 \V1/V3/A3/A1/M3/M2/_0_  (.A1(\V1/V3/A3/A1/M3/s1 ),
    .A2(\V1/V3/A3/A1/c2 ),
    .ZN(\V1/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M3/M2/_1_  (.A(\V1/V3/A3/A1/M3/s1 ),
    .B(\V1/V3/A3/A1/c2 ),
    .Z(\V1/v3 [10]));
 OR2_X1 \V1/V3/A3/A1/M3/_0_  (.A1(\V1/V3/A3/A1/M3/c1 ),
    .A2(\V1/V3/A3/A1/M3/c2 ),
    .ZN(\V1/V3/A3/A1/c3 ));
 AND2_X1 \V1/V3/A3/A1/M4/M1/_0_  (.A1(\V1/V3/v4 [3]),
    .A2(\V1/V3/s2 [7]),
    .ZN(\V1/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M4/M1/_1_  (.A(\V1/V3/v4 [3]),
    .B(\V1/V3/s2 [7]),
    .Z(\V1/V3/A3/A1/M4/s1 ));
 AND2_X1 \V1/V3/A3/A1/M4/M2/_0_  (.A1(\V1/V3/A3/A1/M4/s1 ),
    .A2(\V1/V3/A3/A1/c3 ),
    .ZN(\V1/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M4/M2/_1_  (.A(\V1/V3/A3/A1/M4/s1 ),
    .B(\V1/V3/A3/A1/c3 ),
    .Z(\V1/v3 [11]));
 OR2_X1 \V1/V3/A3/A1/M4/_0_  (.A1(\V1/V3/A3/A1/M4/c1 ),
    .A2(\V1/V3/A3/A1/M4/c2 ),
    .ZN(\V1/V3/A3/c1 ));
 AND2_X1 \V1/V3/A3/A2/M1/M1/_0_  (.A1(\V1/V3/v4 [4]),
    .A2(\V1/V3/c3 ),
    .ZN(\V1/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M1/M1/_1_  (.A(\V1/V3/v4 [4]),
    .B(\V1/V3/c3 ),
    .Z(\V1/V3/A3/A2/M1/s1 ));
 AND2_X1 \V1/V3/A3/A2/M1/M2/_0_  (.A1(\V1/V3/A3/A2/M1/s1 ),
    .A2(\V1/V3/A3/c1 ),
    .ZN(\V1/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M1/M2/_1_  (.A(\V1/V3/A3/A2/M1/s1 ),
    .B(\V1/V3/A3/c1 ),
    .Z(\V1/v3 [12]));
 OR2_X1 \V1/V3/A3/A2/M1/_0_  (.A1(\V1/V3/A3/A2/M1/c1 ),
    .A2(\V1/V3/A3/A2/M1/c2 ),
    .ZN(\V1/V3/A3/A2/c1 ));
 AND2_X1 \V1/V3/A3/A2/M2/M1/_0_  (.A1(\V1/V3/v4 [5]),
    .A2(ground),
    .ZN(\V1/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M2/M1/_1_  (.A(\V1/V3/v4 [5]),
    .B(ground),
    .Z(\V1/V3/A3/A2/M2/s1 ));
 AND2_X1 \V1/V3/A3/A2/M2/M2/_0_  (.A1(\V1/V3/A3/A2/M2/s1 ),
    .A2(\V1/V3/A3/A2/c1 ),
    .ZN(\V1/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M2/M2/_1_  (.A(\V1/V3/A3/A2/M2/s1 ),
    .B(\V1/V3/A3/A2/c1 ),
    .Z(\V1/v3 [13]));
 OR2_X1 \V1/V3/A3/A2/M2/_0_  (.A1(\V1/V3/A3/A2/M2/c1 ),
    .A2(\V1/V3/A3/A2/M2/c2 ),
    .ZN(\V1/V3/A3/A2/c2 ));
 AND2_X1 \V1/V3/A3/A2/M3/M1/_0_  (.A1(\V1/V3/v4 [6]),
    .A2(ground),
    .ZN(\V1/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M3/M1/_1_  (.A(\V1/V3/v4 [6]),
    .B(ground),
    .Z(\V1/V3/A3/A2/M3/s1 ));
 AND2_X1 \V1/V3/A3/A2/M3/M2/_0_  (.A1(\V1/V3/A3/A2/M3/s1 ),
    .A2(\V1/V3/A3/A2/c2 ),
    .ZN(\V1/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M3/M2/_1_  (.A(\V1/V3/A3/A2/M3/s1 ),
    .B(\V1/V3/A3/A2/c2 ),
    .Z(\V1/v3 [14]));
 OR2_X1 \V1/V3/A3/A2/M3/_0_  (.A1(\V1/V3/A3/A2/M3/c1 ),
    .A2(\V1/V3/A3/A2/M3/c2 ),
    .ZN(\V1/V3/A3/A2/c3 ));
 AND2_X1 \V1/V3/A3/A2/M4/M1/_0_  (.A1(\V1/V3/v4 [7]),
    .A2(ground),
    .ZN(\V1/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M4/M1/_1_  (.A(\V1/V3/v4 [7]),
    .B(ground),
    .Z(\V1/V3/A3/A2/M4/s1 ));
 AND2_X1 \V1/V3/A3/A2/M4/M2/_0_  (.A1(\V1/V3/A3/A2/M4/s1 ),
    .A2(\V1/V3/A3/A2/c3 ),
    .ZN(\V1/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M4/M2/_1_  (.A(\V1/V3/A3/A2/M4/s1 ),
    .B(\V1/V3/A3/A2/c3 ),
    .Z(\V1/v3 [15]));
 OR2_X1 \V1/V3/A3/A2/M4/_0_  (.A1(\V1/V3/A3/A2/M4/c1 ),
    .A2(\V1/V3/A3/A2/M4/c2 ),
    .ZN(\V1/V3/overflow ));
 AND2_X1 \V1/V3/V1/A1/M1/M1/_0_  (.A1(\V1/V3/V1/v2 [0]),
    .A2(\V1/V3/V1/v3 [0]),
    .ZN(\V1/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M1/M1/_1_  (.A(\V1/V3/V1/v2 [0]),
    .B(\V1/V3/V1/v3 [0]),
    .Z(\V1/V3/V1/A1/M1/s1 ));
 AND2_X1 \V1/V3/V1/A1/M1/M2/_0_  (.A1(\V1/V3/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M1/M2/_1_  (.A(\V1/V3/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/V1/s1 [0]));
 OR2_X1 \V1/V3/V1/A1/M1/_0_  (.A1(\V1/V3/V1/A1/M1/c1 ),
    .A2(\V1/V3/V1/A1/M1/c2 ),
    .ZN(\V1/V3/V1/A1/c1 ));
 AND2_X1 \V1/V3/V1/A1/M2/M1/_0_  (.A1(\V1/V3/V1/v2 [1]),
    .A2(\V1/V3/V1/v3 [1]),
    .ZN(\V1/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M2/M1/_1_  (.A(\V1/V3/V1/v2 [1]),
    .B(\V1/V3/V1/v3 [1]),
    .Z(\V1/V3/V1/A1/M2/s1 ));
 AND2_X1 \V1/V3/V1/A1/M2/M2/_0_  (.A1(\V1/V3/V1/A1/M2/s1 ),
    .A2(\V1/V3/V1/A1/c1 ),
    .ZN(\V1/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M2/M2/_1_  (.A(\V1/V3/V1/A1/M2/s1 ),
    .B(\V1/V3/V1/A1/c1 ),
    .Z(\V1/V3/V1/s1 [1]));
 OR2_X1 \V1/V3/V1/A1/M2/_0_  (.A1(\V1/V3/V1/A1/M2/c1 ),
    .A2(\V1/V3/V1/A1/M2/c2 ),
    .ZN(\V1/V3/V1/A1/c2 ));
 AND2_X1 \V1/V3/V1/A1/M3/M1/_0_  (.A1(\V1/V3/V1/v2 [2]),
    .A2(\V1/V3/V1/v3 [2]),
    .ZN(\V1/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M3/M1/_1_  (.A(\V1/V3/V1/v2 [2]),
    .B(\V1/V3/V1/v3 [2]),
    .Z(\V1/V3/V1/A1/M3/s1 ));
 AND2_X1 \V1/V3/V1/A1/M3/M2/_0_  (.A1(\V1/V3/V1/A1/M3/s1 ),
    .A2(\V1/V3/V1/A1/c2 ),
    .ZN(\V1/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M3/M2/_1_  (.A(\V1/V3/V1/A1/M3/s1 ),
    .B(\V1/V3/V1/A1/c2 ),
    .Z(\V1/V3/V1/s1 [2]));
 OR2_X1 \V1/V3/V1/A1/M3/_0_  (.A1(\V1/V3/V1/A1/M3/c1 ),
    .A2(\V1/V3/V1/A1/M3/c2 ),
    .ZN(\V1/V3/V1/A1/c3 ));
 AND2_X1 \V1/V3/V1/A1/M4/M1/_0_  (.A1(\V1/V3/V1/v2 [3]),
    .A2(\V1/V3/V1/v3 [3]),
    .ZN(\V1/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M4/M1/_1_  (.A(\V1/V3/V1/v2 [3]),
    .B(\V1/V3/V1/v3 [3]),
    .Z(\V1/V3/V1/A1/M4/s1 ));
 AND2_X1 \V1/V3/V1/A1/M4/M2/_0_  (.A1(\V1/V3/V1/A1/M4/s1 ),
    .A2(\V1/V3/V1/A1/c3 ),
    .ZN(\V1/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M4/M2/_1_  (.A(\V1/V3/V1/A1/M4/s1 ),
    .B(\V1/V3/V1/A1/c3 ),
    .Z(\V1/V3/V1/s1 [3]));
 OR2_X1 \V1/V3/V1/A1/M4/_0_  (.A1(\V1/V3/V1/A1/M4/c1 ),
    .A2(\V1/V3/V1/A1/M4/c2 ),
    .ZN(\V1/V3/V1/c1 ));
 AND2_X1 \V1/V3/V1/A2/M1/M1/_0_  (.A1(\V1/V3/V1/s1 [0]),
    .A2(\V1/V3/V1/v1 [2]),
    .ZN(\V1/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M1/M1/_1_  (.A(\V1/V3/V1/s1 [0]),
    .B(\V1/V3/V1/v1 [2]),
    .Z(\V1/V3/V1/A2/M1/s1 ));
 AND2_X1 \V1/V3/V1/A2/M1/M2/_0_  (.A1(\V1/V3/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M1/M2/_1_  (.A(\V1/V3/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/v3 [2]));
 OR2_X1 \V1/V3/V1/A2/M1/_0_  (.A1(\V1/V3/V1/A2/M1/c1 ),
    .A2(\V1/V3/V1/A2/M1/c2 ),
    .ZN(\V1/V3/V1/A2/c1 ));
 AND2_X1 \V1/V3/V1/A2/M2/M1/_0_  (.A1(\V1/V3/V1/s1 [1]),
    .A2(\V1/V3/V1/v1 [3]),
    .ZN(\V1/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M2/M1/_1_  (.A(\V1/V3/V1/s1 [1]),
    .B(\V1/V3/V1/v1 [3]),
    .Z(\V1/V3/V1/A2/M2/s1 ));
 AND2_X1 \V1/V3/V1/A2/M2/M2/_0_  (.A1(\V1/V3/V1/A2/M2/s1 ),
    .A2(\V1/V3/V1/A2/c1 ),
    .ZN(\V1/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M2/M2/_1_  (.A(\V1/V3/V1/A2/M2/s1 ),
    .B(\V1/V3/V1/A2/c1 ),
    .Z(\V1/v3 [3]));
 OR2_X1 \V1/V3/V1/A2/M2/_0_  (.A1(\V1/V3/V1/A2/M2/c1 ),
    .A2(\V1/V3/V1/A2/M2/c2 ),
    .ZN(\V1/V3/V1/A2/c2 ));
 AND2_X1 \V1/V3/V1/A2/M3/M1/_0_  (.A1(\V1/V3/V1/s1 [2]),
    .A2(ground),
    .ZN(\V1/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M3/M1/_1_  (.A(\V1/V3/V1/s1 [2]),
    .B(ground),
    .Z(\V1/V3/V1/A2/M3/s1 ));
 AND2_X1 \V1/V3/V1/A2/M3/M2/_0_  (.A1(\V1/V3/V1/A2/M3/s1 ),
    .A2(\V1/V3/V1/A2/c2 ),
    .ZN(\V1/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M3/M2/_1_  (.A(\V1/V3/V1/A2/M3/s1 ),
    .B(\V1/V3/V1/A2/c2 ),
    .Z(\V1/V3/V1/s2 [2]));
 OR2_X1 \V1/V3/V1/A2/M3/_0_  (.A1(\V1/V3/V1/A2/M3/c1 ),
    .A2(\V1/V3/V1/A2/M3/c2 ),
    .ZN(\V1/V3/V1/A2/c3 ));
 AND2_X1 \V1/V3/V1/A2/M4/M1/_0_  (.A1(\V1/V3/V1/s1 [3]),
    .A2(ground),
    .ZN(\V1/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M4/M1/_1_  (.A(\V1/V3/V1/s1 [3]),
    .B(ground),
    .Z(\V1/V3/V1/A2/M4/s1 ));
 AND2_X1 \V1/V3/V1/A2/M4/M2/_0_  (.A1(\V1/V3/V1/A2/M4/s1 ),
    .A2(\V1/V3/V1/A2/c3 ),
    .ZN(\V1/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M4/M2/_1_  (.A(\V1/V3/V1/A2/M4/s1 ),
    .B(\V1/V3/V1/A2/c3 ),
    .Z(\V1/V3/V1/s2 [3]));
 OR2_X1 \V1/V3/V1/A2/M4/_0_  (.A1(\V1/V3/V1/A2/M4/c1 ),
    .A2(\V1/V3/V1/A2/M4/c2 ),
    .ZN(\V1/V3/V1/c2 ));
 AND2_X1 \V1/V3/V1/A3/M1/M1/_0_  (.A1(\V1/V3/V1/v4 [0]),
    .A2(\V1/V3/V1/s2 [2]),
    .ZN(\V1/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M1/M1/_1_  (.A(\V1/V3/V1/v4 [0]),
    .B(\V1/V3/V1/s2 [2]),
    .Z(\V1/V3/V1/A3/M1/s1 ));
 AND2_X1 \V1/V3/V1/A3/M1/M2/_0_  (.A1(\V1/V3/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M1/M2/_1_  (.A(\V1/V3/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v1 [4]));
 OR2_X1 \V1/V3/V1/A3/M1/_0_  (.A1(\V1/V3/V1/A3/M1/c1 ),
    .A2(\V1/V3/V1/A3/M1/c2 ),
    .ZN(\V1/V3/V1/A3/c1 ));
 AND2_X1 \V1/V3/V1/A3/M2/M1/_0_  (.A1(\V1/V3/V1/v4 [1]),
    .A2(\V1/V3/V1/s2 [3]),
    .ZN(\V1/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M2/M1/_1_  (.A(\V1/V3/V1/v4 [1]),
    .B(\V1/V3/V1/s2 [3]),
    .Z(\V1/V3/V1/A3/M2/s1 ));
 AND2_X1 \V1/V3/V1/A3/M2/M2/_0_  (.A1(\V1/V3/V1/A3/M2/s1 ),
    .A2(\V1/V3/V1/A3/c1 ),
    .ZN(\V1/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M2/M2/_1_  (.A(\V1/V3/V1/A3/M2/s1 ),
    .B(\V1/V3/V1/A3/c1 ),
    .Z(\V1/V3/v1 [5]));
 OR2_X1 \V1/V3/V1/A3/M2/_0_  (.A1(\V1/V3/V1/A3/M2/c1 ),
    .A2(\V1/V3/V1/A3/M2/c2 ),
    .ZN(\V1/V3/V1/A3/c2 ));
 AND2_X1 \V1/V3/V1/A3/M3/M1/_0_  (.A1(\V1/V3/V1/v4 [2]),
    .A2(\V1/V3/V1/c3 ),
    .ZN(\V1/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M3/M1/_1_  (.A(\V1/V3/V1/v4 [2]),
    .B(\V1/V3/V1/c3 ),
    .Z(\V1/V3/V1/A3/M3/s1 ));
 AND2_X1 \V1/V3/V1/A3/M3/M2/_0_  (.A1(\V1/V3/V1/A3/M3/s1 ),
    .A2(\V1/V3/V1/A3/c2 ),
    .ZN(\V1/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M3/M2/_1_  (.A(\V1/V3/V1/A3/M3/s1 ),
    .B(\V1/V3/V1/A3/c2 ),
    .Z(\V1/V3/v1 [6]));
 OR2_X1 \V1/V3/V1/A3/M3/_0_  (.A1(\V1/V3/V1/A3/M3/c1 ),
    .A2(\V1/V3/V1/A3/M3/c2 ),
    .ZN(\V1/V3/V1/A3/c3 ));
 AND2_X1 \V1/V3/V1/A3/M4/M1/_0_  (.A1(\V1/V3/V1/v4 [3]),
    .A2(ground),
    .ZN(\V1/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M4/M1/_1_  (.A(\V1/V3/V1/v4 [3]),
    .B(ground),
    .Z(\V1/V3/V1/A3/M4/s1 ));
 AND2_X1 \V1/V3/V1/A3/M4/M2/_0_  (.A1(\V1/V3/V1/A3/M4/s1 ),
    .A2(\V1/V3/V1/A3/c3 ),
    .ZN(\V1/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M4/M2/_1_  (.A(\V1/V3/V1/A3/M4/s1 ),
    .B(\V1/V3/V1/A3/c3 ),
    .Z(\V1/V3/v1 [7]));
 OR2_X1 \V1/V3/V1/A3/M4/_0_  (.A1(\V1/V3/V1/A3/M4/c1 ),
    .A2(\V1/V3/V1/A3/M4/c2 ),
    .ZN(\V1/V3/V1/overflow ));
 AND2_X1 \V1/V3/V1/V1/HA1/_0_  (.A1(\V1/V3/V1/V1/w2 ),
    .A2(\V1/V3/V1/V1/w1 ),
    .ZN(\V1/V3/V1/V1/w4 ));
 XOR2_X2 \V1/V3/V1/V1/HA1/_1_  (.A(\V1/V3/V1/V1/w2 ),
    .B(\V1/V3/V1/V1/w1 ),
    .Z(\V1/v3 [1]));
 AND2_X1 \V1/V3/V1/V1/HA2/_0_  (.A1(\V1/V3/V1/V1/w4 ),
    .A2(\V1/V3/V1/V1/w3 ),
    .ZN(\V1/V3/V1/v1 [3]));
 XOR2_X2 \V1/V3/V1/V1/HA2/_1_  (.A(\V1/V3/V1/V1/w4 ),
    .B(\V1/V3/V1/V1/w3 ),
    .Z(\V1/V3/V1/v1 [2]));
 AND2_X1 \V1/V3/V1/V1/_0_  (.A1(A[0]),
    .A2(B[8]),
    .ZN(\V1/v3 [0]));
 AND2_X1 \V1/V3/V1/V1/_1_  (.A1(A[0]),
    .A2(B[9]),
    .ZN(\V1/V3/V1/V1/w1 ));
 AND2_X1 \V1/V3/V1/V1/_2_  (.A1(B[8]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V1/w2 ));
 AND2_X1 \V1/V3/V1/V1/_3_  (.A1(B[9]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V1/w3 ));
 AND2_X1 \V1/V3/V1/V2/HA1/_0_  (.A1(\V1/V3/V1/V2/w2 ),
    .A2(\V1/V3/V1/V2/w1 ),
    .ZN(\V1/V3/V1/V2/w4 ));
 XOR2_X2 \V1/V3/V1/V2/HA1/_1_  (.A(\V1/V3/V1/V2/w2 ),
    .B(\V1/V3/V1/V2/w1 ),
    .Z(\V1/V3/V1/v2 [1]));
 AND2_X1 \V1/V3/V1/V2/HA2/_0_  (.A1(\V1/V3/V1/V2/w4 ),
    .A2(\V1/V3/V1/V2/w3 ),
    .ZN(\V1/V3/V1/v2 [3]));
 XOR2_X2 \V1/V3/V1/V2/HA2/_1_  (.A(\V1/V3/V1/V2/w4 ),
    .B(\V1/V3/V1/V2/w3 ),
    .Z(\V1/V3/V1/v2 [2]));
 AND2_X1 \V1/V3/V1/V2/_0_  (.A1(A[2]),
    .A2(B[8]),
    .ZN(\V1/V3/V1/v2 [0]));
 AND2_X1 \V1/V3/V1/V2/_1_  (.A1(A[2]),
    .A2(B[9]),
    .ZN(\V1/V3/V1/V2/w1 ));
 AND2_X1 \V1/V3/V1/V2/_2_  (.A1(B[8]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V2/w2 ));
 AND2_X1 \V1/V3/V1/V2/_3_  (.A1(B[9]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V2/w3 ));
 AND2_X1 \V1/V3/V1/V3/HA1/_0_  (.A1(\V1/V3/V1/V3/w2 ),
    .A2(\V1/V3/V1/V3/w1 ),
    .ZN(\V1/V3/V1/V3/w4 ));
 XOR2_X2 \V1/V3/V1/V3/HA1/_1_  (.A(\V1/V3/V1/V3/w2 ),
    .B(\V1/V3/V1/V3/w1 ),
    .Z(\V1/V3/V1/v3 [1]));
 AND2_X1 \V1/V3/V1/V3/HA2/_0_  (.A1(\V1/V3/V1/V3/w4 ),
    .A2(\V1/V3/V1/V3/w3 ),
    .ZN(\V1/V3/V1/v3 [3]));
 XOR2_X2 \V1/V3/V1/V3/HA2/_1_  (.A(\V1/V3/V1/V3/w4 ),
    .B(\V1/V3/V1/V3/w3 ),
    .Z(\V1/V3/V1/v3 [2]));
 AND2_X1 \V1/V3/V1/V3/_0_  (.A1(A[0]),
    .A2(B[10]),
    .ZN(\V1/V3/V1/v3 [0]));
 AND2_X1 \V1/V3/V1/V3/_1_  (.A1(A[0]),
    .A2(B[11]),
    .ZN(\V1/V3/V1/V3/w1 ));
 AND2_X1 \V1/V3/V1/V3/_2_  (.A1(B[10]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V3/w2 ));
 AND2_X1 \V1/V3/V1/V3/_3_  (.A1(B[11]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V3/w3 ));
 AND2_X1 \V1/V3/V1/V4/HA1/_0_  (.A1(\V1/V3/V1/V4/w2 ),
    .A2(\V1/V3/V1/V4/w1 ),
    .ZN(\V1/V3/V1/V4/w4 ));
 XOR2_X2 \V1/V3/V1/V4/HA1/_1_  (.A(\V1/V3/V1/V4/w2 ),
    .B(\V1/V3/V1/V4/w1 ),
    .Z(\V1/V3/V1/v4 [1]));
 AND2_X1 \V1/V3/V1/V4/HA2/_0_  (.A1(\V1/V3/V1/V4/w4 ),
    .A2(\V1/V3/V1/V4/w3 ),
    .ZN(\V1/V3/V1/v4 [3]));
 XOR2_X2 \V1/V3/V1/V4/HA2/_1_  (.A(\V1/V3/V1/V4/w4 ),
    .B(\V1/V3/V1/V4/w3 ),
    .Z(\V1/V3/V1/v4 [2]));
 AND2_X1 \V1/V3/V1/V4/_0_  (.A1(A[2]),
    .A2(B[10]),
    .ZN(\V1/V3/V1/v4 [0]));
 AND2_X1 \V1/V3/V1/V4/_1_  (.A1(A[2]),
    .A2(B[11]),
    .ZN(\V1/V3/V1/V4/w1 ));
 AND2_X1 \V1/V3/V1/V4/_2_  (.A1(B[10]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V4/w2 ));
 AND2_X1 \V1/V3/V1/V4/_3_  (.A1(B[11]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V4/w3 ));
 OR2_X1 \V1/V3/V1/_0_  (.A1(\V1/V3/V1/c1 ),
    .A2(\V1/V3/V1/c2 ),
    .ZN(\V1/V3/V1/c3 ));
 AND2_X1 \V1/V3/V2/A1/M1/M1/_0_  (.A1(\V1/V3/V2/v2 [0]),
    .A2(\V1/V3/V2/v3 [0]),
    .ZN(\V1/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M1/M1/_1_  (.A(\V1/V3/V2/v2 [0]),
    .B(\V1/V3/V2/v3 [0]),
    .Z(\V1/V3/V2/A1/M1/s1 ));
 AND2_X1 \V1/V3/V2/A1/M1/M2/_0_  (.A1(\V1/V3/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M1/M2/_1_  (.A(\V1/V3/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/V2/s1 [0]));
 OR2_X1 \V1/V3/V2/A1/M1/_0_  (.A1(\V1/V3/V2/A1/M1/c1 ),
    .A2(\V1/V3/V2/A1/M1/c2 ),
    .ZN(\V1/V3/V2/A1/c1 ));
 AND2_X1 \V1/V3/V2/A1/M2/M1/_0_  (.A1(\V1/V3/V2/v2 [1]),
    .A2(\V1/V3/V2/v3 [1]),
    .ZN(\V1/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M2/M1/_1_  (.A(\V1/V3/V2/v2 [1]),
    .B(\V1/V3/V2/v3 [1]),
    .Z(\V1/V3/V2/A1/M2/s1 ));
 AND2_X1 \V1/V3/V2/A1/M2/M2/_0_  (.A1(\V1/V3/V2/A1/M2/s1 ),
    .A2(\V1/V3/V2/A1/c1 ),
    .ZN(\V1/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M2/M2/_1_  (.A(\V1/V3/V2/A1/M2/s1 ),
    .B(\V1/V3/V2/A1/c1 ),
    .Z(\V1/V3/V2/s1 [1]));
 OR2_X1 \V1/V3/V2/A1/M2/_0_  (.A1(\V1/V3/V2/A1/M2/c1 ),
    .A2(\V1/V3/V2/A1/M2/c2 ),
    .ZN(\V1/V3/V2/A1/c2 ));
 AND2_X1 \V1/V3/V2/A1/M3/M1/_0_  (.A1(\V1/V3/V2/v2 [2]),
    .A2(\V1/V3/V2/v3 [2]),
    .ZN(\V1/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M3/M1/_1_  (.A(\V1/V3/V2/v2 [2]),
    .B(\V1/V3/V2/v3 [2]),
    .Z(\V1/V3/V2/A1/M3/s1 ));
 AND2_X1 \V1/V3/V2/A1/M3/M2/_0_  (.A1(\V1/V3/V2/A1/M3/s1 ),
    .A2(\V1/V3/V2/A1/c2 ),
    .ZN(\V1/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M3/M2/_1_  (.A(\V1/V3/V2/A1/M3/s1 ),
    .B(\V1/V3/V2/A1/c2 ),
    .Z(\V1/V3/V2/s1 [2]));
 OR2_X1 \V1/V3/V2/A1/M3/_0_  (.A1(\V1/V3/V2/A1/M3/c1 ),
    .A2(\V1/V3/V2/A1/M3/c2 ),
    .ZN(\V1/V3/V2/A1/c3 ));
 AND2_X1 \V1/V3/V2/A1/M4/M1/_0_  (.A1(\V1/V3/V2/v2 [3]),
    .A2(\V1/V3/V2/v3 [3]),
    .ZN(\V1/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M4/M1/_1_  (.A(\V1/V3/V2/v2 [3]),
    .B(\V1/V3/V2/v3 [3]),
    .Z(\V1/V3/V2/A1/M4/s1 ));
 AND2_X1 \V1/V3/V2/A1/M4/M2/_0_  (.A1(\V1/V3/V2/A1/M4/s1 ),
    .A2(\V1/V3/V2/A1/c3 ),
    .ZN(\V1/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M4/M2/_1_  (.A(\V1/V3/V2/A1/M4/s1 ),
    .B(\V1/V3/V2/A1/c3 ),
    .Z(\V1/V3/V2/s1 [3]));
 OR2_X1 \V1/V3/V2/A1/M4/_0_  (.A1(\V1/V3/V2/A1/M4/c1 ),
    .A2(\V1/V3/V2/A1/M4/c2 ),
    .ZN(\V1/V3/V2/c1 ));
 AND2_X1 \V1/V3/V2/A2/M1/M1/_0_  (.A1(\V1/V3/V2/s1 [0]),
    .A2(\V1/V3/V2/v1 [2]),
    .ZN(\V1/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M1/M1/_1_  (.A(\V1/V3/V2/s1 [0]),
    .B(\V1/V3/V2/v1 [2]),
    .Z(\V1/V3/V2/A2/M1/s1 ));
 AND2_X1 \V1/V3/V2/A2/M1/M2/_0_  (.A1(\V1/V3/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M1/M2/_1_  (.A(\V1/V3/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v2 [2]));
 OR2_X1 \V1/V3/V2/A2/M1/_0_  (.A1(\V1/V3/V2/A2/M1/c1 ),
    .A2(\V1/V3/V2/A2/M1/c2 ),
    .ZN(\V1/V3/V2/A2/c1 ));
 AND2_X1 \V1/V3/V2/A2/M2/M1/_0_  (.A1(\V1/V3/V2/s1 [1]),
    .A2(\V1/V3/V2/v1 [3]),
    .ZN(\V1/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M2/M1/_1_  (.A(\V1/V3/V2/s1 [1]),
    .B(\V1/V3/V2/v1 [3]),
    .Z(\V1/V3/V2/A2/M2/s1 ));
 AND2_X1 \V1/V3/V2/A2/M2/M2/_0_  (.A1(\V1/V3/V2/A2/M2/s1 ),
    .A2(\V1/V3/V2/A2/c1 ),
    .ZN(\V1/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M2/M2/_1_  (.A(\V1/V3/V2/A2/M2/s1 ),
    .B(\V1/V3/V2/A2/c1 ),
    .Z(\V1/V3/v2 [3]));
 OR2_X1 \V1/V3/V2/A2/M2/_0_  (.A1(\V1/V3/V2/A2/M2/c1 ),
    .A2(\V1/V3/V2/A2/M2/c2 ),
    .ZN(\V1/V3/V2/A2/c2 ));
 AND2_X1 \V1/V3/V2/A2/M3/M1/_0_  (.A1(\V1/V3/V2/s1 [2]),
    .A2(ground),
    .ZN(\V1/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M3/M1/_1_  (.A(\V1/V3/V2/s1 [2]),
    .B(ground),
    .Z(\V1/V3/V2/A2/M3/s1 ));
 AND2_X1 \V1/V3/V2/A2/M3/M2/_0_  (.A1(\V1/V3/V2/A2/M3/s1 ),
    .A2(\V1/V3/V2/A2/c2 ),
    .ZN(\V1/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M3/M2/_1_  (.A(\V1/V3/V2/A2/M3/s1 ),
    .B(\V1/V3/V2/A2/c2 ),
    .Z(\V1/V3/V2/s2 [2]));
 OR2_X1 \V1/V3/V2/A2/M3/_0_  (.A1(\V1/V3/V2/A2/M3/c1 ),
    .A2(\V1/V3/V2/A2/M3/c2 ),
    .ZN(\V1/V3/V2/A2/c3 ));
 AND2_X1 \V1/V3/V2/A2/M4/M1/_0_  (.A1(\V1/V3/V2/s1 [3]),
    .A2(ground),
    .ZN(\V1/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M4/M1/_1_  (.A(\V1/V3/V2/s1 [3]),
    .B(ground),
    .Z(\V1/V3/V2/A2/M4/s1 ));
 AND2_X1 \V1/V3/V2/A2/M4/M2/_0_  (.A1(\V1/V3/V2/A2/M4/s1 ),
    .A2(\V1/V3/V2/A2/c3 ),
    .ZN(\V1/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M4/M2/_1_  (.A(\V1/V3/V2/A2/M4/s1 ),
    .B(\V1/V3/V2/A2/c3 ),
    .Z(\V1/V3/V2/s2 [3]));
 OR2_X1 \V1/V3/V2/A2/M4/_0_  (.A1(\V1/V3/V2/A2/M4/c1 ),
    .A2(\V1/V3/V2/A2/M4/c2 ),
    .ZN(\V1/V3/V2/c2 ));
 AND2_X1 \V1/V3/V2/A3/M1/M1/_0_  (.A1(\V1/V3/V2/v4 [0]),
    .A2(\V1/V3/V2/s2 [2]),
    .ZN(\V1/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M1/M1/_1_  (.A(\V1/V3/V2/v4 [0]),
    .B(\V1/V3/V2/s2 [2]),
    .Z(\V1/V3/V2/A3/M1/s1 ));
 AND2_X1 \V1/V3/V2/A3/M1/M2/_0_  (.A1(\V1/V3/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M1/M2/_1_  (.A(\V1/V3/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v2 [4]));
 OR2_X1 \V1/V3/V2/A3/M1/_0_  (.A1(\V1/V3/V2/A3/M1/c1 ),
    .A2(\V1/V3/V2/A3/M1/c2 ),
    .ZN(\V1/V3/V2/A3/c1 ));
 AND2_X1 \V1/V3/V2/A3/M2/M1/_0_  (.A1(\V1/V3/V2/v4 [1]),
    .A2(\V1/V3/V2/s2 [3]),
    .ZN(\V1/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M2/M1/_1_  (.A(\V1/V3/V2/v4 [1]),
    .B(\V1/V3/V2/s2 [3]),
    .Z(\V1/V3/V2/A3/M2/s1 ));
 AND2_X1 \V1/V3/V2/A3/M2/M2/_0_  (.A1(\V1/V3/V2/A3/M2/s1 ),
    .A2(\V1/V3/V2/A3/c1 ),
    .ZN(\V1/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M2/M2/_1_  (.A(\V1/V3/V2/A3/M2/s1 ),
    .B(\V1/V3/V2/A3/c1 ),
    .Z(\V1/V3/v2 [5]));
 OR2_X1 \V1/V3/V2/A3/M2/_0_  (.A1(\V1/V3/V2/A3/M2/c1 ),
    .A2(\V1/V3/V2/A3/M2/c2 ),
    .ZN(\V1/V3/V2/A3/c2 ));
 AND2_X1 \V1/V3/V2/A3/M3/M1/_0_  (.A1(\V1/V3/V2/v4 [2]),
    .A2(\V1/V3/V2/c3 ),
    .ZN(\V1/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M3/M1/_1_  (.A(\V1/V3/V2/v4 [2]),
    .B(\V1/V3/V2/c3 ),
    .Z(\V1/V3/V2/A3/M3/s1 ));
 AND2_X1 \V1/V3/V2/A3/M3/M2/_0_  (.A1(\V1/V3/V2/A3/M3/s1 ),
    .A2(\V1/V3/V2/A3/c2 ),
    .ZN(\V1/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M3/M2/_1_  (.A(\V1/V3/V2/A3/M3/s1 ),
    .B(\V1/V3/V2/A3/c2 ),
    .Z(\V1/V3/v2 [6]));
 OR2_X1 \V1/V3/V2/A3/M3/_0_  (.A1(\V1/V3/V2/A3/M3/c1 ),
    .A2(\V1/V3/V2/A3/M3/c2 ),
    .ZN(\V1/V3/V2/A3/c3 ));
 AND2_X1 \V1/V3/V2/A3/M4/M1/_0_  (.A1(\V1/V3/V2/v4 [3]),
    .A2(ground),
    .ZN(\V1/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M4/M1/_1_  (.A(\V1/V3/V2/v4 [3]),
    .B(ground),
    .Z(\V1/V3/V2/A3/M4/s1 ));
 AND2_X1 \V1/V3/V2/A3/M4/M2/_0_  (.A1(\V1/V3/V2/A3/M4/s1 ),
    .A2(\V1/V3/V2/A3/c3 ),
    .ZN(\V1/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M4/M2/_1_  (.A(\V1/V3/V2/A3/M4/s1 ),
    .B(\V1/V3/V2/A3/c3 ),
    .Z(\V1/V3/v2 [7]));
 OR2_X1 \V1/V3/V2/A3/M4/_0_  (.A1(\V1/V3/V2/A3/M4/c1 ),
    .A2(\V1/V3/V2/A3/M4/c2 ),
    .ZN(\V1/V3/V2/overflow ));
 AND2_X1 \V1/V3/V2/V1/HA1/_0_  (.A1(\V1/V3/V2/V1/w2 ),
    .A2(\V1/V3/V2/V1/w1 ),
    .ZN(\V1/V3/V2/V1/w4 ));
 XOR2_X2 \V1/V3/V2/V1/HA1/_1_  (.A(\V1/V3/V2/V1/w2 ),
    .B(\V1/V3/V2/V1/w1 ),
    .Z(\V1/V3/v2 [1]));
 AND2_X1 \V1/V3/V2/V1/HA2/_0_  (.A1(\V1/V3/V2/V1/w4 ),
    .A2(\V1/V3/V2/V1/w3 ),
    .ZN(\V1/V3/V2/v1 [3]));
 XOR2_X2 \V1/V3/V2/V1/HA2/_1_  (.A(\V1/V3/V2/V1/w4 ),
    .B(\V1/V3/V2/V1/w3 ),
    .Z(\V1/V3/V2/v1 [2]));
 AND2_X1 \V1/V3/V2/V1/_0_  (.A1(A[4]),
    .A2(B[8]),
    .ZN(\V1/V3/v2 [0]));
 AND2_X1 \V1/V3/V2/V1/_1_  (.A1(A[4]),
    .A2(B[9]),
    .ZN(\V1/V3/V2/V1/w1 ));
 AND2_X1 \V1/V3/V2/V1/_2_  (.A1(B[8]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V1/w2 ));
 AND2_X1 \V1/V3/V2/V1/_3_  (.A1(B[9]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V1/w3 ));
 AND2_X1 \V1/V3/V2/V2/HA1/_0_  (.A1(\V1/V3/V2/V2/w2 ),
    .A2(\V1/V3/V2/V2/w1 ),
    .ZN(\V1/V3/V2/V2/w4 ));
 XOR2_X2 \V1/V3/V2/V2/HA1/_1_  (.A(\V1/V3/V2/V2/w2 ),
    .B(\V1/V3/V2/V2/w1 ),
    .Z(\V1/V3/V2/v2 [1]));
 AND2_X1 \V1/V3/V2/V2/HA2/_0_  (.A1(\V1/V3/V2/V2/w4 ),
    .A2(\V1/V3/V2/V2/w3 ),
    .ZN(\V1/V3/V2/v2 [3]));
 XOR2_X2 \V1/V3/V2/V2/HA2/_1_  (.A(\V1/V3/V2/V2/w4 ),
    .B(\V1/V3/V2/V2/w3 ),
    .Z(\V1/V3/V2/v2 [2]));
 AND2_X1 \V1/V3/V2/V2/_0_  (.A1(A[6]),
    .A2(B[8]),
    .ZN(\V1/V3/V2/v2 [0]));
 AND2_X1 \V1/V3/V2/V2/_1_  (.A1(A[6]),
    .A2(B[9]),
    .ZN(\V1/V3/V2/V2/w1 ));
 AND2_X1 \V1/V3/V2/V2/_2_  (.A1(B[8]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V2/w2 ));
 AND2_X1 \V1/V3/V2/V2/_3_  (.A1(B[9]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V2/w3 ));
 AND2_X1 \V1/V3/V2/V3/HA1/_0_  (.A1(\V1/V3/V2/V3/w2 ),
    .A2(\V1/V3/V2/V3/w1 ),
    .ZN(\V1/V3/V2/V3/w4 ));
 XOR2_X2 \V1/V3/V2/V3/HA1/_1_  (.A(\V1/V3/V2/V3/w2 ),
    .B(\V1/V3/V2/V3/w1 ),
    .Z(\V1/V3/V2/v3 [1]));
 AND2_X1 \V1/V3/V2/V3/HA2/_0_  (.A1(\V1/V3/V2/V3/w4 ),
    .A2(\V1/V3/V2/V3/w3 ),
    .ZN(\V1/V3/V2/v3 [3]));
 XOR2_X2 \V1/V3/V2/V3/HA2/_1_  (.A(\V1/V3/V2/V3/w4 ),
    .B(\V1/V3/V2/V3/w3 ),
    .Z(\V1/V3/V2/v3 [2]));
 AND2_X1 \V1/V3/V2/V3/_0_  (.A1(A[4]),
    .A2(B[10]),
    .ZN(\V1/V3/V2/v3 [0]));
 AND2_X1 \V1/V3/V2/V3/_1_  (.A1(A[4]),
    .A2(B[11]),
    .ZN(\V1/V3/V2/V3/w1 ));
 AND2_X1 \V1/V3/V2/V3/_2_  (.A1(B[10]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V3/w2 ));
 AND2_X1 \V1/V3/V2/V3/_3_  (.A1(B[11]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V3/w3 ));
 AND2_X1 \V1/V3/V2/V4/HA1/_0_  (.A1(\V1/V3/V2/V4/w2 ),
    .A2(\V1/V3/V2/V4/w1 ),
    .ZN(\V1/V3/V2/V4/w4 ));
 XOR2_X2 \V1/V3/V2/V4/HA1/_1_  (.A(\V1/V3/V2/V4/w2 ),
    .B(\V1/V3/V2/V4/w1 ),
    .Z(\V1/V3/V2/v4 [1]));
 AND2_X1 \V1/V3/V2/V4/HA2/_0_  (.A1(\V1/V3/V2/V4/w4 ),
    .A2(\V1/V3/V2/V4/w3 ),
    .ZN(\V1/V3/V2/v4 [3]));
 XOR2_X2 \V1/V3/V2/V4/HA2/_1_  (.A(\V1/V3/V2/V4/w4 ),
    .B(\V1/V3/V2/V4/w3 ),
    .Z(\V1/V3/V2/v4 [2]));
 AND2_X1 \V1/V3/V2/V4/_0_  (.A1(A[6]),
    .A2(B[10]),
    .ZN(\V1/V3/V2/v4 [0]));
 AND2_X1 \V1/V3/V2/V4/_1_  (.A1(A[6]),
    .A2(B[11]),
    .ZN(\V1/V3/V2/V4/w1 ));
 AND2_X1 \V1/V3/V2/V4/_2_  (.A1(B[10]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V4/w2 ));
 AND2_X1 \V1/V3/V2/V4/_3_  (.A1(B[11]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V4/w3 ));
 OR2_X1 \V1/V3/V2/_0_  (.A1(\V1/V3/V2/c1 ),
    .A2(\V1/V3/V2/c2 ),
    .ZN(\V1/V3/V2/c3 ));
 AND2_X1 \V1/V3/V3/A1/M1/M1/_0_  (.A1(\V1/V3/V3/v2 [0]),
    .A2(\V1/V3/V3/v3 [0]),
    .ZN(\V1/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M1/M1/_1_  (.A(\V1/V3/V3/v2 [0]),
    .B(\V1/V3/V3/v3 [0]),
    .Z(\V1/V3/V3/A1/M1/s1 ));
 AND2_X1 \V1/V3/V3/A1/M1/M2/_0_  (.A1(\V1/V3/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M1/M2/_1_  (.A(\V1/V3/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/V3/s1 [0]));
 OR2_X1 \V1/V3/V3/A1/M1/_0_  (.A1(\V1/V3/V3/A1/M1/c1 ),
    .A2(\V1/V3/V3/A1/M1/c2 ),
    .ZN(\V1/V3/V3/A1/c1 ));
 AND2_X1 \V1/V3/V3/A1/M2/M1/_0_  (.A1(\V1/V3/V3/v2 [1]),
    .A2(\V1/V3/V3/v3 [1]),
    .ZN(\V1/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M2/M1/_1_  (.A(\V1/V3/V3/v2 [1]),
    .B(\V1/V3/V3/v3 [1]),
    .Z(\V1/V3/V3/A1/M2/s1 ));
 AND2_X1 \V1/V3/V3/A1/M2/M2/_0_  (.A1(\V1/V3/V3/A1/M2/s1 ),
    .A2(\V1/V3/V3/A1/c1 ),
    .ZN(\V1/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M2/M2/_1_  (.A(\V1/V3/V3/A1/M2/s1 ),
    .B(\V1/V3/V3/A1/c1 ),
    .Z(\V1/V3/V3/s1 [1]));
 OR2_X1 \V1/V3/V3/A1/M2/_0_  (.A1(\V1/V3/V3/A1/M2/c1 ),
    .A2(\V1/V3/V3/A1/M2/c2 ),
    .ZN(\V1/V3/V3/A1/c2 ));
 AND2_X1 \V1/V3/V3/A1/M3/M1/_0_  (.A1(\V1/V3/V3/v2 [2]),
    .A2(\V1/V3/V3/v3 [2]),
    .ZN(\V1/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M3/M1/_1_  (.A(\V1/V3/V3/v2 [2]),
    .B(\V1/V3/V3/v3 [2]),
    .Z(\V1/V3/V3/A1/M3/s1 ));
 AND2_X1 \V1/V3/V3/A1/M3/M2/_0_  (.A1(\V1/V3/V3/A1/M3/s1 ),
    .A2(\V1/V3/V3/A1/c2 ),
    .ZN(\V1/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M3/M2/_1_  (.A(\V1/V3/V3/A1/M3/s1 ),
    .B(\V1/V3/V3/A1/c2 ),
    .Z(\V1/V3/V3/s1 [2]));
 OR2_X1 \V1/V3/V3/A1/M3/_0_  (.A1(\V1/V3/V3/A1/M3/c1 ),
    .A2(\V1/V3/V3/A1/M3/c2 ),
    .ZN(\V1/V3/V3/A1/c3 ));
 AND2_X1 \V1/V3/V3/A1/M4/M1/_0_  (.A1(\V1/V3/V3/v2 [3]),
    .A2(\V1/V3/V3/v3 [3]),
    .ZN(\V1/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M4/M1/_1_  (.A(\V1/V3/V3/v2 [3]),
    .B(\V1/V3/V3/v3 [3]),
    .Z(\V1/V3/V3/A1/M4/s1 ));
 AND2_X1 \V1/V3/V3/A1/M4/M2/_0_  (.A1(\V1/V3/V3/A1/M4/s1 ),
    .A2(\V1/V3/V3/A1/c3 ),
    .ZN(\V1/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M4/M2/_1_  (.A(\V1/V3/V3/A1/M4/s1 ),
    .B(\V1/V3/V3/A1/c3 ),
    .Z(\V1/V3/V3/s1 [3]));
 OR2_X1 \V1/V3/V3/A1/M4/_0_  (.A1(\V1/V3/V3/A1/M4/c1 ),
    .A2(\V1/V3/V3/A1/M4/c2 ),
    .ZN(\V1/V3/V3/c1 ));
 AND2_X1 \V1/V3/V3/A2/M1/M1/_0_  (.A1(\V1/V3/V3/s1 [0]),
    .A2(\V1/V3/V3/v1 [2]),
    .ZN(\V1/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M1/M1/_1_  (.A(\V1/V3/V3/s1 [0]),
    .B(\V1/V3/V3/v1 [2]),
    .Z(\V1/V3/V3/A2/M1/s1 ));
 AND2_X1 \V1/V3/V3/A2/M1/M2/_0_  (.A1(\V1/V3/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M1/M2/_1_  (.A(\V1/V3/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v3 [2]));
 OR2_X1 \V1/V3/V3/A2/M1/_0_  (.A1(\V1/V3/V3/A2/M1/c1 ),
    .A2(\V1/V3/V3/A2/M1/c2 ),
    .ZN(\V1/V3/V3/A2/c1 ));
 AND2_X1 \V1/V3/V3/A2/M2/M1/_0_  (.A1(\V1/V3/V3/s1 [1]),
    .A2(\V1/V3/V3/v1 [3]),
    .ZN(\V1/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M2/M1/_1_  (.A(\V1/V3/V3/s1 [1]),
    .B(\V1/V3/V3/v1 [3]),
    .Z(\V1/V3/V3/A2/M2/s1 ));
 AND2_X1 \V1/V3/V3/A2/M2/M2/_0_  (.A1(\V1/V3/V3/A2/M2/s1 ),
    .A2(\V1/V3/V3/A2/c1 ),
    .ZN(\V1/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M2/M2/_1_  (.A(\V1/V3/V3/A2/M2/s1 ),
    .B(\V1/V3/V3/A2/c1 ),
    .Z(\V1/V3/v3 [3]));
 OR2_X1 \V1/V3/V3/A2/M2/_0_  (.A1(\V1/V3/V3/A2/M2/c1 ),
    .A2(\V1/V3/V3/A2/M2/c2 ),
    .ZN(\V1/V3/V3/A2/c2 ));
 AND2_X1 \V1/V3/V3/A2/M3/M1/_0_  (.A1(\V1/V3/V3/s1 [2]),
    .A2(ground),
    .ZN(\V1/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M3/M1/_1_  (.A(\V1/V3/V3/s1 [2]),
    .B(ground),
    .Z(\V1/V3/V3/A2/M3/s1 ));
 AND2_X1 \V1/V3/V3/A2/M3/M2/_0_  (.A1(\V1/V3/V3/A2/M3/s1 ),
    .A2(\V1/V3/V3/A2/c2 ),
    .ZN(\V1/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M3/M2/_1_  (.A(\V1/V3/V3/A2/M3/s1 ),
    .B(\V1/V3/V3/A2/c2 ),
    .Z(\V1/V3/V3/s2 [2]));
 OR2_X1 \V1/V3/V3/A2/M3/_0_  (.A1(\V1/V3/V3/A2/M3/c1 ),
    .A2(\V1/V3/V3/A2/M3/c2 ),
    .ZN(\V1/V3/V3/A2/c3 ));
 AND2_X1 \V1/V3/V3/A2/M4/M1/_0_  (.A1(\V1/V3/V3/s1 [3]),
    .A2(ground),
    .ZN(\V1/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M4/M1/_1_  (.A(\V1/V3/V3/s1 [3]),
    .B(ground),
    .Z(\V1/V3/V3/A2/M4/s1 ));
 AND2_X1 \V1/V3/V3/A2/M4/M2/_0_  (.A1(\V1/V3/V3/A2/M4/s1 ),
    .A2(\V1/V3/V3/A2/c3 ),
    .ZN(\V1/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M4/M2/_1_  (.A(\V1/V3/V3/A2/M4/s1 ),
    .B(\V1/V3/V3/A2/c3 ),
    .Z(\V1/V3/V3/s2 [3]));
 OR2_X1 \V1/V3/V3/A2/M4/_0_  (.A1(\V1/V3/V3/A2/M4/c1 ),
    .A2(\V1/V3/V3/A2/M4/c2 ),
    .ZN(\V1/V3/V3/c2 ));
 AND2_X1 \V1/V3/V3/A3/M1/M1/_0_  (.A1(\V1/V3/V3/v4 [0]),
    .A2(\V1/V3/V3/s2 [2]),
    .ZN(\V1/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M1/M1/_1_  (.A(\V1/V3/V3/v4 [0]),
    .B(\V1/V3/V3/s2 [2]),
    .Z(\V1/V3/V3/A3/M1/s1 ));
 AND2_X1 \V1/V3/V3/A3/M1/M2/_0_  (.A1(\V1/V3/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M1/M2/_1_  (.A(\V1/V3/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v3 [4]));
 OR2_X1 \V1/V3/V3/A3/M1/_0_  (.A1(\V1/V3/V3/A3/M1/c1 ),
    .A2(\V1/V3/V3/A3/M1/c2 ),
    .ZN(\V1/V3/V3/A3/c1 ));
 AND2_X1 \V1/V3/V3/A3/M2/M1/_0_  (.A1(\V1/V3/V3/v4 [1]),
    .A2(\V1/V3/V3/s2 [3]),
    .ZN(\V1/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M2/M1/_1_  (.A(\V1/V3/V3/v4 [1]),
    .B(\V1/V3/V3/s2 [3]),
    .Z(\V1/V3/V3/A3/M2/s1 ));
 AND2_X1 \V1/V3/V3/A3/M2/M2/_0_  (.A1(\V1/V3/V3/A3/M2/s1 ),
    .A2(\V1/V3/V3/A3/c1 ),
    .ZN(\V1/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M2/M2/_1_  (.A(\V1/V3/V3/A3/M2/s1 ),
    .B(\V1/V3/V3/A3/c1 ),
    .Z(\V1/V3/v3 [5]));
 OR2_X1 \V1/V3/V3/A3/M2/_0_  (.A1(\V1/V3/V3/A3/M2/c1 ),
    .A2(\V1/V3/V3/A3/M2/c2 ),
    .ZN(\V1/V3/V3/A3/c2 ));
 AND2_X1 \V1/V3/V3/A3/M3/M1/_0_  (.A1(\V1/V3/V3/v4 [2]),
    .A2(\V1/V3/V3/c3 ),
    .ZN(\V1/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M3/M1/_1_  (.A(\V1/V3/V3/v4 [2]),
    .B(\V1/V3/V3/c3 ),
    .Z(\V1/V3/V3/A3/M3/s1 ));
 AND2_X1 \V1/V3/V3/A3/M3/M2/_0_  (.A1(\V1/V3/V3/A3/M3/s1 ),
    .A2(\V1/V3/V3/A3/c2 ),
    .ZN(\V1/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M3/M2/_1_  (.A(\V1/V3/V3/A3/M3/s1 ),
    .B(\V1/V3/V3/A3/c2 ),
    .Z(\V1/V3/v3 [6]));
 OR2_X1 \V1/V3/V3/A3/M3/_0_  (.A1(\V1/V3/V3/A3/M3/c1 ),
    .A2(\V1/V3/V3/A3/M3/c2 ),
    .ZN(\V1/V3/V3/A3/c3 ));
 AND2_X1 \V1/V3/V3/A3/M4/M1/_0_  (.A1(\V1/V3/V3/v4 [3]),
    .A2(ground),
    .ZN(\V1/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M4/M1/_1_  (.A(\V1/V3/V3/v4 [3]),
    .B(ground),
    .Z(\V1/V3/V3/A3/M4/s1 ));
 AND2_X1 \V1/V3/V3/A3/M4/M2/_0_  (.A1(\V1/V3/V3/A3/M4/s1 ),
    .A2(\V1/V3/V3/A3/c3 ),
    .ZN(\V1/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M4/M2/_1_  (.A(\V1/V3/V3/A3/M4/s1 ),
    .B(\V1/V3/V3/A3/c3 ),
    .Z(\V1/V3/v3 [7]));
 OR2_X1 \V1/V3/V3/A3/M4/_0_  (.A1(\V1/V3/V3/A3/M4/c1 ),
    .A2(\V1/V3/V3/A3/M4/c2 ),
    .ZN(\V1/V3/V3/overflow ));
 AND2_X1 \V1/V3/V3/V1/HA1/_0_  (.A1(\V1/V3/V3/V1/w2 ),
    .A2(\V1/V3/V3/V1/w1 ),
    .ZN(\V1/V3/V3/V1/w4 ));
 XOR2_X2 \V1/V3/V3/V1/HA1/_1_  (.A(\V1/V3/V3/V1/w2 ),
    .B(\V1/V3/V3/V1/w1 ),
    .Z(\V1/V3/v3 [1]));
 AND2_X1 \V1/V3/V3/V1/HA2/_0_  (.A1(\V1/V3/V3/V1/w4 ),
    .A2(\V1/V3/V3/V1/w3 ),
    .ZN(\V1/V3/V3/v1 [3]));
 XOR2_X2 \V1/V3/V3/V1/HA2/_1_  (.A(\V1/V3/V3/V1/w4 ),
    .B(\V1/V3/V3/V1/w3 ),
    .Z(\V1/V3/V3/v1 [2]));
 AND2_X1 \V1/V3/V3/V1/_0_  (.A1(A[0]),
    .A2(B[12]),
    .ZN(\V1/V3/v3 [0]));
 AND2_X1 \V1/V3/V3/V1/_1_  (.A1(A[0]),
    .A2(B[13]),
    .ZN(\V1/V3/V3/V1/w1 ));
 AND2_X1 \V1/V3/V3/V1/_2_  (.A1(B[12]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V1/w2 ));
 AND2_X1 \V1/V3/V3/V1/_3_  (.A1(B[13]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V1/w3 ));
 AND2_X1 \V1/V3/V3/V2/HA1/_0_  (.A1(\V1/V3/V3/V2/w2 ),
    .A2(\V1/V3/V3/V2/w1 ),
    .ZN(\V1/V3/V3/V2/w4 ));
 XOR2_X2 \V1/V3/V3/V2/HA1/_1_  (.A(\V1/V3/V3/V2/w2 ),
    .B(\V1/V3/V3/V2/w1 ),
    .Z(\V1/V3/V3/v2 [1]));
 AND2_X1 \V1/V3/V3/V2/HA2/_0_  (.A1(\V1/V3/V3/V2/w4 ),
    .A2(\V1/V3/V3/V2/w3 ),
    .ZN(\V1/V3/V3/v2 [3]));
 XOR2_X2 \V1/V3/V3/V2/HA2/_1_  (.A(\V1/V3/V3/V2/w4 ),
    .B(\V1/V3/V3/V2/w3 ),
    .Z(\V1/V3/V3/v2 [2]));
 AND2_X1 \V1/V3/V3/V2/_0_  (.A1(A[2]),
    .A2(B[12]),
    .ZN(\V1/V3/V3/v2 [0]));
 AND2_X1 \V1/V3/V3/V2/_1_  (.A1(A[2]),
    .A2(B[13]),
    .ZN(\V1/V3/V3/V2/w1 ));
 AND2_X1 \V1/V3/V3/V2/_2_  (.A1(B[12]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V2/w2 ));
 AND2_X1 \V1/V3/V3/V2/_3_  (.A1(B[13]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V2/w3 ));
 AND2_X1 \V1/V3/V3/V3/HA1/_0_  (.A1(\V1/V3/V3/V3/w2 ),
    .A2(\V1/V3/V3/V3/w1 ),
    .ZN(\V1/V3/V3/V3/w4 ));
 XOR2_X2 \V1/V3/V3/V3/HA1/_1_  (.A(\V1/V3/V3/V3/w2 ),
    .B(\V1/V3/V3/V3/w1 ),
    .Z(\V1/V3/V3/v3 [1]));
 AND2_X1 \V1/V3/V3/V3/HA2/_0_  (.A1(\V1/V3/V3/V3/w4 ),
    .A2(\V1/V3/V3/V3/w3 ),
    .ZN(\V1/V3/V3/v3 [3]));
 XOR2_X2 \V1/V3/V3/V3/HA2/_1_  (.A(\V1/V3/V3/V3/w4 ),
    .B(\V1/V3/V3/V3/w3 ),
    .Z(\V1/V3/V3/v3 [2]));
 AND2_X1 \V1/V3/V3/V3/_0_  (.A1(A[0]),
    .A2(B[14]),
    .ZN(\V1/V3/V3/v3 [0]));
 AND2_X1 \V1/V3/V3/V3/_1_  (.A1(A[0]),
    .A2(B[15]),
    .ZN(\V1/V3/V3/V3/w1 ));
 AND2_X1 \V1/V3/V3/V3/_2_  (.A1(B[14]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V3/w2 ));
 AND2_X1 \V1/V3/V3/V3/_3_  (.A1(B[15]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V3/w3 ));
 AND2_X1 \V1/V3/V3/V4/HA1/_0_  (.A1(\V1/V3/V3/V4/w2 ),
    .A2(\V1/V3/V3/V4/w1 ),
    .ZN(\V1/V3/V3/V4/w4 ));
 XOR2_X2 \V1/V3/V3/V4/HA1/_1_  (.A(\V1/V3/V3/V4/w2 ),
    .B(\V1/V3/V3/V4/w1 ),
    .Z(\V1/V3/V3/v4 [1]));
 AND2_X1 \V1/V3/V3/V4/HA2/_0_  (.A1(\V1/V3/V3/V4/w4 ),
    .A2(\V1/V3/V3/V4/w3 ),
    .ZN(\V1/V3/V3/v4 [3]));
 XOR2_X2 \V1/V3/V3/V4/HA2/_1_  (.A(\V1/V3/V3/V4/w4 ),
    .B(\V1/V3/V3/V4/w3 ),
    .Z(\V1/V3/V3/v4 [2]));
 AND2_X1 \V1/V3/V3/V4/_0_  (.A1(A[2]),
    .A2(B[14]),
    .ZN(\V1/V3/V3/v4 [0]));
 AND2_X1 \V1/V3/V3/V4/_1_  (.A1(A[2]),
    .A2(B[15]),
    .ZN(\V1/V3/V3/V4/w1 ));
 AND2_X1 \V1/V3/V3/V4/_2_  (.A1(B[14]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V4/w2 ));
 AND2_X1 \V1/V3/V3/V4/_3_  (.A1(B[15]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V4/w3 ));
 OR2_X1 \V1/V3/V3/_0_  (.A1(\V1/V3/V3/c1 ),
    .A2(\V1/V3/V3/c2 ),
    .ZN(\V1/V3/V3/c3 ));
 AND2_X1 \V1/V3/V4/A1/M1/M1/_0_  (.A1(\V1/V3/V4/v2 [0]),
    .A2(\V1/V3/V4/v3 [0]),
    .ZN(\V1/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M1/M1/_1_  (.A(\V1/V3/V4/v2 [0]),
    .B(\V1/V3/V4/v3 [0]),
    .Z(\V1/V3/V4/A1/M1/s1 ));
 AND2_X1 \V1/V3/V4/A1/M1/M2/_0_  (.A1(\V1/V3/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M1/M2/_1_  (.A(\V1/V3/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/V4/s1 [0]));
 OR2_X1 \V1/V3/V4/A1/M1/_0_  (.A1(\V1/V3/V4/A1/M1/c1 ),
    .A2(\V1/V3/V4/A1/M1/c2 ),
    .ZN(\V1/V3/V4/A1/c1 ));
 AND2_X1 \V1/V3/V4/A1/M2/M1/_0_  (.A1(\V1/V3/V4/v2 [1]),
    .A2(\V1/V3/V4/v3 [1]),
    .ZN(\V1/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M2/M1/_1_  (.A(\V1/V3/V4/v2 [1]),
    .B(\V1/V3/V4/v3 [1]),
    .Z(\V1/V3/V4/A1/M2/s1 ));
 AND2_X1 \V1/V3/V4/A1/M2/M2/_0_  (.A1(\V1/V3/V4/A1/M2/s1 ),
    .A2(\V1/V3/V4/A1/c1 ),
    .ZN(\V1/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M2/M2/_1_  (.A(\V1/V3/V4/A1/M2/s1 ),
    .B(\V1/V3/V4/A1/c1 ),
    .Z(\V1/V3/V4/s1 [1]));
 OR2_X1 \V1/V3/V4/A1/M2/_0_  (.A1(\V1/V3/V4/A1/M2/c1 ),
    .A2(\V1/V3/V4/A1/M2/c2 ),
    .ZN(\V1/V3/V4/A1/c2 ));
 AND2_X1 \V1/V3/V4/A1/M3/M1/_0_  (.A1(\V1/V3/V4/v2 [2]),
    .A2(\V1/V3/V4/v3 [2]),
    .ZN(\V1/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M3/M1/_1_  (.A(\V1/V3/V4/v2 [2]),
    .B(\V1/V3/V4/v3 [2]),
    .Z(\V1/V3/V4/A1/M3/s1 ));
 AND2_X1 \V1/V3/V4/A1/M3/M2/_0_  (.A1(\V1/V3/V4/A1/M3/s1 ),
    .A2(\V1/V3/V4/A1/c2 ),
    .ZN(\V1/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M3/M2/_1_  (.A(\V1/V3/V4/A1/M3/s1 ),
    .B(\V1/V3/V4/A1/c2 ),
    .Z(\V1/V3/V4/s1 [2]));
 OR2_X1 \V1/V3/V4/A1/M3/_0_  (.A1(\V1/V3/V4/A1/M3/c1 ),
    .A2(\V1/V3/V4/A1/M3/c2 ),
    .ZN(\V1/V3/V4/A1/c3 ));
 AND2_X1 \V1/V3/V4/A1/M4/M1/_0_  (.A1(\V1/V3/V4/v2 [3]),
    .A2(\V1/V3/V4/v3 [3]),
    .ZN(\V1/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M4/M1/_1_  (.A(\V1/V3/V4/v2 [3]),
    .B(\V1/V3/V4/v3 [3]),
    .Z(\V1/V3/V4/A1/M4/s1 ));
 AND2_X1 \V1/V3/V4/A1/M4/M2/_0_  (.A1(\V1/V3/V4/A1/M4/s1 ),
    .A2(\V1/V3/V4/A1/c3 ),
    .ZN(\V1/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M4/M2/_1_  (.A(\V1/V3/V4/A1/M4/s1 ),
    .B(\V1/V3/V4/A1/c3 ),
    .Z(\V1/V3/V4/s1 [3]));
 OR2_X1 \V1/V3/V4/A1/M4/_0_  (.A1(\V1/V3/V4/A1/M4/c1 ),
    .A2(\V1/V3/V4/A1/M4/c2 ),
    .ZN(\V1/V3/V4/c1 ));
 AND2_X1 \V1/V3/V4/A2/M1/M1/_0_  (.A1(\V1/V3/V4/s1 [0]),
    .A2(\V1/V3/V4/v1 [2]),
    .ZN(\V1/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M1/M1/_1_  (.A(\V1/V3/V4/s1 [0]),
    .B(\V1/V3/V4/v1 [2]),
    .Z(\V1/V3/V4/A2/M1/s1 ));
 AND2_X1 \V1/V3/V4/A2/M1/M2/_0_  (.A1(\V1/V3/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M1/M2/_1_  (.A(\V1/V3/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v4 [2]));
 OR2_X1 \V1/V3/V4/A2/M1/_0_  (.A1(\V1/V3/V4/A2/M1/c1 ),
    .A2(\V1/V3/V4/A2/M1/c2 ),
    .ZN(\V1/V3/V4/A2/c1 ));
 AND2_X1 \V1/V3/V4/A2/M2/M1/_0_  (.A1(\V1/V3/V4/s1 [1]),
    .A2(\V1/V3/V4/v1 [3]),
    .ZN(\V1/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M2/M1/_1_  (.A(\V1/V3/V4/s1 [1]),
    .B(\V1/V3/V4/v1 [3]),
    .Z(\V1/V3/V4/A2/M2/s1 ));
 AND2_X1 \V1/V3/V4/A2/M2/M2/_0_  (.A1(\V1/V3/V4/A2/M2/s1 ),
    .A2(\V1/V3/V4/A2/c1 ),
    .ZN(\V1/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M2/M2/_1_  (.A(\V1/V3/V4/A2/M2/s1 ),
    .B(\V1/V3/V4/A2/c1 ),
    .Z(\V1/V3/v4 [3]));
 OR2_X1 \V1/V3/V4/A2/M2/_0_  (.A1(\V1/V3/V4/A2/M2/c1 ),
    .A2(\V1/V3/V4/A2/M2/c2 ),
    .ZN(\V1/V3/V4/A2/c2 ));
 AND2_X1 \V1/V3/V4/A2/M3/M1/_0_  (.A1(\V1/V3/V4/s1 [2]),
    .A2(ground),
    .ZN(\V1/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M3/M1/_1_  (.A(\V1/V3/V4/s1 [2]),
    .B(ground),
    .Z(\V1/V3/V4/A2/M3/s1 ));
 AND2_X1 \V1/V3/V4/A2/M3/M2/_0_  (.A1(\V1/V3/V4/A2/M3/s1 ),
    .A2(\V1/V3/V4/A2/c2 ),
    .ZN(\V1/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M3/M2/_1_  (.A(\V1/V3/V4/A2/M3/s1 ),
    .B(\V1/V3/V4/A2/c2 ),
    .Z(\V1/V3/V4/s2 [2]));
 OR2_X1 \V1/V3/V4/A2/M3/_0_  (.A1(\V1/V3/V4/A2/M3/c1 ),
    .A2(\V1/V3/V4/A2/M3/c2 ),
    .ZN(\V1/V3/V4/A2/c3 ));
 AND2_X1 \V1/V3/V4/A2/M4/M1/_0_  (.A1(\V1/V3/V4/s1 [3]),
    .A2(ground),
    .ZN(\V1/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M4/M1/_1_  (.A(\V1/V3/V4/s1 [3]),
    .B(ground),
    .Z(\V1/V3/V4/A2/M4/s1 ));
 AND2_X1 \V1/V3/V4/A2/M4/M2/_0_  (.A1(\V1/V3/V4/A2/M4/s1 ),
    .A2(\V1/V3/V4/A2/c3 ),
    .ZN(\V1/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M4/M2/_1_  (.A(\V1/V3/V4/A2/M4/s1 ),
    .B(\V1/V3/V4/A2/c3 ),
    .Z(\V1/V3/V4/s2 [3]));
 OR2_X1 \V1/V3/V4/A2/M4/_0_  (.A1(\V1/V3/V4/A2/M4/c1 ),
    .A2(\V1/V3/V4/A2/M4/c2 ),
    .ZN(\V1/V3/V4/c2 ));
 AND2_X1 \V1/V3/V4/A3/M1/M1/_0_  (.A1(\V1/V3/V4/v4 [0]),
    .A2(\V1/V3/V4/s2 [2]),
    .ZN(\V1/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M1/M1/_1_  (.A(\V1/V3/V4/v4 [0]),
    .B(\V1/V3/V4/s2 [2]),
    .Z(\V1/V3/V4/A3/M1/s1 ));
 AND2_X1 \V1/V3/V4/A3/M1/M2/_0_  (.A1(\V1/V3/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M1/M2/_1_  (.A(\V1/V3/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V3/v4 [4]));
 OR2_X1 \V1/V3/V4/A3/M1/_0_  (.A1(\V1/V3/V4/A3/M1/c1 ),
    .A2(\V1/V3/V4/A3/M1/c2 ),
    .ZN(\V1/V3/V4/A3/c1 ));
 AND2_X1 \V1/V3/V4/A3/M2/M1/_0_  (.A1(\V1/V3/V4/v4 [1]),
    .A2(\V1/V3/V4/s2 [3]),
    .ZN(\V1/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M2/M1/_1_  (.A(\V1/V3/V4/v4 [1]),
    .B(\V1/V3/V4/s2 [3]),
    .Z(\V1/V3/V4/A3/M2/s1 ));
 AND2_X1 \V1/V3/V4/A3/M2/M2/_0_  (.A1(\V1/V3/V4/A3/M2/s1 ),
    .A2(\V1/V3/V4/A3/c1 ),
    .ZN(\V1/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M2/M2/_1_  (.A(\V1/V3/V4/A3/M2/s1 ),
    .B(\V1/V3/V4/A3/c1 ),
    .Z(\V1/V3/v4 [5]));
 OR2_X1 \V1/V3/V4/A3/M2/_0_  (.A1(\V1/V3/V4/A3/M2/c1 ),
    .A2(\V1/V3/V4/A3/M2/c2 ),
    .ZN(\V1/V3/V4/A3/c2 ));
 AND2_X1 \V1/V3/V4/A3/M3/M1/_0_  (.A1(\V1/V3/V4/v4 [2]),
    .A2(\V1/V3/V4/c3 ),
    .ZN(\V1/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M3/M1/_1_  (.A(\V1/V3/V4/v4 [2]),
    .B(\V1/V3/V4/c3 ),
    .Z(\V1/V3/V4/A3/M3/s1 ));
 AND2_X1 \V1/V3/V4/A3/M3/M2/_0_  (.A1(\V1/V3/V4/A3/M3/s1 ),
    .A2(\V1/V3/V4/A3/c2 ),
    .ZN(\V1/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M3/M2/_1_  (.A(\V1/V3/V4/A3/M3/s1 ),
    .B(\V1/V3/V4/A3/c2 ),
    .Z(\V1/V3/v4 [6]));
 OR2_X1 \V1/V3/V4/A3/M3/_0_  (.A1(\V1/V3/V4/A3/M3/c1 ),
    .A2(\V1/V3/V4/A3/M3/c2 ),
    .ZN(\V1/V3/V4/A3/c3 ));
 AND2_X1 \V1/V3/V4/A3/M4/M1/_0_  (.A1(\V1/V3/V4/v4 [3]),
    .A2(ground),
    .ZN(\V1/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M4/M1/_1_  (.A(\V1/V3/V4/v4 [3]),
    .B(ground),
    .Z(\V1/V3/V4/A3/M4/s1 ));
 AND2_X1 \V1/V3/V4/A3/M4/M2/_0_  (.A1(\V1/V3/V4/A3/M4/s1 ),
    .A2(\V1/V3/V4/A3/c3 ),
    .ZN(\V1/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M4/M2/_1_  (.A(\V1/V3/V4/A3/M4/s1 ),
    .B(\V1/V3/V4/A3/c3 ),
    .Z(\V1/V3/v4 [7]));
 OR2_X1 \V1/V3/V4/A3/M4/_0_  (.A1(\V1/V3/V4/A3/M4/c1 ),
    .A2(\V1/V3/V4/A3/M4/c2 ),
    .ZN(\V1/V3/V4/overflow ));
 AND2_X1 \V1/V3/V4/V1/HA1/_0_  (.A1(\V1/V3/V4/V1/w2 ),
    .A2(\V1/V3/V4/V1/w1 ),
    .ZN(\V1/V3/V4/V1/w4 ));
 XOR2_X2 \V1/V3/V4/V1/HA1/_1_  (.A(\V1/V3/V4/V1/w2 ),
    .B(\V1/V3/V4/V1/w1 ),
    .Z(\V1/V3/v4 [1]));
 AND2_X1 \V1/V3/V4/V1/HA2/_0_  (.A1(\V1/V3/V4/V1/w4 ),
    .A2(\V1/V3/V4/V1/w3 ),
    .ZN(\V1/V3/V4/v1 [3]));
 XOR2_X2 \V1/V3/V4/V1/HA2/_1_  (.A(\V1/V3/V4/V1/w4 ),
    .B(\V1/V3/V4/V1/w3 ),
    .Z(\V1/V3/V4/v1 [2]));
 AND2_X1 \V1/V3/V4/V1/_0_  (.A1(A[4]),
    .A2(B[12]),
    .ZN(\V1/V3/v4 [0]));
 AND2_X1 \V1/V3/V4/V1/_1_  (.A1(A[4]),
    .A2(B[13]),
    .ZN(\V1/V3/V4/V1/w1 ));
 AND2_X1 \V1/V3/V4/V1/_2_  (.A1(B[12]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V1/w2 ));
 AND2_X1 \V1/V3/V4/V1/_3_  (.A1(B[13]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V1/w3 ));
 AND2_X1 \V1/V3/V4/V2/HA1/_0_  (.A1(\V1/V3/V4/V2/w2 ),
    .A2(\V1/V3/V4/V2/w1 ),
    .ZN(\V1/V3/V4/V2/w4 ));
 XOR2_X2 \V1/V3/V4/V2/HA1/_1_  (.A(\V1/V3/V4/V2/w2 ),
    .B(\V1/V3/V4/V2/w1 ),
    .Z(\V1/V3/V4/v2 [1]));
 AND2_X1 \V1/V3/V4/V2/HA2/_0_  (.A1(\V1/V3/V4/V2/w4 ),
    .A2(\V1/V3/V4/V2/w3 ),
    .ZN(\V1/V3/V4/v2 [3]));
 XOR2_X2 \V1/V3/V4/V2/HA2/_1_  (.A(\V1/V3/V4/V2/w4 ),
    .B(\V1/V3/V4/V2/w3 ),
    .Z(\V1/V3/V4/v2 [2]));
 AND2_X1 \V1/V3/V4/V2/_0_  (.A1(A[6]),
    .A2(B[12]),
    .ZN(\V1/V3/V4/v2 [0]));
 AND2_X1 \V1/V3/V4/V2/_1_  (.A1(A[6]),
    .A2(B[13]),
    .ZN(\V1/V3/V4/V2/w1 ));
 AND2_X1 \V1/V3/V4/V2/_2_  (.A1(B[12]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V2/w2 ));
 AND2_X1 \V1/V3/V4/V2/_3_  (.A1(B[13]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V2/w3 ));
 AND2_X1 \V1/V3/V4/V3/HA1/_0_  (.A1(\V1/V3/V4/V3/w2 ),
    .A2(\V1/V3/V4/V3/w1 ),
    .ZN(\V1/V3/V4/V3/w4 ));
 XOR2_X2 \V1/V3/V4/V3/HA1/_1_  (.A(\V1/V3/V4/V3/w2 ),
    .B(\V1/V3/V4/V3/w1 ),
    .Z(\V1/V3/V4/v3 [1]));
 AND2_X1 \V1/V3/V4/V3/HA2/_0_  (.A1(\V1/V3/V4/V3/w4 ),
    .A2(\V1/V3/V4/V3/w3 ),
    .ZN(\V1/V3/V4/v3 [3]));
 XOR2_X2 \V1/V3/V4/V3/HA2/_1_  (.A(\V1/V3/V4/V3/w4 ),
    .B(\V1/V3/V4/V3/w3 ),
    .Z(\V1/V3/V4/v3 [2]));
 AND2_X1 \V1/V3/V4/V3/_0_  (.A1(A[4]),
    .A2(B[14]),
    .ZN(\V1/V3/V4/v3 [0]));
 AND2_X1 \V1/V3/V4/V3/_1_  (.A1(A[4]),
    .A2(B[15]),
    .ZN(\V1/V3/V4/V3/w1 ));
 AND2_X1 \V1/V3/V4/V3/_2_  (.A1(B[14]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V3/w2 ));
 AND2_X1 \V1/V3/V4/V3/_3_  (.A1(B[15]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V3/w3 ));
 AND2_X1 \V1/V3/V4/V4/HA1/_0_  (.A1(\V1/V3/V4/V4/w2 ),
    .A2(\V1/V3/V4/V4/w1 ),
    .ZN(\V1/V3/V4/V4/w4 ));
 XOR2_X2 \V1/V3/V4/V4/HA1/_1_  (.A(\V1/V3/V4/V4/w2 ),
    .B(\V1/V3/V4/V4/w1 ),
    .Z(\V1/V3/V4/v4 [1]));
 AND2_X1 \V1/V3/V4/V4/HA2/_0_  (.A1(\V1/V3/V4/V4/w4 ),
    .A2(\V1/V3/V4/V4/w3 ),
    .ZN(\V1/V3/V4/v4 [3]));
 XOR2_X2 \V1/V3/V4/V4/HA2/_1_  (.A(\V1/V3/V4/V4/w4 ),
    .B(\V1/V3/V4/V4/w3 ),
    .Z(\V1/V3/V4/v4 [2]));
 AND2_X1 \V1/V3/V4/V4/_0_  (.A1(A[6]),
    .A2(B[14]),
    .ZN(\V1/V3/V4/v4 [0]));
 AND2_X1 \V1/V3/V4/V4/_1_  (.A1(A[6]),
    .A2(B[15]),
    .ZN(\V1/V3/V4/V4/w1 ));
 AND2_X1 \V1/V3/V4/V4/_2_  (.A1(B[14]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V4/w2 ));
 AND2_X1 \V1/V3/V4/V4/_3_  (.A1(B[15]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V4/w3 ));
 OR2_X1 \V1/V3/V4/_0_  (.A1(\V1/V3/V4/c1 ),
    .A2(\V1/V3/V4/c2 ),
    .ZN(\V1/V3/V4/c3 ));
 OR2_X1 \V1/V3/_0_  (.A1(\V1/V3/c1 ),
    .A2(\V1/V3/c2 ),
    .ZN(\V1/V3/c3 ));
 AND2_X1 \V1/V4/A1/A1/M1/M1/_0_  (.A1(\V1/V4/v2 [0]),
    .A2(\V1/V4/v3 [0]),
    .ZN(\V1/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M1/M1/_1_  (.A(\V1/V4/v2 [0]),
    .B(\V1/V4/v3 [0]),
    .Z(\V1/V4/A1/A1/M1/s1 ));
 AND2_X1 \V1/V4/A1/A1/M1/M2/_0_  (.A1(\V1/V4/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M1/M2/_1_  (.A(\V1/V4/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/s1 [0]));
 OR2_X1 \V1/V4/A1/A1/M1/_0_  (.A1(\V1/V4/A1/A1/M1/c1 ),
    .A2(\V1/V4/A1/A1/M1/c2 ),
    .ZN(\V1/V4/A1/A1/c1 ));
 AND2_X1 \V1/V4/A1/A1/M2/M1/_0_  (.A1(\V1/V4/v2 [1]),
    .A2(\V1/V4/v3 [1]),
    .ZN(\V1/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M2/M1/_1_  (.A(\V1/V4/v2 [1]),
    .B(\V1/V4/v3 [1]),
    .Z(\V1/V4/A1/A1/M2/s1 ));
 AND2_X1 \V1/V4/A1/A1/M2/M2/_0_  (.A1(\V1/V4/A1/A1/M2/s1 ),
    .A2(\V1/V4/A1/A1/c1 ),
    .ZN(\V1/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M2/M2/_1_  (.A(\V1/V4/A1/A1/M2/s1 ),
    .B(\V1/V4/A1/A1/c1 ),
    .Z(\V1/V4/s1 [1]));
 OR2_X1 \V1/V4/A1/A1/M2/_0_  (.A1(\V1/V4/A1/A1/M2/c1 ),
    .A2(\V1/V4/A1/A1/M2/c2 ),
    .ZN(\V1/V4/A1/A1/c2 ));
 AND2_X1 \V1/V4/A1/A1/M3/M1/_0_  (.A1(\V1/V4/v2 [2]),
    .A2(\V1/V4/v3 [2]),
    .ZN(\V1/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M3/M1/_1_  (.A(\V1/V4/v2 [2]),
    .B(\V1/V4/v3 [2]),
    .Z(\V1/V4/A1/A1/M3/s1 ));
 AND2_X1 \V1/V4/A1/A1/M3/M2/_0_  (.A1(\V1/V4/A1/A1/M3/s1 ),
    .A2(\V1/V4/A1/A1/c2 ),
    .ZN(\V1/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M3/M2/_1_  (.A(\V1/V4/A1/A1/M3/s1 ),
    .B(\V1/V4/A1/A1/c2 ),
    .Z(\V1/V4/s1 [2]));
 OR2_X1 \V1/V4/A1/A1/M3/_0_  (.A1(\V1/V4/A1/A1/M3/c1 ),
    .A2(\V1/V4/A1/A1/M3/c2 ),
    .ZN(\V1/V4/A1/A1/c3 ));
 AND2_X1 \V1/V4/A1/A1/M4/M1/_0_  (.A1(\V1/V4/v2 [3]),
    .A2(\V1/V4/v3 [3]),
    .ZN(\V1/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M4/M1/_1_  (.A(\V1/V4/v2 [3]),
    .B(\V1/V4/v3 [3]),
    .Z(\V1/V4/A1/A1/M4/s1 ));
 AND2_X1 \V1/V4/A1/A1/M4/M2/_0_  (.A1(\V1/V4/A1/A1/M4/s1 ),
    .A2(\V1/V4/A1/A1/c3 ),
    .ZN(\V1/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M4/M2/_1_  (.A(\V1/V4/A1/A1/M4/s1 ),
    .B(\V1/V4/A1/A1/c3 ),
    .Z(\V1/V4/s1 [3]));
 OR2_X1 \V1/V4/A1/A1/M4/_0_  (.A1(\V1/V4/A1/A1/M4/c1 ),
    .A2(\V1/V4/A1/A1/M4/c2 ),
    .ZN(\V1/V4/A1/c1 ));
 AND2_X1 \V1/V4/A1/A2/M1/M1/_0_  (.A1(\V1/V4/v2 [4]),
    .A2(\V1/V4/v3 [4]),
    .ZN(\V1/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M1/M1/_1_  (.A(\V1/V4/v2 [4]),
    .B(\V1/V4/v3 [4]),
    .Z(\V1/V4/A1/A2/M1/s1 ));
 AND2_X1 \V1/V4/A1/A2/M1/M2/_0_  (.A1(\V1/V4/A1/A2/M1/s1 ),
    .A2(\V1/V4/A1/c1 ),
    .ZN(\V1/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M1/M2/_1_  (.A(\V1/V4/A1/A2/M1/s1 ),
    .B(\V1/V4/A1/c1 ),
    .Z(\V1/V4/s1 [4]));
 OR2_X1 \V1/V4/A1/A2/M1/_0_  (.A1(\V1/V4/A1/A2/M1/c1 ),
    .A2(\V1/V4/A1/A2/M1/c2 ),
    .ZN(\V1/V4/A1/A2/c1 ));
 AND2_X1 \V1/V4/A1/A2/M2/M1/_0_  (.A1(\V1/V4/v2 [5]),
    .A2(\V1/V4/v3 [5]),
    .ZN(\V1/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M2/M1/_1_  (.A(\V1/V4/v2 [5]),
    .B(\V1/V4/v3 [5]),
    .Z(\V1/V4/A1/A2/M2/s1 ));
 AND2_X1 \V1/V4/A1/A2/M2/M2/_0_  (.A1(\V1/V4/A1/A2/M2/s1 ),
    .A2(\V1/V4/A1/A2/c1 ),
    .ZN(\V1/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M2/M2/_1_  (.A(\V1/V4/A1/A2/M2/s1 ),
    .B(\V1/V4/A1/A2/c1 ),
    .Z(\V1/V4/s1 [5]));
 OR2_X1 \V1/V4/A1/A2/M2/_0_  (.A1(\V1/V4/A1/A2/M2/c1 ),
    .A2(\V1/V4/A1/A2/M2/c2 ),
    .ZN(\V1/V4/A1/A2/c2 ));
 AND2_X1 \V1/V4/A1/A2/M3/M1/_0_  (.A1(\V1/V4/v2 [6]),
    .A2(\V1/V4/v3 [6]),
    .ZN(\V1/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M3/M1/_1_  (.A(\V1/V4/v2 [6]),
    .B(\V1/V4/v3 [6]),
    .Z(\V1/V4/A1/A2/M3/s1 ));
 AND2_X1 \V1/V4/A1/A2/M3/M2/_0_  (.A1(\V1/V4/A1/A2/M3/s1 ),
    .A2(\V1/V4/A1/A2/c2 ),
    .ZN(\V1/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M3/M2/_1_  (.A(\V1/V4/A1/A2/M3/s1 ),
    .B(\V1/V4/A1/A2/c2 ),
    .Z(\V1/V4/s1 [6]));
 OR2_X1 \V1/V4/A1/A2/M3/_0_  (.A1(\V1/V4/A1/A2/M3/c1 ),
    .A2(\V1/V4/A1/A2/M3/c2 ),
    .ZN(\V1/V4/A1/A2/c3 ));
 AND2_X1 \V1/V4/A1/A2/M4/M1/_0_  (.A1(\V1/V4/v2 [7]),
    .A2(\V1/V4/v3 [7]),
    .ZN(\V1/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M4/M1/_1_  (.A(\V1/V4/v2 [7]),
    .B(\V1/V4/v3 [7]),
    .Z(\V1/V4/A1/A2/M4/s1 ));
 AND2_X1 \V1/V4/A1/A2/M4/M2/_0_  (.A1(\V1/V4/A1/A2/M4/s1 ),
    .A2(\V1/V4/A1/A2/c3 ),
    .ZN(\V1/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M4/M2/_1_  (.A(\V1/V4/A1/A2/M4/s1 ),
    .B(\V1/V4/A1/A2/c3 ),
    .Z(\V1/V4/s1 [7]));
 OR2_X1 \V1/V4/A1/A2/M4/_0_  (.A1(\V1/V4/A1/A2/M4/c1 ),
    .A2(\V1/V4/A1/A2/M4/c2 ),
    .ZN(\V1/V4/c1 ));
 AND2_X1 \V1/V4/A2/A1/M1/M1/_0_  (.A1(\V1/V4/s1 [0]),
    .A2(\V1/V4/v1 [4]),
    .ZN(\V1/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M1/M1/_1_  (.A(\V1/V4/s1 [0]),
    .B(\V1/V4/v1 [4]),
    .Z(\V1/V4/A2/A1/M1/s1 ));
 AND2_X1 \V1/V4/A2/A1/M1/M2/_0_  (.A1(\V1/V4/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M1/M2/_1_  (.A(\V1/V4/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v4 [4]));
 OR2_X1 \V1/V4/A2/A1/M1/_0_  (.A1(\V1/V4/A2/A1/M1/c1 ),
    .A2(\V1/V4/A2/A1/M1/c2 ),
    .ZN(\V1/V4/A2/A1/c1 ));
 AND2_X1 \V1/V4/A2/A1/M2/M1/_0_  (.A1(\V1/V4/s1 [1]),
    .A2(\V1/V4/v1 [5]),
    .ZN(\V1/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M2/M1/_1_  (.A(\V1/V4/s1 [1]),
    .B(\V1/V4/v1 [5]),
    .Z(\V1/V4/A2/A1/M2/s1 ));
 AND2_X1 \V1/V4/A2/A1/M2/M2/_0_  (.A1(\V1/V4/A2/A1/M2/s1 ),
    .A2(\V1/V4/A2/A1/c1 ),
    .ZN(\V1/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M2/M2/_1_  (.A(\V1/V4/A2/A1/M2/s1 ),
    .B(\V1/V4/A2/A1/c1 ),
    .Z(\V1/v4 [5]));
 OR2_X1 \V1/V4/A2/A1/M2/_0_  (.A1(\V1/V4/A2/A1/M2/c1 ),
    .A2(\V1/V4/A2/A1/M2/c2 ),
    .ZN(\V1/V4/A2/A1/c2 ));
 AND2_X1 \V1/V4/A2/A1/M3/M1/_0_  (.A1(\V1/V4/s1 [2]),
    .A2(\V1/V4/v1 [6]),
    .ZN(\V1/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M3/M1/_1_  (.A(\V1/V4/s1 [2]),
    .B(\V1/V4/v1 [6]),
    .Z(\V1/V4/A2/A1/M3/s1 ));
 AND2_X1 \V1/V4/A2/A1/M3/M2/_0_  (.A1(\V1/V4/A2/A1/M3/s1 ),
    .A2(\V1/V4/A2/A1/c2 ),
    .ZN(\V1/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M3/M2/_1_  (.A(\V1/V4/A2/A1/M3/s1 ),
    .B(\V1/V4/A2/A1/c2 ),
    .Z(\V1/v4 [6]));
 OR2_X1 \V1/V4/A2/A1/M3/_0_  (.A1(\V1/V4/A2/A1/M3/c1 ),
    .A2(\V1/V4/A2/A1/M3/c2 ),
    .ZN(\V1/V4/A2/A1/c3 ));
 AND2_X1 \V1/V4/A2/A1/M4/M1/_0_  (.A1(\V1/V4/s1 [3]),
    .A2(\V1/V4/v1 [7]),
    .ZN(\V1/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M4/M1/_1_  (.A(\V1/V4/s1 [3]),
    .B(\V1/V4/v1 [7]),
    .Z(\V1/V4/A2/A1/M4/s1 ));
 AND2_X1 \V1/V4/A2/A1/M4/M2/_0_  (.A1(\V1/V4/A2/A1/M4/s1 ),
    .A2(\V1/V4/A2/A1/c3 ),
    .ZN(\V1/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M4/M2/_1_  (.A(\V1/V4/A2/A1/M4/s1 ),
    .B(\V1/V4/A2/A1/c3 ),
    .Z(\V1/v4 [7]));
 OR2_X1 \V1/V4/A2/A1/M4/_0_  (.A1(\V1/V4/A2/A1/M4/c1 ),
    .A2(\V1/V4/A2/A1/M4/c2 ),
    .ZN(\V1/V4/A2/c1 ));
 AND2_X1 \V1/V4/A2/A2/M1/M1/_0_  (.A1(\V1/V4/s1 [4]),
    .A2(ground),
    .ZN(\V1/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M1/M1/_1_  (.A(\V1/V4/s1 [4]),
    .B(ground),
    .Z(\V1/V4/A2/A2/M1/s1 ));
 AND2_X1 \V1/V4/A2/A2/M1/M2/_0_  (.A1(\V1/V4/A2/A2/M1/s1 ),
    .A2(\V1/V4/A2/c1 ),
    .ZN(\V1/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M1/M2/_1_  (.A(\V1/V4/A2/A2/M1/s1 ),
    .B(\V1/V4/A2/c1 ),
    .Z(\V1/V4/s2 [4]));
 OR2_X1 \V1/V4/A2/A2/M1/_0_  (.A1(\V1/V4/A2/A2/M1/c1 ),
    .A2(\V1/V4/A2/A2/M1/c2 ),
    .ZN(\V1/V4/A2/A2/c1 ));
 AND2_X1 \V1/V4/A2/A2/M2/M1/_0_  (.A1(\V1/V4/s1 [5]),
    .A2(ground),
    .ZN(\V1/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M2/M1/_1_  (.A(\V1/V4/s1 [5]),
    .B(ground),
    .Z(\V1/V4/A2/A2/M2/s1 ));
 AND2_X1 \V1/V4/A2/A2/M2/M2/_0_  (.A1(\V1/V4/A2/A2/M2/s1 ),
    .A2(\V1/V4/A2/A2/c1 ),
    .ZN(\V1/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M2/M2/_1_  (.A(\V1/V4/A2/A2/M2/s1 ),
    .B(\V1/V4/A2/A2/c1 ),
    .Z(\V1/V4/s2 [5]));
 OR2_X1 \V1/V4/A2/A2/M2/_0_  (.A1(\V1/V4/A2/A2/M2/c1 ),
    .A2(\V1/V4/A2/A2/M2/c2 ),
    .ZN(\V1/V4/A2/A2/c2 ));
 AND2_X1 \V1/V4/A2/A2/M3/M1/_0_  (.A1(\V1/V4/s1 [6]),
    .A2(ground),
    .ZN(\V1/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M3/M1/_1_  (.A(\V1/V4/s1 [6]),
    .B(ground),
    .Z(\V1/V4/A2/A2/M3/s1 ));
 AND2_X1 \V1/V4/A2/A2/M3/M2/_0_  (.A1(\V1/V4/A2/A2/M3/s1 ),
    .A2(\V1/V4/A2/A2/c2 ),
    .ZN(\V1/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M3/M2/_1_  (.A(\V1/V4/A2/A2/M3/s1 ),
    .B(\V1/V4/A2/A2/c2 ),
    .Z(\V1/V4/s2 [6]));
 OR2_X1 \V1/V4/A2/A2/M3/_0_  (.A1(\V1/V4/A2/A2/M3/c1 ),
    .A2(\V1/V4/A2/A2/M3/c2 ),
    .ZN(\V1/V4/A2/A2/c3 ));
 AND2_X1 \V1/V4/A2/A2/M4/M1/_0_  (.A1(\V1/V4/s1 [7]),
    .A2(ground),
    .ZN(\V1/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M4/M1/_1_  (.A(\V1/V4/s1 [7]),
    .B(ground),
    .Z(\V1/V4/A2/A2/M4/s1 ));
 AND2_X1 \V1/V4/A2/A2/M4/M2/_0_  (.A1(\V1/V4/A2/A2/M4/s1 ),
    .A2(\V1/V4/A2/A2/c3 ),
    .ZN(\V1/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M4/M2/_1_  (.A(\V1/V4/A2/A2/M4/s1 ),
    .B(\V1/V4/A2/A2/c3 ),
    .Z(\V1/V4/s2 [7]));
 OR2_X1 \V1/V4/A2/A2/M4/_0_  (.A1(\V1/V4/A2/A2/M4/c1 ),
    .A2(\V1/V4/A2/A2/M4/c2 ),
    .ZN(\V1/V4/c2 ));
 AND2_X1 \V1/V4/A3/A1/M1/M1/_0_  (.A1(\V1/V4/v4 [0]),
    .A2(\V1/V4/s2 [4]),
    .ZN(\V1/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M1/M1/_1_  (.A(\V1/V4/v4 [0]),
    .B(\V1/V4/s2 [4]),
    .Z(\V1/V4/A3/A1/M1/s1 ));
 AND2_X1 \V1/V4/A3/A1/M1/M2/_0_  (.A1(\V1/V4/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M1/M2/_1_  (.A(\V1/V4/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/v4 [8]));
 OR2_X1 \V1/V4/A3/A1/M1/_0_  (.A1(\V1/V4/A3/A1/M1/c1 ),
    .A2(\V1/V4/A3/A1/M1/c2 ),
    .ZN(\V1/V4/A3/A1/c1 ));
 AND2_X1 \V1/V4/A3/A1/M2/M1/_0_  (.A1(\V1/V4/v4 [1]),
    .A2(\V1/V4/s2 [5]),
    .ZN(\V1/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M2/M1/_1_  (.A(\V1/V4/v4 [1]),
    .B(\V1/V4/s2 [5]),
    .Z(\V1/V4/A3/A1/M2/s1 ));
 AND2_X1 \V1/V4/A3/A1/M2/M2/_0_  (.A1(\V1/V4/A3/A1/M2/s1 ),
    .A2(\V1/V4/A3/A1/c1 ),
    .ZN(\V1/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M2/M2/_1_  (.A(\V1/V4/A3/A1/M2/s1 ),
    .B(\V1/V4/A3/A1/c1 ),
    .Z(\V1/v4 [9]));
 OR2_X1 \V1/V4/A3/A1/M2/_0_  (.A1(\V1/V4/A3/A1/M2/c1 ),
    .A2(\V1/V4/A3/A1/M2/c2 ),
    .ZN(\V1/V4/A3/A1/c2 ));
 AND2_X1 \V1/V4/A3/A1/M3/M1/_0_  (.A1(\V1/V4/v4 [2]),
    .A2(\V1/V4/s2 [6]),
    .ZN(\V1/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M3/M1/_1_  (.A(\V1/V4/v4 [2]),
    .B(\V1/V4/s2 [6]),
    .Z(\V1/V4/A3/A1/M3/s1 ));
 AND2_X1 \V1/V4/A3/A1/M3/M2/_0_  (.A1(\V1/V4/A3/A1/M3/s1 ),
    .A2(\V1/V4/A3/A1/c2 ),
    .ZN(\V1/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M3/M2/_1_  (.A(\V1/V4/A3/A1/M3/s1 ),
    .B(\V1/V4/A3/A1/c2 ),
    .Z(\V1/v4 [10]));
 OR2_X1 \V1/V4/A3/A1/M3/_0_  (.A1(\V1/V4/A3/A1/M3/c1 ),
    .A2(\V1/V4/A3/A1/M3/c2 ),
    .ZN(\V1/V4/A3/A1/c3 ));
 AND2_X1 \V1/V4/A3/A1/M4/M1/_0_  (.A1(\V1/V4/v4 [3]),
    .A2(\V1/V4/s2 [7]),
    .ZN(\V1/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M4/M1/_1_  (.A(\V1/V4/v4 [3]),
    .B(\V1/V4/s2 [7]),
    .Z(\V1/V4/A3/A1/M4/s1 ));
 AND2_X1 \V1/V4/A3/A1/M4/M2/_0_  (.A1(\V1/V4/A3/A1/M4/s1 ),
    .A2(\V1/V4/A3/A1/c3 ),
    .ZN(\V1/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M4/M2/_1_  (.A(\V1/V4/A3/A1/M4/s1 ),
    .B(\V1/V4/A3/A1/c3 ),
    .Z(\V1/v4 [11]));
 OR2_X1 \V1/V4/A3/A1/M4/_0_  (.A1(\V1/V4/A3/A1/M4/c1 ),
    .A2(\V1/V4/A3/A1/M4/c2 ),
    .ZN(\V1/V4/A3/c1 ));
 AND2_X1 \V1/V4/A3/A2/M1/M1/_0_  (.A1(\V1/V4/v4 [4]),
    .A2(\V1/V4/c3 ),
    .ZN(\V1/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M1/M1/_1_  (.A(\V1/V4/v4 [4]),
    .B(\V1/V4/c3 ),
    .Z(\V1/V4/A3/A2/M1/s1 ));
 AND2_X1 \V1/V4/A3/A2/M1/M2/_0_  (.A1(\V1/V4/A3/A2/M1/s1 ),
    .A2(\V1/V4/A3/c1 ),
    .ZN(\V1/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M1/M2/_1_  (.A(\V1/V4/A3/A2/M1/s1 ),
    .B(\V1/V4/A3/c1 ),
    .Z(\V1/v4 [12]));
 OR2_X1 \V1/V4/A3/A2/M1/_0_  (.A1(\V1/V4/A3/A2/M1/c1 ),
    .A2(\V1/V4/A3/A2/M1/c2 ),
    .ZN(\V1/V4/A3/A2/c1 ));
 AND2_X1 \V1/V4/A3/A2/M2/M1/_0_  (.A1(\V1/V4/v4 [5]),
    .A2(ground),
    .ZN(\V1/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M2/M1/_1_  (.A(\V1/V4/v4 [5]),
    .B(ground),
    .Z(\V1/V4/A3/A2/M2/s1 ));
 AND2_X1 \V1/V4/A3/A2/M2/M2/_0_  (.A1(\V1/V4/A3/A2/M2/s1 ),
    .A2(\V1/V4/A3/A2/c1 ),
    .ZN(\V1/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M2/M2/_1_  (.A(\V1/V4/A3/A2/M2/s1 ),
    .B(\V1/V4/A3/A2/c1 ),
    .Z(\V1/v4 [13]));
 OR2_X1 \V1/V4/A3/A2/M2/_0_  (.A1(\V1/V4/A3/A2/M2/c1 ),
    .A2(\V1/V4/A3/A2/M2/c2 ),
    .ZN(\V1/V4/A3/A2/c2 ));
 AND2_X1 \V1/V4/A3/A2/M3/M1/_0_  (.A1(\V1/V4/v4 [6]),
    .A2(ground),
    .ZN(\V1/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M3/M1/_1_  (.A(\V1/V4/v4 [6]),
    .B(ground),
    .Z(\V1/V4/A3/A2/M3/s1 ));
 AND2_X1 \V1/V4/A3/A2/M3/M2/_0_  (.A1(\V1/V4/A3/A2/M3/s1 ),
    .A2(\V1/V4/A3/A2/c2 ),
    .ZN(\V1/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M3/M2/_1_  (.A(\V1/V4/A3/A2/M3/s1 ),
    .B(\V1/V4/A3/A2/c2 ),
    .Z(\V1/v4 [14]));
 OR2_X1 \V1/V4/A3/A2/M3/_0_  (.A1(\V1/V4/A3/A2/M3/c1 ),
    .A2(\V1/V4/A3/A2/M3/c2 ),
    .ZN(\V1/V4/A3/A2/c3 ));
 AND2_X1 \V1/V4/A3/A2/M4/M1/_0_  (.A1(\V1/V4/v4 [7]),
    .A2(ground),
    .ZN(\V1/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M4/M1/_1_  (.A(\V1/V4/v4 [7]),
    .B(ground),
    .Z(\V1/V4/A3/A2/M4/s1 ));
 AND2_X1 \V1/V4/A3/A2/M4/M2/_0_  (.A1(\V1/V4/A3/A2/M4/s1 ),
    .A2(\V1/V4/A3/A2/c3 ),
    .ZN(\V1/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M4/M2/_1_  (.A(\V1/V4/A3/A2/M4/s1 ),
    .B(\V1/V4/A3/A2/c3 ),
    .Z(\V1/v4 [15]));
 OR2_X1 \V1/V4/A3/A2/M4/_0_  (.A1(\V1/V4/A3/A2/M4/c1 ),
    .A2(\V1/V4/A3/A2/M4/c2 ),
    .ZN(\V1/V4/overflow ));
 AND2_X1 \V1/V4/V1/A1/M1/M1/_0_  (.A1(\V1/V4/V1/v2 [0]),
    .A2(\V1/V4/V1/v3 [0]),
    .ZN(\V1/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M1/M1/_1_  (.A(\V1/V4/V1/v2 [0]),
    .B(\V1/V4/V1/v3 [0]),
    .Z(\V1/V4/V1/A1/M1/s1 ));
 AND2_X1 \V1/V4/V1/A1/M1/M2/_0_  (.A1(\V1/V4/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M1/M2/_1_  (.A(\V1/V4/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/V1/s1 [0]));
 OR2_X1 \V1/V4/V1/A1/M1/_0_  (.A1(\V1/V4/V1/A1/M1/c1 ),
    .A2(\V1/V4/V1/A1/M1/c2 ),
    .ZN(\V1/V4/V1/A1/c1 ));
 AND2_X1 \V1/V4/V1/A1/M2/M1/_0_  (.A1(\V1/V4/V1/v2 [1]),
    .A2(\V1/V4/V1/v3 [1]),
    .ZN(\V1/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M2/M1/_1_  (.A(\V1/V4/V1/v2 [1]),
    .B(\V1/V4/V1/v3 [1]),
    .Z(\V1/V4/V1/A1/M2/s1 ));
 AND2_X1 \V1/V4/V1/A1/M2/M2/_0_  (.A1(\V1/V4/V1/A1/M2/s1 ),
    .A2(\V1/V4/V1/A1/c1 ),
    .ZN(\V1/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M2/M2/_1_  (.A(\V1/V4/V1/A1/M2/s1 ),
    .B(\V1/V4/V1/A1/c1 ),
    .Z(\V1/V4/V1/s1 [1]));
 OR2_X1 \V1/V4/V1/A1/M2/_0_  (.A1(\V1/V4/V1/A1/M2/c1 ),
    .A2(\V1/V4/V1/A1/M2/c2 ),
    .ZN(\V1/V4/V1/A1/c2 ));
 AND2_X1 \V1/V4/V1/A1/M3/M1/_0_  (.A1(\V1/V4/V1/v2 [2]),
    .A2(\V1/V4/V1/v3 [2]),
    .ZN(\V1/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M3/M1/_1_  (.A(\V1/V4/V1/v2 [2]),
    .B(\V1/V4/V1/v3 [2]),
    .Z(\V1/V4/V1/A1/M3/s1 ));
 AND2_X1 \V1/V4/V1/A1/M3/M2/_0_  (.A1(\V1/V4/V1/A1/M3/s1 ),
    .A2(\V1/V4/V1/A1/c2 ),
    .ZN(\V1/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M3/M2/_1_  (.A(\V1/V4/V1/A1/M3/s1 ),
    .B(\V1/V4/V1/A1/c2 ),
    .Z(\V1/V4/V1/s1 [2]));
 OR2_X1 \V1/V4/V1/A1/M3/_0_  (.A1(\V1/V4/V1/A1/M3/c1 ),
    .A2(\V1/V4/V1/A1/M3/c2 ),
    .ZN(\V1/V4/V1/A1/c3 ));
 AND2_X1 \V1/V4/V1/A1/M4/M1/_0_  (.A1(\V1/V4/V1/v2 [3]),
    .A2(\V1/V4/V1/v3 [3]),
    .ZN(\V1/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M4/M1/_1_  (.A(\V1/V4/V1/v2 [3]),
    .B(\V1/V4/V1/v3 [3]),
    .Z(\V1/V4/V1/A1/M4/s1 ));
 AND2_X1 \V1/V4/V1/A1/M4/M2/_0_  (.A1(\V1/V4/V1/A1/M4/s1 ),
    .A2(\V1/V4/V1/A1/c3 ),
    .ZN(\V1/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M4/M2/_1_  (.A(\V1/V4/V1/A1/M4/s1 ),
    .B(\V1/V4/V1/A1/c3 ),
    .Z(\V1/V4/V1/s1 [3]));
 OR2_X1 \V1/V4/V1/A1/M4/_0_  (.A1(\V1/V4/V1/A1/M4/c1 ),
    .A2(\V1/V4/V1/A1/M4/c2 ),
    .ZN(\V1/V4/V1/c1 ));
 AND2_X1 \V1/V4/V1/A2/M1/M1/_0_  (.A1(\V1/V4/V1/s1 [0]),
    .A2(\V1/V4/V1/v1 [2]),
    .ZN(\V1/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M1/M1/_1_  (.A(\V1/V4/V1/s1 [0]),
    .B(\V1/V4/V1/v1 [2]),
    .Z(\V1/V4/V1/A2/M1/s1 ));
 AND2_X1 \V1/V4/V1/A2/M1/M2/_0_  (.A1(\V1/V4/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M1/M2/_1_  (.A(\V1/V4/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/v4 [2]));
 OR2_X1 \V1/V4/V1/A2/M1/_0_  (.A1(\V1/V4/V1/A2/M1/c1 ),
    .A2(\V1/V4/V1/A2/M1/c2 ),
    .ZN(\V1/V4/V1/A2/c1 ));
 AND2_X1 \V1/V4/V1/A2/M2/M1/_0_  (.A1(\V1/V4/V1/s1 [1]),
    .A2(\V1/V4/V1/v1 [3]),
    .ZN(\V1/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M2/M1/_1_  (.A(\V1/V4/V1/s1 [1]),
    .B(\V1/V4/V1/v1 [3]),
    .Z(\V1/V4/V1/A2/M2/s1 ));
 AND2_X1 \V1/V4/V1/A2/M2/M2/_0_  (.A1(\V1/V4/V1/A2/M2/s1 ),
    .A2(\V1/V4/V1/A2/c1 ),
    .ZN(\V1/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M2/M2/_1_  (.A(\V1/V4/V1/A2/M2/s1 ),
    .B(\V1/V4/V1/A2/c1 ),
    .Z(\V1/v4 [3]));
 OR2_X1 \V1/V4/V1/A2/M2/_0_  (.A1(\V1/V4/V1/A2/M2/c1 ),
    .A2(\V1/V4/V1/A2/M2/c2 ),
    .ZN(\V1/V4/V1/A2/c2 ));
 AND2_X1 \V1/V4/V1/A2/M3/M1/_0_  (.A1(\V1/V4/V1/s1 [2]),
    .A2(ground),
    .ZN(\V1/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M3/M1/_1_  (.A(\V1/V4/V1/s1 [2]),
    .B(ground),
    .Z(\V1/V4/V1/A2/M3/s1 ));
 AND2_X1 \V1/V4/V1/A2/M3/M2/_0_  (.A1(\V1/V4/V1/A2/M3/s1 ),
    .A2(\V1/V4/V1/A2/c2 ),
    .ZN(\V1/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M3/M2/_1_  (.A(\V1/V4/V1/A2/M3/s1 ),
    .B(\V1/V4/V1/A2/c2 ),
    .Z(\V1/V4/V1/s2 [2]));
 OR2_X1 \V1/V4/V1/A2/M3/_0_  (.A1(\V1/V4/V1/A2/M3/c1 ),
    .A2(\V1/V4/V1/A2/M3/c2 ),
    .ZN(\V1/V4/V1/A2/c3 ));
 AND2_X1 \V1/V4/V1/A2/M4/M1/_0_  (.A1(\V1/V4/V1/s1 [3]),
    .A2(ground),
    .ZN(\V1/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M4/M1/_1_  (.A(\V1/V4/V1/s1 [3]),
    .B(ground),
    .Z(\V1/V4/V1/A2/M4/s1 ));
 AND2_X1 \V1/V4/V1/A2/M4/M2/_0_  (.A1(\V1/V4/V1/A2/M4/s1 ),
    .A2(\V1/V4/V1/A2/c3 ),
    .ZN(\V1/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M4/M2/_1_  (.A(\V1/V4/V1/A2/M4/s1 ),
    .B(\V1/V4/V1/A2/c3 ),
    .Z(\V1/V4/V1/s2 [3]));
 OR2_X1 \V1/V4/V1/A2/M4/_0_  (.A1(\V1/V4/V1/A2/M4/c1 ),
    .A2(\V1/V4/V1/A2/M4/c2 ),
    .ZN(\V1/V4/V1/c2 ));
 AND2_X1 \V1/V4/V1/A3/M1/M1/_0_  (.A1(\V1/V4/V1/v4 [0]),
    .A2(\V1/V4/V1/s2 [2]),
    .ZN(\V1/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M1/M1/_1_  (.A(\V1/V4/V1/v4 [0]),
    .B(\V1/V4/V1/s2 [2]),
    .Z(\V1/V4/V1/A3/M1/s1 ));
 AND2_X1 \V1/V4/V1/A3/M1/M2/_0_  (.A1(\V1/V4/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M1/M2/_1_  (.A(\V1/V4/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v1 [4]));
 OR2_X1 \V1/V4/V1/A3/M1/_0_  (.A1(\V1/V4/V1/A3/M1/c1 ),
    .A2(\V1/V4/V1/A3/M1/c2 ),
    .ZN(\V1/V4/V1/A3/c1 ));
 AND2_X1 \V1/V4/V1/A3/M2/M1/_0_  (.A1(\V1/V4/V1/v4 [1]),
    .A2(\V1/V4/V1/s2 [3]),
    .ZN(\V1/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M2/M1/_1_  (.A(\V1/V4/V1/v4 [1]),
    .B(\V1/V4/V1/s2 [3]),
    .Z(\V1/V4/V1/A3/M2/s1 ));
 AND2_X1 \V1/V4/V1/A3/M2/M2/_0_  (.A1(\V1/V4/V1/A3/M2/s1 ),
    .A2(\V1/V4/V1/A3/c1 ),
    .ZN(\V1/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M2/M2/_1_  (.A(\V1/V4/V1/A3/M2/s1 ),
    .B(\V1/V4/V1/A3/c1 ),
    .Z(\V1/V4/v1 [5]));
 OR2_X1 \V1/V4/V1/A3/M2/_0_  (.A1(\V1/V4/V1/A3/M2/c1 ),
    .A2(\V1/V4/V1/A3/M2/c2 ),
    .ZN(\V1/V4/V1/A3/c2 ));
 AND2_X1 \V1/V4/V1/A3/M3/M1/_0_  (.A1(\V1/V4/V1/v4 [2]),
    .A2(\V1/V4/V1/c3 ),
    .ZN(\V1/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M3/M1/_1_  (.A(\V1/V4/V1/v4 [2]),
    .B(\V1/V4/V1/c3 ),
    .Z(\V1/V4/V1/A3/M3/s1 ));
 AND2_X1 \V1/V4/V1/A3/M3/M2/_0_  (.A1(\V1/V4/V1/A3/M3/s1 ),
    .A2(\V1/V4/V1/A3/c2 ),
    .ZN(\V1/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M3/M2/_1_  (.A(\V1/V4/V1/A3/M3/s1 ),
    .B(\V1/V4/V1/A3/c2 ),
    .Z(\V1/V4/v1 [6]));
 OR2_X1 \V1/V4/V1/A3/M3/_0_  (.A1(\V1/V4/V1/A3/M3/c1 ),
    .A2(\V1/V4/V1/A3/M3/c2 ),
    .ZN(\V1/V4/V1/A3/c3 ));
 AND2_X1 \V1/V4/V1/A3/M4/M1/_0_  (.A1(\V1/V4/V1/v4 [3]),
    .A2(ground),
    .ZN(\V1/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M4/M1/_1_  (.A(\V1/V4/V1/v4 [3]),
    .B(ground),
    .Z(\V1/V4/V1/A3/M4/s1 ));
 AND2_X1 \V1/V4/V1/A3/M4/M2/_0_  (.A1(\V1/V4/V1/A3/M4/s1 ),
    .A2(\V1/V4/V1/A3/c3 ),
    .ZN(\V1/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M4/M2/_1_  (.A(\V1/V4/V1/A3/M4/s1 ),
    .B(\V1/V4/V1/A3/c3 ),
    .Z(\V1/V4/v1 [7]));
 OR2_X1 \V1/V4/V1/A3/M4/_0_  (.A1(\V1/V4/V1/A3/M4/c1 ),
    .A2(\V1/V4/V1/A3/M4/c2 ),
    .ZN(\V1/V4/V1/overflow ));
 AND2_X1 \V1/V4/V1/V1/HA1/_0_  (.A1(\V1/V4/V1/V1/w2 ),
    .A2(\V1/V4/V1/V1/w1 ),
    .ZN(\V1/V4/V1/V1/w4 ));
 XOR2_X2 \V1/V4/V1/V1/HA1/_1_  (.A(\V1/V4/V1/V1/w2 ),
    .B(\V1/V4/V1/V1/w1 ),
    .Z(\V1/v4 [1]));
 AND2_X1 \V1/V4/V1/V1/HA2/_0_  (.A1(\V1/V4/V1/V1/w4 ),
    .A2(\V1/V4/V1/V1/w3 ),
    .ZN(\V1/V4/V1/v1 [3]));
 XOR2_X2 \V1/V4/V1/V1/HA2/_1_  (.A(\V1/V4/V1/V1/w4 ),
    .B(\V1/V4/V1/V1/w3 ),
    .Z(\V1/V4/V1/v1 [2]));
 AND2_X1 \V1/V4/V1/V1/_0_  (.A1(A[8]),
    .A2(B[8]),
    .ZN(\V1/v4 [0]));
 AND2_X1 \V1/V4/V1/V1/_1_  (.A1(A[8]),
    .A2(B[9]),
    .ZN(\V1/V4/V1/V1/w1 ));
 AND2_X1 \V1/V4/V1/V1/_2_  (.A1(B[8]),
    .A2(A[9]),
    .ZN(\V1/V4/V1/V1/w2 ));
 AND2_X1 \V1/V4/V1/V1/_3_  (.A1(B[9]),
    .A2(A[9]),
    .ZN(\V1/V4/V1/V1/w3 ));
 AND2_X1 \V1/V4/V1/V2/HA1/_0_  (.A1(\V1/V4/V1/V2/w2 ),
    .A2(\V1/V4/V1/V2/w1 ),
    .ZN(\V1/V4/V1/V2/w4 ));
 XOR2_X2 \V1/V4/V1/V2/HA1/_1_  (.A(\V1/V4/V1/V2/w2 ),
    .B(\V1/V4/V1/V2/w1 ),
    .Z(\V1/V4/V1/v2 [1]));
 AND2_X1 \V1/V4/V1/V2/HA2/_0_  (.A1(\V1/V4/V1/V2/w4 ),
    .A2(\V1/V4/V1/V2/w3 ),
    .ZN(\V1/V4/V1/v2 [3]));
 XOR2_X2 \V1/V4/V1/V2/HA2/_1_  (.A(\V1/V4/V1/V2/w4 ),
    .B(\V1/V4/V1/V2/w3 ),
    .Z(\V1/V4/V1/v2 [2]));
 AND2_X1 \V1/V4/V1/V2/_0_  (.A1(A[10]),
    .A2(B[8]),
    .ZN(\V1/V4/V1/v2 [0]));
 AND2_X1 \V1/V4/V1/V2/_1_  (.A1(A[10]),
    .A2(B[9]),
    .ZN(\V1/V4/V1/V2/w1 ));
 AND2_X1 \V1/V4/V1/V2/_2_  (.A1(B[8]),
    .A2(A[11]),
    .ZN(\V1/V4/V1/V2/w2 ));
 AND2_X1 \V1/V4/V1/V2/_3_  (.A1(B[9]),
    .A2(A[11]),
    .ZN(\V1/V4/V1/V2/w3 ));
 AND2_X1 \V1/V4/V1/V3/HA1/_0_  (.A1(\V1/V4/V1/V3/w2 ),
    .A2(\V1/V4/V1/V3/w1 ),
    .ZN(\V1/V4/V1/V3/w4 ));
 XOR2_X2 \V1/V4/V1/V3/HA1/_1_  (.A(\V1/V4/V1/V3/w2 ),
    .B(\V1/V4/V1/V3/w1 ),
    .Z(\V1/V4/V1/v3 [1]));
 AND2_X1 \V1/V4/V1/V3/HA2/_0_  (.A1(\V1/V4/V1/V3/w4 ),
    .A2(\V1/V4/V1/V3/w3 ),
    .ZN(\V1/V4/V1/v3 [3]));
 XOR2_X2 \V1/V4/V1/V3/HA2/_1_  (.A(\V1/V4/V1/V3/w4 ),
    .B(\V1/V4/V1/V3/w3 ),
    .Z(\V1/V4/V1/v3 [2]));
 AND2_X1 \V1/V4/V1/V3/_0_  (.A1(A[8]),
    .A2(B[10]),
    .ZN(\V1/V4/V1/v3 [0]));
 AND2_X1 \V1/V4/V1/V3/_1_  (.A1(A[8]),
    .A2(B[11]),
    .ZN(\V1/V4/V1/V3/w1 ));
 AND2_X1 \V1/V4/V1/V3/_2_  (.A1(B[10]),
    .A2(A[9]),
    .ZN(\V1/V4/V1/V3/w2 ));
 AND2_X1 \V1/V4/V1/V3/_3_  (.A1(B[11]),
    .A2(A[9]),
    .ZN(\V1/V4/V1/V3/w3 ));
 AND2_X1 \V1/V4/V1/V4/HA1/_0_  (.A1(\V1/V4/V1/V4/w2 ),
    .A2(\V1/V4/V1/V4/w1 ),
    .ZN(\V1/V4/V1/V4/w4 ));
 XOR2_X2 \V1/V4/V1/V4/HA1/_1_  (.A(\V1/V4/V1/V4/w2 ),
    .B(\V1/V4/V1/V4/w1 ),
    .Z(\V1/V4/V1/v4 [1]));
 AND2_X1 \V1/V4/V1/V4/HA2/_0_  (.A1(\V1/V4/V1/V4/w4 ),
    .A2(\V1/V4/V1/V4/w3 ),
    .ZN(\V1/V4/V1/v4 [3]));
 XOR2_X2 \V1/V4/V1/V4/HA2/_1_  (.A(\V1/V4/V1/V4/w4 ),
    .B(\V1/V4/V1/V4/w3 ),
    .Z(\V1/V4/V1/v4 [2]));
 AND2_X1 \V1/V4/V1/V4/_0_  (.A1(A[10]),
    .A2(B[10]),
    .ZN(\V1/V4/V1/v4 [0]));
 AND2_X1 \V1/V4/V1/V4/_1_  (.A1(A[10]),
    .A2(B[11]),
    .ZN(\V1/V4/V1/V4/w1 ));
 AND2_X1 \V1/V4/V1/V4/_2_  (.A1(B[10]),
    .A2(A[11]),
    .ZN(\V1/V4/V1/V4/w2 ));
 AND2_X1 \V1/V4/V1/V4/_3_  (.A1(B[11]),
    .A2(A[11]),
    .ZN(\V1/V4/V1/V4/w3 ));
 OR2_X1 \V1/V4/V1/_0_  (.A1(\V1/V4/V1/c1 ),
    .A2(\V1/V4/V1/c2 ),
    .ZN(\V1/V4/V1/c3 ));
 AND2_X1 \V1/V4/V2/A1/M1/M1/_0_  (.A1(\V1/V4/V2/v2 [0]),
    .A2(\V1/V4/V2/v3 [0]),
    .ZN(\V1/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M1/M1/_1_  (.A(\V1/V4/V2/v2 [0]),
    .B(\V1/V4/V2/v3 [0]),
    .Z(\V1/V4/V2/A1/M1/s1 ));
 AND2_X1 \V1/V4/V2/A1/M1/M2/_0_  (.A1(\V1/V4/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M1/M2/_1_  (.A(\V1/V4/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/V2/s1 [0]));
 OR2_X1 \V1/V4/V2/A1/M1/_0_  (.A1(\V1/V4/V2/A1/M1/c1 ),
    .A2(\V1/V4/V2/A1/M1/c2 ),
    .ZN(\V1/V4/V2/A1/c1 ));
 AND2_X1 \V1/V4/V2/A1/M2/M1/_0_  (.A1(\V1/V4/V2/v2 [1]),
    .A2(\V1/V4/V2/v3 [1]),
    .ZN(\V1/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M2/M1/_1_  (.A(\V1/V4/V2/v2 [1]),
    .B(\V1/V4/V2/v3 [1]),
    .Z(\V1/V4/V2/A1/M2/s1 ));
 AND2_X1 \V1/V4/V2/A1/M2/M2/_0_  (.A1(\V1/V4/V2/A1/M2/s1 ),
    .A2(\V1/V4/V2/A1/c1 ),
    .ZN(\V1/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M2/M2/_1_  (.A(\V1/V4/V2/A1/M2/s1 ),
    .B(\V1/V4/V2/A1/c1 ),
    .Z(\V1/V4/V2/s1 [1]));
 OR2_X1 \V1/V4/V2/A1/M2/_0_  (.A1(\V1/V4/V2/A1/M2/c1 ),
    .A2(\V1/V4/V2/A1/M2/c2 ),
    .ZN(\V1/V4/V2/A1/c2 ));
 AND2_X1 \V1/V4/V2/A1/M3/M1/_0_  (.A1(\V1/V4/V2/v2 [2]),
    .A2(\V1/V4/V2/v3 [2]),
    .ZN(\V1/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M3/M1/_1_  (.A(\V1/V4/V2/v2 [2]),
    .B(\V1/V4/V2/v3 [2]),
    .Z(\V1/V4/V2/A1/M3/s1 ));
 AND2_X1 \V1/V4/V2/A1/M3/M2/_0_  (.A1(\V1/V4/V2/A1/M3/s1 ),
    .A2(\V1/V4/V2/A1/c2 ),
    .ZN(\V1/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M3/M2/_1_  (.A(\V1/V4/V2/A1/M3/s1 ),
    .B(\V1/V4/V2/A1/c2 ),
    .Z(\V1/V4/V2/s1 [2]));
 OR2_X1 \V1/V4/V2/A1/M3/_0_  (.A1(\V1/V4/V2/A1/M3/c1 ),
    .A2(\V1/V4/V2/A1/M3/c2 ),
    .ZN(\V1/V4/V2/A1/c3 ));
 AND2_X1 \V1/V4/V2/A1/M4/M1/_0_  (.A1(\V1/V4/V2/v2 [3]),
    .A2(\V1/V4/V2/v3 [3]),
    .ZN(\V1/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M4/M1/_1_  (.A(\V1/V4/V2/v2 [3]),
    .B(\V1/V4/V2/v3 [3]),
    .Z(\V1/V4/V2/A1/M4/s1 ));
 AND2_X1 \V1/V4/V2/A1/M4/M2/_0_  (.A1(\V1/V4/V2/A1/M4/s1 ),
    .A2(\V1/V4/V2/A1/c3 ),
    .ZN(\V1/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M4/M2/_1_  (.A(\V1/V4/V2/A1/M4/s1 ),
    .B(\V1/V4/V2/A1/c3 ),
    .Z(\V1/V4/V2/s1 [3]));
 OR2_X1 \V1/V4/V2/A1/M4/_0_  (.A1(\V1/V4/V2/A1/M4/c1 ),
    .A2(\V1/V4/V2/A1/M4/c2 ),
    .ZN(\V1/V4/V2/c1 ));
 AND2_X1 \V1/V4/V2/A2/M1/M1/_0_  (.A1(\V1/V4/V2/s1 [0]),
    .A2(\V1/V4/V2/v1 [2]),
    .ZN(\V1/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M1/M1/_1_  (.A(\V1/V4/V2/s1 [0]),
    .B(\V1/V4/V2/v1 [2]),
    .Z(\V1/V4/V2/A2/M1/s1 ));
 AND2_X1 \V1/V4/V2/A2/M1/M2/_0_  (.A1(\V1/V4/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M1/M2/_1_  (.A(\V1/V4/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v2 [2]));
 OR2_X1 \V1/V4/V2/A2/M1/_0_  (.A1(\V1/V4/V2/A2/M1/c1 ),
    .A2(\V1/V4/V2/A2/M1/c2 ),
    .ZN(\V1/V4/V2/A2/c1 ));
 AND2_X1 \V1/V4/V2/A2/M2/M1/_0_  (.A1(\V1/V4/V2/s1 [1]),
    .A2(\V1/V4/V2/v1 [3]),
    .ZN(\V1/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M2/M1/_1_  (.A(\V1/V4/V2/s1 [1]),
    .B(\V1/V4/V2/v1 [3]),
    .Z(\V1/V4/V2/A2/M2/s1 ));
 AND2_X1 \V1/V4/V2/A2/M2/M2/_0_  (.A1(\V1/V4/V2/A2/M2/s1 ),
    .A2(\V1/V4/V2/A2/c1 ),
    .ZN(\V1/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M2/M2/_1_  (.A(\V1/V4/V2/A2/M2/s1 ),
    .B(\V1/V4/V2/A2/c1 ),
    .Z(\V1/V4/v2 [3]));
 OR2_X1 \V1/V4/V2/A2/M2/_0_  (.A1(\V1/V4/V2/A2/M2/c1 ),
    .A2(\V1/V4/V2/A2/M2/c2 ),
    .ZN(\V1/V4/V2/A2/c2 ));
 AND2_X1 \V1/V4/V2/A2/M3/M1/_0_  (.A1(\V1/V4/V2/s1 [2]),
    .A2(ground),
    .ZN(\V1/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M3/M1/_1_  (.A(\V1/V4/V2/s1 [2]),
    .B(ground),
    .Z(\V1/V4/V2/A2/M3/s1 ));
 AND2_X1 \V1/V4/V2/A2/M3/M2/_0_  (.A1(\V1/V4/V2/A2/M3/s1 ),
    .A2(\V1/V4/V2/A2/c2 ),
    .ZN(\V1/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M3/M2/_1_  (.A(\V1/V4/V2/A2/M3/s1 ),
    .B(\V1/V4/V2/A2/c2 ),
    .Z(\V1/V4/V2/s2 [2]));
 OR2_X1 \V1/V4/V2/A2/M3/_0_  (.A1(\V1/V4/V2/A2/M3/c1 ),
    .A2(\V1/V4/V2/A2/M3/c2 ),
    .ZN(\V1/V4/V2/A2/c3 ));
 AND2_X1 \V1/V4/V2/A2/M4/M1/_0_  (.A1(\V1/V4/V2/s1 [3]),
    .A2(ground),
    .ZN(\V1/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M4/M1/_1_  (.A(\V1/V4/V2/s1 [3]),
    .B(ground),
    .Z(\V1/V4/V2/A2/M4/s1 ));
 AND2_X1 \V1/V4/V2/A2/M4/M2/_0_  (.A1(\V1/V4/V2/A2/M4/s1 ),
    .A2(\V1/V4/V2/A2/c3 ),
    .ZN(\V1/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M4/M2/_1_  (.A(\V1/V4/V2/A2/M4/s1 ),
    .B(\V1/V4/V2/A2/c3 ),
    .Z(\V1/V4/V2/s2 [3]));
 OR2_X1 \V1/V4/V2/A2/M4/_0_  (.A1(\V1/V4/V2/A2/M4/c1 ),
    .A2(\V1/V4/V2/A2/M4/c2 ),
    .ZN(\V1/V4/V2/c2 ));
 AND2_X1 \V1/V4/V2/A3/M1/M1/_0_  (.A1(\V1/V4/V2/v4 [0]),
    .A2(\V1/V4/V2/s2 [2]),
    .ZN(\V1/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M1/M1/_1_  (.A(\V1/V4/V2/v4 [0]),
    .B(\V1/V4/V2/s2 [2]),
    .Z(\V1/V4/V2/A3/M1/s1 ));
 AND2_X1 \V1/V4/V2/A3/M1/M2/_0_  (.A1(\V1/V4/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M1/M2/_1_  (.A(\V1/V4/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v2 [4]));
 OR2_X1 \V1/V4/V2/A3/M1/_0_  (.A1(\V1/V4/V2/A3/M1/c1 ),
    .A2(\V1/V4/V2/A3/M1/c2 ),
    .ZN(\V1/V4/V2/A3/c1 ));
 AND2_X1 \V1/V4/V2/A3/M2/M1/_0_  (.A1(\V1/V4/V2/v4 [1]),
    .A2(\V1/V4/V2/s2 [3]),
    .ZN(\V1/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M2/M1/_1_  (.A(\V1/V4/V2/v4 [1]),
    .B(\V1/V4/V2/s2 [3]),
    .Z(\V1/V4/V2/A3/M2/s1 ));
 AND2_X1 \V1/V4/V2/A3/M2/M2/_0_  (.A1(\V1/V4/V2/A3/M2/s1 ),
    .A2(\V1/V4/V2/A3/c1 ),
    .ZN(\V1/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M2/M2/_1_  (.A(\V1/V4/V2/A3/M2/s1 ),
    .B(\V1/V4/V2/A3/c1 ),
    .Z(\V1/V4/v2 [5]));
 OR2_X1 \V1/V4/V2/A3/M2/_0_  (.A1(\V1/V4/V2/A3/M2/c1 ),
    .A2(\V1/V4/V2/A3/M2/c2 ),
    .ZN(\V1/V4/V2/A3/c2 ));
 AND2_X1 \V1/V4/V2/A3/M3/M1/_0_  (.A1(\V1/V4/V2/v4 [2]),
    .A2(\V1/V4/V2/c3 ),
    .ZN(\V1/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M3/M1/_1_  (.A(\V1/V4/V2/v4 [2]),
    .B(\V1/V4/V2/c3 ),
    .Z(\V1/V4/V2/A3/M3/s1 ));
 AND2_X1 \V1/V4/V2/A3/M3/M2/_0_  (.A1(\V1/V4/V2/A3/M3/s1 ),
    .A2(\V1/V4/V2/A3/c2 ),
    .ZN(\V1/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M3/M2/_1_  (.A(\V1/V4/V2/A3/M3/s1 ),
    .B(\V1/V4/V2/A3/c2 ),
    .Z(\V1/V4/v2 [6]));
 OR2_X1 \V1/V4/V2/A3/M3/_0_  (.A1(\V1/V4/V2/A3/M3/c1 ),
    .A2(\V1/V4/V2/A3/M3/c2 ),
    .ZN(\V1/V4/V2/A3/c3 ));
 AND2_X1 \V1/V4/V2/A3/M4/M1/_0_  (.A1(\V1/V4/V2/v4 [3]),
    .A2(ground),
    .ZN(\V1/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M4/M1/_1_  (.A(\V1/V4/V2/v4 [3]),
    .B(ground),
    .Z(\V1/V4/V2/A3/M4/s1 ));
 AND2_X1 \V1/V4/V2/A3/M4/M2/_0_  (.A1(\V1/V4/V2/A3/M4/s1 ),
    .A2(\V1/V4/V2/A3/c3 ),
    .ZN(\V1/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M4/M2/_1_  (.A(\V1/V4/V2/A3/M4/s1 ),
    .B(\V1/V4/V2/A3/c3 ),
    .Z(\V1/V4/v2 [7]));
 OR2_X1 \V1/V4/V2/A3/M4/_0_  (.A1(\V1/V4/V2/A3/M4/c1 ),
    .A2(\V1/V4/V2/A3/M4/c2 ),
    .ZN(\V1/V4/V2/overflow ));
 AND2_X1 \V1/V4/V2/V1/HA1/_0_  (.A1(\V1/V4/V2/V1/w2 ),
    .A2(\V1/V4/V2/V1/w1 ),
    .ZN(\V1/V4/V2/V1/w4 ));
 XOR2_X2 \V1/V4/V2/V1/HA1/_1_  (.A(\V1/V4/V2/V1/w2 ),
    .B(\V1/V4/V2/V1/w1 ),
    .Z(\V1/V4/v2 [1]));
 AND2_X1 \V1/V4/V2/V1/HA2/_0_  (.A1(\V1/V4/V2/V1/w4 ),
    .A2(\V1/V4/V2/V1/w3 ),
    .ZN(\V1/V4/V2/v1 [3]));
 XOR2_X2 \V1/V4/V2/V1/HA2/_1_  (.A(\V1/V4/V2/V1/w4 ),
    .B(\V1/V4/V2/V1/w3 ),
    .Z(\V1/V4/V2/v1 [2]));
 AND2_X1 \V1/V4/V2/V1/_0_  (.A1(A[12]),
    .A2(B[8]),
    .ZN(\V1/V4/v2 [0]));
 AND2_X1 \V1/V4/V2/V1/_1_  (.A1(A[12]),
    .A2(B[9]),
    .ZN(\V1/V4/V2/V1/w1 ));
 AND2_X1 \V1/V4/V2/V1/_2_  (.A1(B[8]),
    .A2(A[13]),
    .ZN(\V1/V4/V2/V1/w2 ));
 AND2_X1 \V1/V4/V2/V1/_3_  (.A1(B[9]),
    .A2(A[13]),
    .ZN(\V1/V4/V2/V1/w3 ));
 AND2_X1 \V1/V4/V2/V2/HA1/_0_  (.A1(\V1/V4/V2/V2/w2 ),
    .A2(\V1/V4/V2/V2/w1 ),
    .ZN(\V1/V4/V2/V2/w4 ));
 XOR2_X2 \V1/V4/V2/V2/HA1/_1_  (.A(\V1/V4/V2/V2/w2 ),
    .B(\V1/V4/V2/V2/w1 ),
    .Z(\V1/V4/V2/v2 [1]));
 AND2_X1 \V1/V4/V2/V2/HA2/_0_  (.A1(\V1/V4/V2/V2/w4 ),
    .A2(\V1/V4/V2/V2/w3 ),
    .ZN(\V1/V4/V2/v2 [3]));
 XOR2_X2 \V1/V4/V2/V2/HA2/_1_  (.A(\V1/V4/V2/V2/w4 ),
    .B(\V1/V4/V2/V2/w3 ),
    .Z(\V1/V4/V2/v2 [2]));
 AND2_X1 \V1/V4/V2/V2/_0_  (.A1(A[14]),
    .A2(B[8]),
    .ZN(\V1/V4/V2/v2 [0]));
 AND2_X1 \V1/V4/V2/V2/_1_  (.A1(A[14]),
    .A2(B[9]),
    .ZN(\V1/V4/V2/V2/w1 ));
 AND2_X1 \V1/V4/V2/V2/_2_  (.A1(B[8]),
    .A2(A[15]),
    .ZN(\V1/V4/V2/V2/w2 ));
 AND2_X1 \V1/V4/V2/V2/_3_  (.A1(B[9]),
    .A2(A[15]),
    .ZN(\V1/V4/V2/V2/w3 ));
 AND2_X1 \V1/V4/V2/V3/HA1/_0_  (.A1(\V1/V4/V2/V3/w2 ),
    .A2(\V1/V4/V2/V3/w1 ),
    .ZN(\V1/V4/V2/V3/w4 ));
 XOR2_X2 \V1/V4/V2/V3/HA1/_1_  (.A(\V1/V4/V2/V3/w2 ),
    .B(\V1/V4/V2/V3/w1 ),
    .Z(\V1/V4/V2/v3 [1]));
 AND2_X1 \V1/V4/V2/V3/HA2/_0_  (.A1(\V1/V4/V2/V3/w4 ),
    .A2(\V1/V4/V2/V3/w3 ),
    .ZN(\V1/V4/V2/v3 [3]));
 XOR2_X2 \V1/V4/V2/V3/HA2/_1_  (.A(\V1/V4/V2/V3/w4 ),
    .B(\V1/V4/V2/V3/w3 ),
    .Z(\V1/V4/V2/v3 [2]));
 AND2_X1 \V1/V4/V2/V3/_0_  (.A1(A[12]),
    .A2(B[10]),
    .ZN(\V1/V4/V2/v3 [0]));
 AND2_X1 \V1/V4/V2/V3/_1_  (.A1(A[12]),
    .A2(B[11]),
    .ZN(\V1/V4/V2/V3/w1 ));
 AND2_X1 \V1/V4/V2/V3/_2_  (.A1(B[10]),
    .A2(A[13]),
    .ZN(\V1/V4/V2/V3/w2 ));
 AND2_X1 \V1/V4/V2/V3/_3_  (.A1(B[11]),
    .A2(A[13]),
    .ZN(\V1/V4/V2/V3/w3 ));
 AND2_X1 \V1/V4/V2/V4/HA1/_0_  (.A1(\V1/V4/V2/V4/w2 ),
    .A2(\V1/V4/V2/V4/w1 ),
    .ZN(\V1/V4/V2/V4/w4 ));
 XOR2_X2 \V1/V4/V2/V4/HA1/_1_  (.A(\V1/V4/V2/V4/w2 ),
    .B(\V1/V4/V2/V4/w1 ),
    .Z(\V1/V4/V2/v4 [1]));
 AND2_X1 \V1/V4/V2/V4/HA2/_0_  (.A1(\V1/V4/V2/V4/w4 ),
    .A2(\V1/V4/V2/V4/w3 ),
    .ZN(\V1/V4/V2/v4 [3]));
 XOR2_X2 \V1/V4/V2/V4/HA2/_1_  (.A(\V1/V4/V2/V4/w4 ),
    .B(\V1/V4/V2/V4/w3 ),
    .Z(\V1/V4/V2/v4 [2]));
 AND2_X1 \V1/V4/V2/V4/_0_  (.A1(A[14]),
    .A2(B[10]),
    .ZN(\V1/V4/V2/v4 [0]));
 AND2_X1 \V1/V4/V2/V4/_1_  (.A1(A[14]),
    .A2(B[11]),
    .ZN(\V1/V4/V2/V4/w1 ));
 AND2_X1 \V1/V4/V2/V4/_2_  (.A1(B[10]),
    .A2(A[15]),
    .ZN(\V1/V4/V2/V4/w2 ));
 AND2_X1 \V1/V4/V2/V4/_3_  (.A1(B[11]),
    .A2(A[15]),
    .ZN(\V1/V4/V2/V4/w3 ));
 OR2_X1 \V1/V4/V2/_0_  (.A1(\V1/V4/V2/c1 ),
    .A2(\V1/V4/V2/c2 ),
    .ZN(\V1/V4/V2/c3 ));
 AND2_X1 \V1/V4/V3/A1/M1/M1/_0_  (.A1(\V1/V4/V3/v2 [0]),
    .A2(\V1/V4/V3/v3 [0]),
    .ZN(\V1/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M1/M1/_1_  (.A(\V1/V4/V3/v2 [0]),
    .B(\V1/V4/V3/v3 [0]),
    .Z(\V1/V4/V3/A1/M1/s1 ));
 AND2_X1 \V1/V4/V3/A1/M1/M2/_0_  (.A1(\V1/V4/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M1/M2/_1_  (.A(\V1/V4/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/V3/s1 [0]));
 OR2_X1 \V1/V4/V3/A1/M1/_0_  (.A1(\V1/V4/V3/A1/M1/c1 ),
    .A2(\V1/V4/V3/A1/M1/c2 ),
    .ZN(\V1/V4/V3/A1/c1 ));
 AND2_X1 \V1/V4/V3/A1/M2/M1/_0_  (.A1(\V1/V4/V3/v2 [1]),
    .A2(\V1/V4/V3/v3 [1]),
    .ZN(\V1/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M2/M1/_1_  (.A(\V1/V4/V3/v2 [1]),
    .B(\V1/V4/V3/v3 [1]),
    .Z(\V1/V4/V3/A1/M2/s1 ));
 AND2_X1 \V1/V4/V3/A1/M2/M2/_0_  (.A1(\V1/V4/V3/A1/M2/s1 ),
    .A2(\V1/V4/V3/A1/c1 ),
    .ZN(\V1/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M2/M2/_1_  (.A(\V1/V4/V3/A1/M2/s1 ),
    .B(\V1/V4/V3/A1/c1 ),
    .Z(\V1/V4/V3/s1 [1]));
 OR2_X1 \V1/V4/V3/A1/M2/_0_  (.A1(\V1/V4/V3/A1/M2/c1 ),
    .A2(\V1/V4/V3/A1/M2/c2 ),
    .ZN(\V1/V4/V3/A1/c2 ));
 AND2_X1 \V1/V4/V3/A1/M3/M1/_0_  (.A1(\V1/V4/V3/v2 [2]),
    .A2(\V1/V4/V3/v3 [2]),
    .ZN(\V1/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M3/M1/_1_  (.A(\V1/V4/V3/v2 [2]),
    .B(\V1/V4/V3/v3 [2]),
    .Z(\V1/V4/V3/A1/M3/s1 ));
 AND2_X1 \V1/V4/V3/A1/M3/M2/_0_  (.A1(\V1/V4/V3/A1/M3/s1 ),
    .A2(\V1/V4/V3/A1/c2 ),
    .ZN(\V1/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M3/M2/_1_  (.A(\V1/V4/V3/A1/M3/s1 ),
    .B(\V1/V4/V3/A1/c2 ),
    .Z(\V1/V4/V3/s1 [2]));
 OR2_X1 \V1/V4/V3/A1/M3/_0_  (.A1(\V1/V4/V3/A1/M3/c1 ),
    .A2(\V1/V4/V3/A1/M3/c2 ),
    .ZN(\V1/V4/V3/A1/c3 ));
 AND2_X1 \V1/V4/V3/A1/M4/M1/_0_  (.A1(\V1/V4/V3/v2 [3]),
    .A2(\V1/V4/V3/v3 [3]),
    .ZN(\V1/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M4/M1/_1_  (.A(\V1/V4/V3/v2 [3]),
    .B(\V1/V4/V3/v3 [3]),
    .Z(\V1/V4/V3/A1/M4/s1 ));
 AND2_X1 \V1/V4/V3/A1/M4/M2/_0_  (.A1(\V1/V4/V3/A1/M4/s1 ),
    .A2(\V1/V4/V3/A1/c3 ),
    .ZN(\V1/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M4/M2/_1_  (.A(\V1/V4/V3/A1/M4/s1 ),
    .B(\V1/V4/V3/A1/c3 ),
    .Z(\V1/V4/V3/s1 [3]));
 OR2_X1 \V1/V4/V3/A1/M4/_0_  (.A1(\V1/V4/V3/A1/M4/c1 ),
    .A2(\V1/V4/V3/A1/M4/c2 ),
    .ZN(\V1/V4/V3/c1 ));
 AND2_X1 \V1/V4/V3/A2/M1/M1/_0_  (.A1(\V1/V4/V3/s1 [0]),
    .A2(\V1/V4/V3/v1 [2]),
    .ZN(\V1/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M1/M1/_1_  (.A(\V1/V4/V3/s1 [0]),
    .B(\V1/V4/V3/v1 [2]),
    .Z(\V1/V4/V3/A2/M1/s1 ));
 AND2_X1 \V1/V4/V3/A2/M1/M2/_0_  (.A1(\V1/V4/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M1/M2/_1_  (.A(\V1/V4/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v3 [2]));
 OR2_X1 \V1/V4/V3/A2/M1/_0_  (.A1(\V1/V4/V3/A2/M1/c1 ),
    .A2(\V1/V4/V3/A2/M1/c2 ),
    .ZN(\V1/V4/V3/A2/c1 ));
 AND2_X1 \V1/V4/V3/A2/M2/M1/_0_  (.A1(\V1/V4/V3/s1 [1]),
    .A2(\V1/V4/V3/v1 [3]),
    .ZN(\V1/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M2/M1/_1_  (.A(\V1/V4/V3/s1 [1]),
    .B(\V1/V4/V3/v1 [3]),
    .Z(\V1/V4/V3/A2/M2/s1 ));
 AND2_X1 \V1/V4/V3/A2/M2/M2/_0_  (.A1(\V1/V4/V3/A2/M2/s1 ),
    .A2(\V1/V4/V3/A2/c1 ),
    .ZN(\V1/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M2/M2/_1_  (.A(\V1/V4/V3/A2/M2/s1 ),
    .B(\V1/V4/V3/A2/c1 ),
    .Z(\V1/V4/v3 [3]));
 OR2_X1 \V1/V4/V3/A2/M2/_0_  (.A1(\V1/V4/V3/A2/M2/c1 ),
    .A2(\V1/V4/V3/A2/M2/c2 ),
    .ZN(\V1/V4/V3/A2/c2 ));
 AND2_X1 \V1/V4/V3/A2/M3/M1/_0_  (.A1(\V1/V4/V3/s1 [2]),
    .A2(ground),
    .ZN(\V1/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M3/M1/_1_  (.A(\V1/V4/V3/s1 [2]),
    .B(ground),
    .Z(\V1/V4/V3/A2/M3/s1 ));
 AND2_X1 \V1/V4/V3/A2/M3/M2/_0_  (.A1(\V1/V4/V3/A2/M3/s1 ),
    .A2(\V1/V4/V3/A2/c2 ),
    .ZN(\V1/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M3/M2/_1_  (.A(\V1/V4/V3/A2/M3/s1 ),
    .B(\V1/V4/V3/A2/c2 ),
    .Z(\V1/V4/V3/s2 [2]));
 OR2_X1 \V1/V4/V3/A2/M3/_0_  (.A1(\V1/V4/V3/A2/M3/c1 ),
    .A2(\V1/V4/V3/A2/M3/c2 ),
    .ZN(\V1/V4/V3/A2/c3 ));
 AND2_X1 \V1/V4/V3/A2/M4/M1/_0_  (.A1(\V1/V4/V3/s1 [3]),
    .A2(ground),
    .ZN(\V1/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M4/M1/_1_  (.A(\V1/V4/V3/s1 [3]),
    .B(ground),
    .Z(\V1/V4/V3/A2/M4/s1 ));
 AND2_X1 \V1/V4/V3/A2/M4/M2/_0_  (.A1(\V1/V4/V3/A2/M4/s1 ),
    .A2(\V1/V4/V3/A2/c3 ),
    .ZN(\V1/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M4/M2/_1_  (.A(\V1/V4/V3/A2/M4/s1 ),
    .B(\V1/V4/V3/A2/c3 ),
    .Z(\V1/V4/V3/s2 [3]));
 OR2_X1 \V1/V4/V3/A2/M4/_0_  (.A1(\V1/V4/V3/A2/M4/c1 ),
    .A2(\V1/V4/V3/A2/M4/c2 ),
    .ZN(\V1/V4/V3/c2 ));
 AND2_X1 \V1/V4/V3/A3/M1/M1/_0_  (.A1(\V1/V4/V3/v4 [0]),
    .A2(\V1/V4/V3/s2 [2]),
    .ZN(\V1/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M1/M1/_1_  (.A(\V1/V4/V3/v4 [0]),
    .B(\V1/V4/V3/s2 [2]),
    .Z(\V1/V4/V3/A3/M1/s1 ));
 AND2_X1 \V1/V4/V3/A3/M1/M2/_0_  (.A1(\V1/V4/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M1/M2/_1_  (.A(\V1/V4/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v3 [4]));
 OR2_X1 \V1/V4/V3/A3/M1/_0_  (.A1(\V1/V4/V3/A3/M1/c1 ),
    .A2(\V1/V4/V3/A3/M1/c2 ),
    .ZN(\V1/V4/V3/A3/c1 ));
 AND2_X1 \V1/V4/V3/A3/M2/M1/_0_  (.A1(\V1/V4/V3/v4 [1]),
    .A2(\V1/V4/V3/s2 [3]),
    .ZN(\V1/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M2/M1/_1_  (.A(\V1/V4/V3/v4 [1]),
    .B(\V1/V4/V3/s2 [3]),
    .Z(\V1/V4/V3/A3/M2/s1 ));
 AND2_X1 \V1/V4/V3/A3/M2/M2/_0_  (.A1(\V1/V4/V3/A3/M2/s1 ),
    .A2(\V1/V4/V3/A3/c1 ),
    .ZN(\V1/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M2/M2/_1_  (.A(\V1/V4/V3/A3/M2/s1 ),
    .B(\V1/V4/V3/A3/c1 ),
    .Z(\V1/V4/v3 [5]));
 OR2_X1 \V1/V4/V3/A3/M2/_0_  (.A1(\V1/V4/V3/A3/M2/c1 ),
    .A2(\V1/V4/V3/A3/M2/c2 ),
    .ZN(\V1/V4/V3/A3/c2 ));
 AND2_X1 \V1/V4/V3/A3/M3/M1/_0_  (.A1(\V1/V4/V3/v4 [2]),
    .A2(\V1/V4/V3/c3 ),
    .ZN(\V1/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M3/M1/_1_  (.A(\V1/V4/V3/v4 [2]),
    .B(\V1/V4/V3/c3 ),
    .Z(\V1/V4/V3/A3/M3/s1 ));
 AND2_X1 \V1/V4/V3/A3/M3/M2/_0_  (.A1(\V1/V4/V3/A3/M3/s1 ),
    .A2(\V1/V4/V3/A3/c2 ),
    .ZN(\V1/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M3/M2/_1_  (.A(\V1/V4/V3/A3/M3/s1 ),
    .B(\V1/V4/V3/A3/c2 ),
    .Z(\V1/V4/v3 [6]));
 OR2_X1 \V1/V4/V3/A3/M3/_0_  (.A1(\V1/V4/V3/A3/M3/c1 ),
    .A2(\V1/V4/V3/A3/M3/c2 ),
    .ZN(\V1/V4/V3/A3/c3 ));
 AND2_X1 \V1/V4/V3/A3/M4/M1/_0_  (.A1(\V1/V4/V3/v4 [3]),
    .A2(ground),
    .ZN(\V1/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M4/M1/_1_  (.A(\V1/V4/V3/v4 [3]),
    .B(ground),
    .Z(\V1/V4/V3/A3/M4/s1 ));
 AND2_X1 \V1/V4/V3/A3/M4/M2/_0_  (.A1(\V1/V4/V3/A3/M4/s1 ),
    .A2(\V1/V4/V3/A3/c3 ),
    .ZN(\V1/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M4/M2/_1_  (.A(\V1/V4/V3/A3/M4/s1 ),
    .B(\V1/V4/V3/A3/c3 ),
    .Z(\V1/V4/v3 [7]));
 OR2_X1 \V1/V4/V3/A3/M4/_0_  (.A1(\V1/V4/V3/A3/M4/c1 ),
    .A2(\V1/V4/V3/A3/M4/c2 ),
    .ZN(\V1/V4/V3/overflow ));
 AND2_X1 \V1/V4/V3/V1/HA1/_0_  (.A1(\V1/V4/V3/V1/w2 ),
    .A2(\V1/V4/V3/V1/w1 ),
    .ZN(\V1/V4/V3/V1/w4 ));
 XOR2_X2 \V1/V4/V3/V1/HA1/_1_  (.A(\V1/V4/V3/V1/w2 ),
    .B(\V1/V4/V3/V1/w1 ),
    .Z(\V1/V4/v3 [1]));
 AND2_X1 \V1/V4/V3/V1/HA2/_0_  (.A1(\V1/V4/V3/V1/w4 ),
    .A2(\V1/V4/V3/V1/w3 ),
    .ZN(\V1/V4/V3/v1 [3]));
 XOR2_X2 \V1/V4/V3/V1/HA2/_1_  (.A(\V1/V4/V3/V1/w4 ),
    .B(\V1/V4/V3/V1/w3 ),
    .Z(\V1/V4/V3/v1 [2]));
 AND2_X1 \V1/V4/V3/V1/_0_  (.A1(A[8]),
    .A2(B[12]),
    .ZN(\V1/V4/v3 [0]));
 AND2_X1 \V1/V4/V3/V1/_1_  (.A1(A[8]),
    .A2(B[13]),
    .ZN(\V1/V4/V3/V1/w1 ));
 AND2_X1 \V1/V4/V3/V1/_2_  (.A1(B[12]),
    .A2(A[9]),
    .ZN(\V1/V4/V3/V1/w2 ));
 AND2_X1 \V1/V4/V3/V1/_3_  (.A1(B[13]),
    .A2(A[9]),
    .ZN(\V1/V4/V3/V1/w3 ));
 AND2_X1 \V1/V4/V3/V2/HA1/_0_  (.A1(\V1/V4/V3/V2/w2 ),
    .A2(\V1/V4/V3/V2/w1 ),
    .ZN(\V1/V4/V3/V2/w4 ));
 XOR2_X2 \V1/V4/V3/V2/HA1/_1_  (.A(\V1/V4/V3/V2/w2 ),
    .B(\V1/V4/V3/V2/w1 ),
    .Z(\V1/V4/V3/v2 [1]));
 AND2_X1 \V1/V4/V3/V2/HA2/_0_  (.A1(\V1/V4/V3/V2/w4 ),
    .A2(\V1/V4/V3/V2/w3 ),
    .ZN(\V1/V4/V3/v2 [3]));
 XOR2_X2 \V1/V4/V3/V2/HA2/_1_  (.A(\V1/V4/V3/V2/w4 ),
    .B(\V1/V4/V3/V2/w3 ),
    .Z(\V1/V4/V3/v2 [2]));
 AND2_X1 \V1/V4/V3/V2/_0_  (.A1(A[10]),
    .A2(B[12]),
    .ZN(\V1/V4/V3/v2 [0]));
 AND2_X1 \V1/V4/V3/V2/_1_  (.A1(A[10]),
    .A2(B[13]),
    .ZN(\V1/V4/V3/V2/w1 ));
 AND2_X1 \V1/V4/V3/V2/_2_  (.A1(B[12]),
    .A2(A[11]),
    .ZN(\V1/V4/V3/V2/w2 ));
 AND2_X1 \V1/V4/V3/V2/_3_  (.A1(B[13]),
    .A2(A[11]),
    .ZN(\V1/V4/V3/V2/w3 ));
 AND2_X1 \V1/V4/V3/V3/HA1/_0_  (.A1(\V1/V4/V3/V3/w2 ),
    .A2(\V1/V4/V3/V3/w1 ),
    .ZN(\V1/V4/V3/V3/w4 ));
 XOR2_X2 \V1/V4/V3/V3/HA1/_1_  (.A(\V1/V4/V3/V3/w2 ),
    .B(\V1/V4/V3/V3/w1 ),
    .Z(\V1/V4/V3/v3 [1]));
 AND2_X1 \V1/V4/V3/V3/HA2/_0_  (.A1(\V1/V4/V3/V3/w4 ),
    .A2(\V1/V4/V3/V3/w3 ),
    .ZN(\V1/V4/V3/v3 [3]));
 XOR2_X2 \V1/V4/V3/V3/HA2/_1_  (.A(\V1/V4/V3/V3/w4 ),
    .B(\V1/V4/V3/V3/w3 ),
    .Z(\V1/V4/V3/v3 [2]));
 AND2_X1 \V1/V4/V3/V3/_0_  (.A1(A[8]),
    .A2(B[14]),
    .ZN(\V1/V4/V3/v3 [0]));
 AND2_X1 \V1/V4/V3/V3/_1_  (.A1(A[8]),
    .A2(B[15]),
    .ZN(\V1/V4/V3/V3/w1 ));
 AND2_X1 \V1/V4/V3/V3/_2_  (.A1(B[14]),
    .A2(A[9]),
    .ZN(\V1/V4/V3/V3/w2 ));
 AND2_X1 \V1/V4/V3/V3/_3_  (.A1(B[15]),
    .A2(A[9]),
    .ZN(\V1/V4/V3/V3/w3 ));
 AND2_X1 \V1/V4/V3/V4/HA1/_0_  (.A1(\V1/V4/V3/V4/w2 ),
    .A2(\V1/V4/V3/V4/w1 ),
    .ZN(\V1/V4/V3/V4/w4 ));
 XOR2_X2 \V1/V4/V3/V4/HA1/_1_  (.A(\V1/V4/V3/V4/w2 ),
    .B(\V1/V4/V3/V4/w1 ),
    .Z(\V1/V4/V3/v4 [1]));
 AND2_X1 \V1/V4/V3/V4/HA2/_0_  (.A1(\V1/V4/V3/V4/w4 ),
    .A2(\V1/V4/V3/V4/w3 ),
    .ZN(\V1/V4/V3/v4 [3]));
 XOR2_X2 \V1/V4/V3/V4/HA2/_1_  (.A(\V1/V4/V3/V4/w4 ),
    .B(\V1/V4/V3/V4/w3 ),
    .Z(\V1/V4/V3/v4 [2]));
 AND2_X1 \V1/V4/V3/V4/_0_  (.A1(A[10]),
    .A2(B[14]),
    .ZN(\V1/V4/V3/v4 [0]));
 AND2_X1 \V1/V4/V3/V4/_1_  (.A1(A[10]),
    .A2(B[15]),
    .ZN(\V1/V4/V3/V4/w1 ));
 AND2_X1 \V1/V4/V3/V4/_2_  (.A1(B[14]),
    .A2(A[11]),
    .ZN(\V1/V4/V3/V4/w2 ));
 AND2_X1 \V1/V4/V3/V4/_3_  (.A1(B[15]),
    .A2(A[11]),
    .ZN(\V1/V4/V3/V4/w3 ));
 OR2_X1 \V1/V4/V3/_0_  (.A1(\V1/V4/V3/c1 ),
    .A2(\V1/V4/V3/c2 ),
    .ZN(\V1/V4/V3/c3 ));
 AND2_X1 \V1/V4/V4/A1/M1/M1/_0_  (.A1(\V1/V4/V4/v2 [0]),
    .A2(\V1/V4/V4/v3 [0]),
    .ZN(\V1/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M1/M1/_1_  (.A(\V1/V4/V4/v2 [0]),
    .B(\V1/V4/V4/v3 [0]),
    .Z(\V1/V4/V4/A1/M1/s1 ));
 AND2_X1 \V1/V4/V4/A1/M1/M2/_0_  (.A1(\V1/V4/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M1/M2/_1_  (.A(\V1/V4/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/V4/s1 [0]));
 OR2_X1 \V1/V4/V4/A1/M1/_0_  (.A1(\V1/V4/V4/A1/M1/c1 ),
    .A2(\V1/V4/V4/A1/M1/c2 ),
    .ZN(\V1/V4/V4/A1/c1 ));
 AND2_X1 \V1/V4/V4/A1/M2/M1/_0_  (.A1(\V1/V4/V4/v2 [1]),
    .A2(\V1/V4/V4/v3 [1]),
    .ZN(\V1/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M2/M1/_1_  (.A(\V1/V4/V4/v2 [1]),
    .B(\V1/V4/V4/v3 [1]),
    .Z(\V1/V4/V4/A1/M2/s1 ));
 AND2_X1 \V1/V4/V4/A1/M2/M2/_0_  (.A1(\V1/V4/V4/A1/M2/s1 ),
    .A2(\V1/V4/V4/A1/c1 ),
    .ZN(\V1/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M2/M2/_1_  (.A(\V1/V4/V4/A1/M2/s1 ),
    .B(\V1/V4/V4/A1/c1 ),
    .Z(\V1/V4/V4/s1 [1]));
 OR2_X1 \V1/V4/V4/A1/M2/_0_  (.A1(\V1/V4/V4/A1/M2/c1 ),
    .A2(\V1/V4/V4/A1/M2/c2 ),
    .ZN(\V1/V4/V4/A1/c2 ));
 AND2_X1 \V1/V4/V4/A1/M3/M1/_0_  (.A1(\V1/V4/V4/v2 [2]),
    .A2(\V1/V4/V4/v3 [2]),
    .ZN(\V1/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M3/M1/_1_  (.A(\V1/V4/V4/v2 [2]),
    .B(\V1/V4/V4/v3 [2]),
    .Z(\V1/V4/V4/A1/M3/s1 ));
 AND2_X1 \V1/V4/V4/A1/M3/M2/_0_  (.A1(\V1/V4/V4/A1/M3/s1 ),
    .A2(\V1/V4/V4/A1/c2 ),
    .ZN(\V1/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M3/M2/_1_  (.A(\V1/V4/V4/A1/M3/s1 ),
    .B(\V1/V4/V4/A1/c2 ),
    .Z(\V1/V4/V4/s1 [2]));
 OR2_X1 \V1/V4/V4/A1/M3/_0_  (.A1(\V1/V4/V4/A1/M3/c1 ),
    .A2(\V1/V4/V4/A1/M3/c2 ),
    .ZN(\V1/V4/V4/A1/c3 ));
 AND2_X1 \V1/V4/V4/A1/M4/M1/_0_  (.A1(\V1/V4/V4/v2 [3]),
    .A2(\V1/V4/V4/v3 [3]),
    .ZN(\V1/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M4/M1/_1_  (.A(\V1/V4/V4/v2 [3]),
    .B(\V1/V4/V4/v3 [3]),
    .Z(\V1/V4/V4/A1/M4/s1 ));
 AND2_X1 \V1/V4/V4/A1/M4/M2/_0_  (.A1(\V1/V4/V4/A1/M4/s1 ),
    .A2(\V1/V4/V4/A1/c3 ),
    .ZN(\V1/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M4/M2/_1_  (.A(\V1/V4/V4/A1/M4/s1 ),
    .B(\V1/V4/V4/A1/c3 ),
    .Z(\V1/V4/V4/s1 [3]));
 OR2_X1 \V1/V4/V4/A1/M4/_0_  (.A1(\V1/V4/V4/A1/M4/c1 ),
    .A2(\V1/V4/V4/A1/M4/c2 ),
    .ZN(\V1/V4/V4/c1 ));
 AND2_X1 \V1/V4/V4/A2/M1/M1/_0_  (.A1(\V1/V4/V4/s1 [0]),
    .A2(\V1/V4/V4/v1 [2]),
    .ZN(\V1/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M1/M1/_1_  (.A(\V1/V4/V4/s1 [0]),
    .B(\V1/V4/V4/v1 [2]),
    .Z(\V1/V4/V4/A2/M1/s1 ));
 AND2_X1 \V1/V4/V4/A2/M1/M2/_0_  (.A1(\V1/V4/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M1/M2/_1_  (.A(\V1/V4/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v4 [2]));
 OR2_X1 \V1/V4/V4/A2/M1/_0_  (.A1(\V1/V4/V4/A2/M1/c1 ),
    .A2(\V1/V4/V4/A2/M1/c2 ),
    .ZN(\V1/V4/V4/A2/c1 ));
 AND2_X1 \V1/V4/V4/A2/M2/M1/_0_  (.A1(\V1/V4/V4/s1 [1]),
    .A2(\V1/V4/V4/v1 [3]),
    .ZN(\V1/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M2/M1/_1_  (.A(\V1/V4/V4/s1 [1]),
    .B(\V1/V4/V4/v1 [3]),
    .Z(\V1/V4/V4/A2/M2/s1 ));
 AND2_X1 \V1/V4/V4/A2/M2/M2/_0_  (.A1(\V1/V4/V4/A2/M2/s1 ),
    .A2(\V1/V4/V4/A2/c1 ),
    .ZN(\V1/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M2/M2/_1_  (.A(\V1/V4/V4/A2/M2/s1 ),
    .B(\V1/V4/V4/A2/c1 ),
    .Z(\V1/V4/v4 [3]));
 OR2_X1 \V1/V4/V4/A2/M2/_0_  (.A1(\V1/V4/V4/A2/M2/c1 ),
    .A2(\V1/V4/V4/A2/M2/c2 ),
    .ZN(\V1/V4/V4/A2/c2 ));
 AND2_X1 \V1/V4/V4/A2/M3/M1/_0_  (.A1(\V1/V4/V4/s1 [2]),
    .A2(ground),
    .ZN(\V1/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M3/M1/_1_  (.A(\V1/V4/V4/s1 [2]),
    .B(ground),
    .Z(\V1/V4/V4/A2/M3/s1 ));
 AND2_X1 \V1/V4/V4/A2/M3/M2/_0_  (.A1(\V1/V4/V4/A2/M3/s1 ),
    .A2(\V1/V4/V4/A2/c2 ),
    .ZN(\V1/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M3/M2/_1_  (.A(\V1/V4/V4/A2/M3/s1 ),
    .B(\V1/V4/V4/A2/c2 ),
    .Z(\V1/V4/V4/s2 [2]));
 OR2_X1 \V1/V4/V4/A2/M3/_0_  (.A1(\V1/V4/V4/A2/M3/c1 ),
    .A2(\V1/V4/V4/A2/M3/c2 ),
    .ZN(\V1/V4/V4/A2/c3 ));
 AND2_X1 \V1/V4/V4/A2/M4/M1/_0_  (.A1(\V1/V4/V4/s1 [3]),
    .A2(ground),
    .ZN(\V1/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M4/M1/_1_  (.A(\V1/V4/V4/s1 [3]),
    .B(ground),
    .Z(\V1/V4/V4/A2/M4/s1 ));
 AND2_X1 \V1/V4/V4/A2/M4/M2/_0_  (.A1(\V1/V4/V4/A2/M4/s1 ),
    .A2(\V1/V4/V4/A2/c3 ),
    .ZN(\V1/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M4/M2/_1_  (.A(\V1/V4/V4/A2/M4/s1 ),
    .B(\V1/V4/V4/A2/c3 ),
    .Z(\V1/V4/V4/s2 [3]));
 OR2_X1 \V1/V4/V4/A2/M4/_0_  (.A1(\V1/V4/V4/A2/M4/c1 ),
    .A2(\V1/V4/V4/A2/M4/c2 ),
    .ZN(\V1/V4/V4/c2 ));
 AND2_X1 \V1/V4/V4/A3/M1/M1/_0_  (.A1(\V1/V4/V4/v4 [0]),
    .A2(\V1/V4/V4/s2 [2]),
    .ZN(\V1/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M1/M1/_1_  (.A(\V1/V4/V4/v4 [0]),
    .B(\V1/V4/V4/s2 [2]),
    .Z(\V1/V4/V4/A3/M1/s1 ));
 AND2_X1 \V1/V4/V4/A3/M1/M2/_0_  (.A1(\V1/V4/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V1/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M1/M2/_1_  (.A(\V1/V4/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V1/V4/v4 [4]));
 OR2_X1 \V1/V4/V4/A3/M1/_0_  (.A1(\V1/V4/V4/A3/M1/c1 ),
    .A2(\V1/V4/V4/A3/M1/c2 ),
    .ZN(\V1/V4/V4/A3/c1 ));
 AND2_X1 \V1/V4/V4/A3/M2/M1/_0_  (.A1(\V1/V4/V4/v4 [1]),
    .A2(\V1/V4/V4/s2 [3]),
    .ZN(\V1/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M2/M1/_1_  (.A(\V1/V4/V4/v4 [1]),
    .B(\V1/V4/V4/s2 [3]),
    .Z(\V1/V4/V4/A3/M2/s1 ));
 AND2_X1 \V1/V4/V4/A3/M2/M2/_0_  (.A1(\V1/V4/V4/A3/M2/s1 ),
    .A2(\V1/V4/V4/A3/c1 ),
    .ZN(\V1/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M2/M2/_1_  (.A(\V1/V4/V4/A3/M2/s1 ),
    .B(\V1/V4/V4/A3/c1 ),
    .Z(\V1/V4/v4 [5]));
 OR2_X1 \V1/V4/V4/A3/M2/_0_  (.A1(\V1/V4/V4/A3/M2/c1 ),
    .A2(\V1/V4/V4/A3/M2/c2 ),
    .ZN(\V1/V4/V4/A3/c2 ));
 AND2_X1 \V1/V4/V4/A3/M3/M1/_0_  (.A1(\V1/V4/V4/v4 [2]),
    .A2(\V1/V4/V4/c3 ),
    .ZN(\V1/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M3/M1/_1_  (.A(\V1/V4/V4/v4 [2]),
    .B(\V1/V4/V4/c3 ),
    .Z(\V1/V4/V4/A3/M3/s1 ));
 AND2_X1 \V1/V4/V4/A3/M3/M2/_0_  (.A1(\V1/V4/V4/A3/M3/s1 ),
    .A2(\V1/V4/V4/A3/c2 ),
    .ZN(\V1/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M3/M2/_1_  (.A(\V1/V4/V4/A3/M3/s1 ),
    .B(\V1/V4/V4/A3/c2 ),
    .Z(\V1/V4/v4 [6]));
 OR2_X1 \V1/V4/V4/A3/M3/_0_  (.A1(\V1/V4/V4/A3/M3/c1 ),
    .A2(\V1/V4/V4/A3/M3/c2 ),
    .ZN(\V1/V4/V4/A3/c3 ));
 AND2_X1 \V1/V4/V4/A3/M4/M1/_0_  (.A1(\V1/V4/V4/v4 [3]),
    .A2(ground),
    .ZN(\V1/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M4/M1/_1_  (.A(\V1/V4/V4/v4 [3]),
    .B(ground),
    .Z(\V1/V4/V4/A3/M4/s1 ));
 AND2_X1 \V1/V4/V4/A3/M4/M2/_0_  (.A1(\V1/V4/V4/A3/M4/s1 ),
    .A2(\V1/V4/V4/A3/c3 ),
    .ZN(\V1/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M4/M2/_1_  (.A(\V1/V4/V4/A3/M4/s1 ),
    .B(\V1/V4/V4/A3/c3 ),
    .Z(\V1/V4/v4 [7]));
 OR2_X1 \V1/V4/V4/A3/M4/_0_  (.A1(\V1/V4/V4/A3/M4/c1 ),
    .A2(\V1/V4/V4/A3/M4/c2 ),
    .ZN(\V1/V4/V4/overflow ));
 AND2_X1 \V1/V4/V4/V1/HA1/_0_  (.A1(\V1/V4/V4/V1/w2 ),
    .A2(\V1/V4/V4/V1/w1 ),
    .ZN(\V1/V4/V4/V1/w4 ));
 XOR2_X2 \V1/V4/V4/V1/HA1/_1_  (.A(\V1/V4/V4/V1/w2 ),
    .B(\V1/V4/V4/V1/w1 ),
    .Z(\V1/V4/v4 [1]));
 AND2_X1 \V1/V4/V4/V1/HA2/_0_  (.A1(\V1/V4/V4/V1/w4 ),
    .A2(\V1/V4/V4/V1/w3 ),
    .ZN(\V1/V4/V4/v1 [3]));
 XOR2_X2 \V1/V4/V4/V1/HA2/_1_  (.A(\V1/V4/V4/V1/w4 ),
    .B(\V1/V4/V4/V1/w3 ),
    .Z(\V1/V4/V4/v1 [2]));
 AND2_X1 \V1/V4/V4/V1/_0_  (.A1(A[12]),
    .A2(B[12]),
    .ZN(\V1/V4/v4 [0]));
 AND2_X1 \V1/V4/V4/V1/_1_  (.A1(A[12]),
    .A2(B[13]),
    .ZN(\V1/V4/V4/V1/w1 ));
 AND2_X1 \V1/V4/V4/V1/_2_  (.A1(B[12]),
    .A2(A[13]),
    .ZN(\V1/V4/V4/V1/w2 ));
 AND2_X1 \V1/V4/V4/V1/_3_  (.A1(B[13]),
    .A2(A[13]),
    .ZN(\V1/V4/V4/V1/w3 ));
 AND2_X1 \V1/V4/V4/V2/HA1/_0_  (.A1(\V1/V4/V4/V2/w2 ),
    .A2(\V1/V4/V4/V2/w1 ),
    .ZN(\V1/V4/V4/V2/w4 ));
 XOR2_X2 \V1/V4/V4/V2/HA1/_1_  (.A(\V1/V4/V4/V2/w2 ),
    .B(\V1/V4/V4/V2/w1 ),
    .Z(\V1/V4/V4/v2 [1]));
 AND2_X1 \V1/V4/V4/V2/HA2/_0_  (.A1(\V1/V4/V4/V2/w4 ),
    .A2(\V1/V4/V4/V2/w3 ),
    .ZN(\V1/V4/V4/v2 [3]));
 XOR2_X2 \V1/V4/V4/V2/HA2/_1_  (.A(\V1/V4/V4/V2/w4 ),
    .B(\V1/V4/V4/V2/w3 ),
    .Z(\V1/V4/V4/v2 [2]));
 AND2_X1 \V1/V4/V4/V2/_0_  (.A1(A[14]),
    .A2(B[12]),
    .ZN(\V1/V4/V4/v2 [0]));
 AND2_X1 \V1/V4/V4/V2/_1_  (.A1(A[14]),
    .A2(B[13]),
    .ZN(\V1/V4/V4/V2/w1 ));
 AND2_X1 \V1/V4/V4/V2/_2_  (.A1(B[12]),
    .A2(A[15]),
    .ZN(\V1/V4/V4/V2/w2 ));
 AND2_X1 \V1/V4/V4/V2/_3_  (.A1(B[13]),
    .A2(A[15]),
    .ZN(\V1/V4/V4/V2/w3 ));
 AND2_X1 \V1/V4/V4/V3/HA1/_0_  (.A1(\V1/V4/V4/V3/w2 ),
    .A2(\V1/V4/V4/V3/w1 ),
    .ZN(\V1/V4/V4/V3/w4 ));
 XOR2_X2 \V1/V4/V4/V3/HA1/_1_  (.A(\V1/V4/V4/V3/w2 ),
    .B(\V1/V4/V4/V3/w1 ),
    .Z(\V1/V4/V4/v3 [1]));
 AND2_X1 \V1/V4/V4/V3/HA2/_0_  (.A1(\V1/V4/V4/V3/w4 ),
    .A2(\V1/V4/V4/V3/w3 ),
    .ZN(\V1/V4/V4/v3 [3]));
 XOR2_X2 \V1/V4/V4/V3/HA2/_1_  (.A(\V1/V4/V4/V3/w4 ),
    .B(\V1/V4/V4/V3/w3 ),
    .Z(\V1/V4/V4/v3 [2]));
 AND2_X1 \V1/V4/V4/V3/_0_  (.A1(A[12]),
    .A2(B[14]),
    .ZN(\V1/V4/V4/v3 [0]));
 AND2_X1 \V1/V4/V4/V3/_1_  (.A1(A[12]),
    .A2(B[15]),
    .ZN(\V1/V4/V4/V3/w1 ));
 AND2_X1 \V1/V4/V4/V3/_2_  (.A1(B[14]),
    .A2(A[13]),
    .ZN(\V1/V4/V4/V3/w2 ));
 AND2_X1 \V1/V4/V4/V3/_3_  (.A1(B[15]),
    .A2(A[13]),
    .ZN(\V1/V4/V4/V3/w3 ));
 AND2_X1 \V1/V4/V4/V4/HA1/_0_  (.A1(\V1/V4/V4/V4/w2 ),
    .A2(\V1/V4/V4/V4/w1 ),
    .ZN(\V1/V4/V4/V4/w4 ));
 XOR2_X2 \V1/V4/V4/V4/HA1/_1_  (.A(\V1/V4/V4/V4/w2 ),
    .B(\V1/V4/V4/V4/w1 ),
    .Z(\V1/V4/V4/v4 [1]));
 AND2_X1 \V1/V4/V4/V4/HA2/_0_  (.A1(\V1/V4/V4/V4/w4 ),
    .A2(\V1/V4/V4/V4/w3 ),
    .ZN(\V1/V4/V4/v4 [3]));
 XOR2_X2 \V1/V4/V4/V4/HA2/_1_  (.A(\V1/V4/V4/V4/w4 ),
    .B(\V1/V4/V4/V4/w3 ),
    .Z(\V1/V4/V4/v4 [2]));
 AND2_X1 \V1/V4/V4/V4/_0_  (.A1(A[14]),
    .A2(B[14]),
    .ZN(\V1/V4/V4/v4 [0]));
 AND2_X1 \V1/V4/V4/V4/_1_  (.A1(A[14]),
    .A2(B[15]),
    .ZN(\V1/V4/V4/V4/w1 ));
 AND2_X1 \V1/V4/V4/V4/_2_  (.A1(B[14]),
    .A2(A[15]),
    .ZN(\V1/V4/V4/V4/w2 ));
 AND2_X1 \V1/V4/V4/V4/_3_  (.A1(B[15]),
    .A2(A[15]),
    .ZN(\V1/V4/V4/V4/w3 ));
 OR2_X1 \V1/V4/V4/_0_  (.A1(\V1/V4/V4/c1 ),
    .A2(\V1/V4/V4/c2 ),
    .ZN(\V1/V4/V4/c3 ));
 OR2_X1 \V1/V4/_0_  (.A1(\V1/V4/c1 ),
    .A2(\V1/V4/c2 ),
    .ZN(\V1/V4/c3 ));
 OR2_X1 \V1/_0_  (.A1(\V1/c1 ),
    .A2(\V1/c2 ),
    .ZN(\V1/c3 ));
 AND2_X1 \V2/A1/A1/A1/M1/M1/_0_  (.A1(\V2/v2 [0]),
    .A2(\V2/v3 [0]),
    .ZN(\V2/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M1/M1/_1_  (.A(\V2/v2 [0]),
    .B(\V2/v3 [0]),
    .Z(\V2/A1/A1/A1/M1/s1 ));
 AND2_X1 \V2/A1/A1/A1/M1/M2/_0_  (.A1(\V2/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M1/M2/_1_  (.A(\V2/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/s1 [0]));
 OR2_X1 \V2/A1/A1/A1/M1/_0_  (.A1(\V2/A1/A1/A1/M1/c1 ),
    .A2(\V2/A1/A1/A1/M1/c2 ),
    .ZN(\V2/A1/A1/A1/c1 ));
 AND2_X1 \V2/A1/A1/A1/M2/M1/_0_  (.A1(\V2/v2 [1]),
    .A2(\V2/v3 [1]),
    .ZN(\V2/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M2/M1/_1_  (.A(\V2/v2 [1]),
    .B(\V2/v3 [1]),
    .Z(\V2/A1/A1/A1/M2/s1 ));
 AND2_X1 \V2/A1/A1/A1/M2/M2/_0_  (.A1(\V2/A1/A1/A1/M2/s1 ),
    .A2(\V2/A1/A1/A1/c1 ),
    .ZN(\V2/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M2/M2/_1_  (.A(\V2/A1/A1/A1/M2/s1 ),
    .B(\V2/A1/A1/A1/c1 ),
    .Z(\V2/s1 [1]));
 OR2_X1 \V2/A1/A1/A1/M2/_0_  (.A1(\V2/A1/A1/A1/M2/c1 ),
    .A2(\V2/A1/A1/A1/M2/c2 ),
    .ZN(\V2/A1/A1/A1/c2 ));
 AND2_X1 \V2/A1/A1/A1/M3/M1/_0_  (.A1(\V2/v2 [2]),
    .A2(\V2/v3 [2]),
    .ZN(\V2/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M3/M1/_1_  (.A(\V2/v2 [2]),
    .B(\V2/v3 [2]),
    .Z(\V2/A1/A1/A1/M3/s1 ));
 AND2_X1 \V2/A1/A1/A1/M3/M2/_0_  (.A1(\V2/A1/A1/A1/M3/s1 ),
    .A2(\V2/A1/A1/A1/c2 ),
    .ZN(\V2/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M3/M2/_1_  (.A(\V2/A1/A1/A1/M3/s1 ),
    .B(\V2/A1/A1/A1/c2 ),
    .Z(\V2/s1 [2]));
 OR2_X1 \V2/A1/A1/A1/M3/_0_  (.A1(\V2/A1/A1/A1/M3/c1 ),
    .A2(\V2/A1/A1/A1/M3/c2 ),
    .ZN(\V2/A1/A1/A1/c3 ));
 AND2_X1 \V2/A1/A1/A1/M4/M1/_0_  (.A1(\V2/v2 [3]),
    .A2(\V2/v3 [3]),
    .ZN(\V2/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M4/M1/_1_  (.A(\V2/v2 [3]),
    .B(\V2/v3 [3]),
    .Z(\V2/A1/A1/A1/M4/s1 ));
 AND2_X1 \V2/A1/A1/A1/M4/M2/_0_  (.A1(\V2/A1/A1/A1/M4/s1 ),
    .A2(\V2/A1/A1/A1/c3 ),
    .ZN(\V2/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M4/M2/_1_  (.A(\V2/A1/A1/A1/M4/s1 ),
    .B(\V2/A1/A1/A1/c3 ),
    .Z(\V2/s1 [3]));
 OR2_X1 \V2/A1/A1/A1/M4/_0_  (.A1(\V2/A1/A1/A1/M4/c1 ),
    .A2(\V2/A1/A1/A1/M4/c2 ),
    .ZN(\V2/A1/A1/c1 ));
 AND2_X1 \V2/A1/A1/A2/M1/M1/_0_  (.A1(\V2/v2 [4]),
    .A2(\V2/v3 [4]),
    .ZN(\V2/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M1/M1/_1_  (.A(\V2/v2 [4]),
    .B(\V2/v3 [4]),
    .Z(\V2/A1/A1/A2/M1/s1 ));
 AND2_X1 \V2/A1/A1/A2/M1/M2/_0_  (.A1(\V2/A1/A1/A2/M1/s1 ),
    .A2(\V2/A1/A1/c1 ),
    .ZN(\V2/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M1/M2/_1_  (.A(\V2/A1/A1/A2/M1/s1 ),
    .B(\V2/A1/A1/c1 ),
    .Z(\V2/s1 [4]));
 OR2_X1 \V2/A1/A1/A2/M1/_0_  (.A1(\V2/A1/A1/A2/M1/c1 ),
    .A2(\V2/A1/A1/A2/M1/c2 ),
    .ZN(\V2/A1/A1/A2/c1 ));
 AND2_X1 \V2/A1/A1/A2/M2/M1/_0_  (.A1(\V2/v2 [5]),
    .A2(\V2/v3 [5]),
    .ZN(\V2/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M2/M1/_1_  (.A(\V2/v2 [5]),
    .B(\V2/v3 [5]),
    .Z(\V2/A1/A1/A2/M2/s1 ));
 AND2_X1 \V2/A1/A1/A2/M2/M2/_0_  (.A1(\V2/A1/A1/A2/M2/s1 ),
    .A2(\V2/A1/A1/A2/c1 ),
    .ZN(\V2/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M2/M2/_1_  (.A(\V2/A1/A1/A2/M2/s1 ),
    .B(\V2/A1/A1/A2/c1 ),
    .Z(\V2/s1 [5]));
 OR2_X1 \V2/A1/A1/A2/M2/_0_  (.A1(\V2/A1/A1/A2/M2/c1 ),
    .A2(\V2/A1/A1/A2/M2/c2 ),
    .ZN(\V2/A1/A1/A2/c2 ));
 AND2_X1 \V2/A1/A1/A2/M3/M1/_0_  (.A1(\V2/v2 [6]),
    .A2(\V2/v3 [6]),
    .ZN(\V2/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M3/M1/_1_  (.A(\V2/v2 [6]),
    .B(\V2/v3 [6]),
    .Z(\V2/A1/A1/A2/M3/s1 ));
 AND2_X1 \V2/A1/A1/A2/M3/M2/_0_  (.A1(\V2/A1/A1/A2/M3/s1 ),
    .A2(\V2/A1/A1/A2/c2 ),
    .ZN(\V2/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M3/M2/_1_  (.A(\V2/A1/A1/A2/M3/s1 ),
    .B(\V2/A1/A1/A2/c2 ),
    .Z(\V2/s1 [6]));
 OR2_X1 \V2/A1/A1/A2/M3/_0_  (.A1(\V2/A1/A1/A2/M3/c1 ),
    .A2(\V2/A1/A1/A2/M3/c2 ),
    .ZN(\V2/A1/A1/A2/c3 ));
 AND2_X1 \V2/A1/A1/A2/M4/M1/_0_  (.A1(\V2/v2 [7]),
    .A2(\V2/v3 [7]),
    .ZN(\V2/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M4/M1/_1_  (.A(\V2/v2 [7]),
    .B(\V2/v3 [7]),
    .Z(\V2/A1/A1/A2/M4/s1 ));
 AND2_X1 \V2/A1/A1/A2/M4/M2/_0_  (.A1(\V2/A1/A1/A2/M4/s1 ),
    .A2(\V2/A1/A1/A2/c3 ),
    .ZN(\V2/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M4/M2/_1_  (.A(\V2/A1/A1/A2/M4/s1 ),
    .B(\V2/A1/A1/A2/c3 ),
    .Z(\V2/s1 [7]));
 OR2_X1 \V2/A1/A1/A2/M4/_0_  (.A1(\V2/A1/A1/A2/M4/c1 ),
    .A2(\V2/A1/A1/A2/M4/c2 ),
    .ZN(\V2/A1/c1 ));
 AND2_X1 \V2/A1/A2/A1/M1/M1/_0_  (.A1(\V2/v2 [8]),
    .A2(\V2/v3 [8]),
    .ZN(\V2/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M1/M1/_1_  (.A(\V2/v2 [8]),
    .B(\V2/v3 [8]),
    .Z(\V2/A1/A2/A1/M1/s1 ));
 AND2_X1 \V2/A1/A2/A1/M1/M2/_0_  (.A1(\V2/A1/A2/A1/M1/s1 ),
    .A2(\V2/A1/c1 ),
    .ZN(\V2/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M1/M2/_1_  (.A(\V2/A1/A2/A1/M1/s1 ),
    .B(\V2/A1/c1 ),
    .Z(\V2/s1 [8]));
 OR2_X1 \V2/A1/A2/A1/M1/_0_  (.A1(\V2/A1/A2/A1/M1/c1 ),
    .A2(\V2/A1/A2/A1/M1/c2 ),
    .ZN(\V2/A1/A2/A1/c1 ));
 AND2_X1 \V2/A1/A2/A1/M2/M1/_0_  (.A1(\V2/v2 [9]),
    .A2(\V2/v3 [9]),
    .ZN(\V2/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M2/M1/_1_  (.A(\V2/v2 [9]),
    .B(\V2/v3 [9]),
    .Z(\V2/A1/A2/A1/M2/s1 ));
 AND2_X1 \V2/A1/A2/A1/M2/M2/_0_  (.A1(\V2/A1/A2/A1/M2/s1 ),
    .A2(\V2/A1/A2/A1/c1 ),
    .ZN(\V2/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M2/M2/_1_  (.A(\V2/A1/A2/A1/M2/s1 ),
    .B(\V2/A1/A2/A1/c1 ),
    .Z(\V2/s1 [9]));
 OR2_X1 \V2/A1/A2/A1/M2/_0_  (.A1(\V2/A1/A2/A1/M2/c1 ),
    .A2(\V2/A1/A2/A1/M2/c2 ),
    .ZN(\V2/A1/A2/A1/c2 ));
 AND2_X1 \V2/A1/A2/A1/M3/M1/_0_  (.A1(\V2/v2 [10]),
    .A2(\V2/v3 [10]),
    .ZN(\V2/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M3/M1/_1_  (.A(\V2/v2 [10]),
    .B(\V2/v3 [10]),
    .Z(\V2/A1/A2/A1/M3/s1 ));
 AND2_X1 \V2/A1/A2/A1/M3/M2/_0_  (.A1(\V2/A1/A2/A1/M3/s1 ),
    .A2(\V2/A1/A2/A1/c2 ),
    .ZN(\V2/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M3/M2/_1_  (.A(\V2/A1/A2/A1/M3/s1 ),
    .B(\V2/A1/A2/A1/c2 ),
    .Z(\V2/s1 [10]));
 OR2_X1 \V2/A1/A2/A1/M3/_0_  (.A1(\V2/A1/A2/A1/M3/c1 ),
    .A2(\V2/A1/A2/A1/M3/c2 ),
    .ZN(\V2/A1/A2/A1/c3 ));
 AND2_X1 \V2/A1/A2/A1/M4/M1/_0_  (.A1(\V2/v2 [11]),
    .A2(\V2/v3 [11]),
    .ZN(\V2/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M4/M1/_1_  (.A(\V2/v2 [11]),
    .B(\V2/v3 [11]),
    .Z(\V2/A1/A2/A1/M4/s1 ));
 AND2_X1 \V2/A1/A2/A1/M4/M2/_0_  (.A1(\V2/A1/A2/A1/M4/s1 ),
    .A2(\V2/A1/A2/A1/c3 ),
    .ZN(\V2/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M4/M2/_1_  (.A(\V2/A1/A2/A1/M4/s1 ),
    .B(\V2/A1/A2/A1/c3 ),
    .Z(\V2/s1 [11]));
 OR2_X1 \V2/A1/A2/A1/M4/_0_  (.A1(\V2/A1/A2/A1/M4/c1 ),
    .A2(\V2/A1/A2/A1/M4/c2 ),
    .ZN(\V2/A1/A2/c1 ));
 AND2_X1 \V2/A1/A2/A2/M1/M1/_0_  (.A1(\V2/v2 [12]),
    .A2(\V2/v3 [12]),
    .ZN(\V2/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M1/M1/_1_  (.A(\V2/v2 [12]),
    .B(\V2/v3 [12]),
    .Z(\V2/A1/A2/A2/M1/s1 ));
 AND2_X1 \V2/A1/A2/A2/M1/M2/_0_  (.A1(\V2/A1/A2/A2/M1/s1 ),
    .A2(\V2/A1/A2/c1 ),
    .ZN(\V2/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M1/M2/_1_  (.A(\V2/A1/A2/A2/M1/s1 ),
    .B(\V2/A1/A2/c1 ),
    .Z(\V2/s1 [12]));
 OR2_X1 \V2/A1/A2/A2/M1/_0_  (.A1(\V2/A1/A2/A2/M1/c1 ),
    .A2(\V2/A1/A2/A2/M1/c2 ),
    .ZN(\V2/A1/A2/A2/c1 ));
 AND2_X1 \V2/A1/A2/A2/M2/M1/_0_  (.A1(\V2/v2 [13]),
    .A2(\V2/v3 [13]),
    .ZN(\V2/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M2/M1/_1_  (.A(\V2/v2 [13]),
    .B(\V2/v3 [13]),
    .Z(\V2/A1/A2/A2/M2/s1 ));
 AND2_X1 \V2/A1/A2/A2/M2/M2/_0_  (.A1(\V2/A1/A2/A2/M2/s1 ),
    .A2(\V2/A1/A2/A2/c1 ),
    .ZN(\V2/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M2/M2/_1_  (.A(\V2/A1/A2/A2/M2/s1 ),
    .B(\V2/A1/A2/A2/c1 ),
    .Z(\V2/s1 [13]));
 OR2_X1 \V2/A1/A2/A2/M2/_0_  (.A1(\V2/A1/A2/A2/M2/c1 ),
    .A2(\V2/A1/A2/A2/M2/c2 ),
    .ZN(\V2/A1/A2/A2/c2 ));
 AND2_X1 \V2/A1/A2/A2/M3/M1/_0_  (.A1(\V2/v2 [14]),
    .A2(\V2/v3 [14]),
    .ZN(\V2/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M3/M1/_1_  (.A(\V2/v2 [14]),
    .B(\V2/v3 [14]),
    .Z(\V2/A1/A2/A2/M3/s1 ));
 AND2_X1 \V2/A1/A2/A2/M3/M2/_0_  (.A1(\V2/A1/A2/A2/M3/s1 ),
    .A2(\V2/A1/A2/A2/c2 ),
    .ZN(\V2/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M3/M2/_1_  (.A(\V2/A1/A2/A2/M3/s1 ),
    .B(\V2/A1/A2/A2/c2 ),
    .Z(\V2/s1 [14]));
 OR2_X1 \V2/A1/A2/A2/M3/_0_  (.A1(\V2/A1/A2/A2/M3/c1 ),
    .A2(\V2/A1/A2/A2/M3/c2 ),
    .ZN(\V2/A1/A2/A2/c3 ));
 AND2_X1 \V2/A1/A2/A2/M4/M1/_0_  (.A1(\V2/v2 [15]),
    .A2(\V2/v3 [15]),
    .ZN(\V2/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M4/M1/_1_  (.A(\V2/v2 [15]),
    .B(\V2/v3 [15]),
    .Z(\V2/A1/A2/A2/M4/s1 ));
 AND2_X1 \V2/A1/A2/A2/M4/M2/_0_  (.A1(\V2/A1/A2/A2/M4/s1 ),
    .A2(\V2/A1/A2/A2/c3 ),
    .ZN(\V2/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M4/M2/_1_  (.A(\V2/A1/A2/A2/M4/s1 ),
    .B(\V2/A1/A2/A2/c3 ),
    .Z(\V2/s1 [15]));
 OR2_X1 \V2/A1/A2/A2/M4/_0_  (.A1(\V2/A1/A2/A2/M4/c1 ),
    .A2(\V2/A1/A2/A2/M4/c2 ),
    .ZN(\V2/c1 ));
 AND2_X1 \V2/A2/A1/A1/M1/M1/_0_  (.A1(\V2/s1 [0]),
    .A2(\V2/v1 [8]),
    .ZN(\V2/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M1/M1/_1_  (.A(\V2/s1 [0]),
    .B(\V2/v1 [8]),
    .Z(\V2/A2/A1/A1/M1/s1 ));
 AND2_X1 \V2/A2/A1/A1/M1/M2/_0_  (.A1(\V2/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M1/M2/_1_  (.A(\V2/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v2[8]));
 OR2_X1 \V2/A2/A1/A1/M1/_0_  (.A1(\V2/A2/A1/A1/M1/c1 ),
    .A2(\V2/A2/A1/A1/M1/c2 ),
    .ZN(\V2/A2/A1/A1/c1 ));
 AND2_X1 \V2/A2/A1/A1/M2/M1/_0_  (.A1(\V2/s1 [1]),
    .A2(\V2/v1 [9]),
    .ZN(\V2/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M2/M1/_1_  (.A(\V2/s1 [1]),
    .B(\V2/v1 [9]),
    .Z(\V2/A2/A1/A1/M2/s1 ));
 AND2_X1 \V2/A2/A1/A1/M2/M2/_0_  (.A1(\V2/A2/A1/A1/M2/s1 ),
    .A2(\V2/A2/A1/A1/c1 ),
    .ZN(\V2/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M2/M2/_1_  (.A(\V2/A2/A1/A1/M2/s1 ),
    .B(\V2/A2/A1/A1/c1 ),
    .Z(v2[9]));
 OR2_X1 \V2/A2/A1/A1/M2/_0_  (.A1(\V2/A2/A1/A1/M2/c1 ),
    .A2(\V2/A2/A1/A1/M2/c2 ),
    .ZN(\V2/A2/A1/A1/c2 ));
 AND2_X1 \V2/A2/A1/A1/M3/M1/_0_  (.A1(\V2/s1 [2]),
    .A2(\V2/v1 [10]),
    .ZN(\V2/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M3/M1/_1_  (.A(\V2/s1 [2]),
    .B(\V2/v1 [10]),
    .Z(\V2/A2/A1/A1/M3/s1 ));
 AND2_X1 \V2/A2/A1/A1/M3/M2/_0_  (.A1(\V2/A2/A1/A1/M3/s1 ),
    .A2(\V2/A2/A1/A1/c2 ),
    .ZN(\V2/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M3/M2/_1_  (.A(\V2/A2/A1/A1/M3/s1 ),
    .B(\V2/A2/A1/A1/c2 ),
    .Z(v2[10]));
 OR2_X1 \V2/A2/A1/A1/M3/_0_  (.A1(\V2/A2/A1/A1/M3/c1 ),
    .A2(\V2/A2/A1/A1/M3/c2 ),
    .ZN(\V2/A2/A1/A1/c3 ));
 AND2_X1 \V2/A2/A1/A1/M4/M1/_0_  (.A1(\V2/s1 [3]),
    .A2(\V2/v1 [11]),
    .ZN(\V2/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M4/M1/_1_  (.A(\V2/s1 [3]),
    .B(\V2/v1 [11]),
    .Z(\V2/A2/A1/A1/M4/s1 ));
 AND2_X1 \V2/A2/A1/A1/M4/M2/_0_  (.A1(\V2/A2/A1/A1/M4/s1 ),
    .A2(\V2/A2/A1/A1/c3 ),
    .ZN(\V2/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M4/M2/_1_  (.A(\V2/A2/A1/A1/M4/s1 ),
    .B(\V2/A2/A1/A1/c3 ),
    .Z(v2[11]));
 OR2_X1 \V2/A2/A1/A1/M4/_0_  (.A1(\V2/A2/A1/A1/M4/c1 ),
    .A2(\V2/A2/A1/A1/M4/c2 ),
    .ZN(\V2/A2/A1/c1 ));
 AND2_X1 \V2/A2/A1/A2/M1/M1/_0_  (.A1(\V2/s1 [4]),
    .A2(\V2/v1 [12]),
    .ZN(\V2/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M1/M1/_1_  (.A(\V2/s1 [4]),
    .B(\V2/v1 [12]),
    .Z(\V2/A2/A1/A2/M1/s1 ));
 AND2_X1 \V2/A2/A1/A2/M1/M2/_0_  (.A1(\V2/A2/A1/A2/M1/s1 ),
    .A2(\V2/A2/A1/c1 ),
    .ZN(\V2/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M1/M2/_1_  (.A(\V2/A2/A1/A2/M1/s1 ),
    .B(\V2/A2/A1/c1 ),
    .Z(v2[12]));
 OR2_X1 \V2/A2/A1/A2/M1/_0_  (.A1(\V2/A2/A1/A2/M1/c1 ),
    .A2(\V2/A2/A1/A2/M1/c2 ),
    .ZN(\V2/A2/A1/A2/c1 ));
 AND2_X1 \V2/A2/A1/A2/M2/M1/_0_  (.A1(\V2/s1 [5]),
    .A2(\V2/v1 [13]),
    .ZN(\V2/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M2/M1/_1_  (.A(\V2/s1 [5]),
    .B(\V2/v1 [13]),
    .Z(\V2/A2/A1/A2/M2/s1 ));
 AND2_X1 \V2/A2/A1/A2/M2/M2/_0_  (.A1(\V2/A2/A1/A2/M2/s1 ),
    .A2(\V2/A2/A1/A2/c1 ),
    .ZN(\V2/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M2/M2/_1_  (.A(\V2/A2/A1/A2/M2/s1 ),
    .B(\V2/A2/A1/A2/c1 ),
    .Z(v2[13]));
 OR2_X1 \V2/A2/A1/A2/M2/_0_  (.A1(\V2/A2/A1/A2/M2/c1 ),
    .A2(\V2/A2/A1/A2/M2/c2 ),
    .ZN(\V2/A2/A1/A2/c2 ));
 AND2_X1 \V2/A2/A1/A2/M3/M1/_0_  (.A1(\V2/s1 [6]),
    .A2(\V2/v1 [14]),
    .ZN(\V2/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M3/M1/_1_  (.A(\V2/s1 [6]),
    .B(\V2/v1 [14]),
    .Z(\V2/A2/A1/A2/M3/s1 ));
 AND2_X1 \V2/A2/A1/A2/M3/M2/_0_  (.A1(\V2/A2/A1/A2/M3/s1 ),
    .A2(\V2/A2/A1/A2/c2 ),
    .ZN(\V2/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M3/M2/_1_  (.A(\V2/A2/A1/A2/M3/s1 ),
    .B(\V2/A2/A1/A2/c2 ),
    .Z(v2[14]));
 OR2_X1 \V2/A2/A1/A2/M3/_0_  (.A1(\V2/A2/A1/A2/M3/c1 ),
    .A2(\V2/A2/A1/A2/M3/c2 ),
    .ZN(\V2/A2/A1/A2/c3 ));
 AND2_X1 \V2/A2/A1/A2/M4/M1/_0_  (.A1(\V2/s1 [7]),
    .A2(\V2/v1 [15]),
    .ZN(\V2/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M4/M1/_1_  (.A(\V2/s1 [7]),
    .B(\V2/v1 [15]),
    .Z(\V2/A2/A1/A2/M4/s1 ));
 AND2_X1 \V2/A2/A1/A2/M4/M2/_0_  (.A1(\V2/A2/A1/A2/M4/s1 ),
    .A2(\V2/A2/A1/A2/c3 ),
    .ZN(\V2/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M4/M2/_1_  (.A(\V2/A2/A1/A2/M4/s1 ),
    .B(\V2/A2/A1/A2/c3 ),
    .Z(v2[15]));
 OR2_X1 \V2/A2/A1/A2/M4/_0_  (.A1(\V2/A2/A1/A2/M4/c1 ),
    .A2(\V2/A2/A1/A2/M4/c2 ),
    .ZN(\V2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A1/M1/M1/_0_  (.A1(\V2/s1 [8]),
    .A2(ground),
    .ZN(\V2/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M1/M1/_1_  (.A(\V2/s1 [8]),
    .B(ground),
    .Z(\V2/A2/A2/A1/M1/s1 ));
 AND2_X1 \V2/A2/A2/A1/M1/M2/_0_  (.A1(\V2/A2/A2/A1/M1/s1 ),
    .A2(\V2/A2/c1 ),
    .ZN(\V2/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M1/M2/_1_  (.A(\V2/A2/A2/A1/M1/s1 ),
    .B(\V2/A2/c1 ),
    .Z(\V2/s2 [8]));
 OR2_X1 \V2/A2/A2/A1/M1/_0_  (.A1(\V2/A2/A2/A1/M1/c1 ),
    .A2(\V2/A2/A2/A1/M1/c2 ),
    .ZN(\V2/A2/A2/A1/c1 ));
 AND2_X1 \V2/A2/A2/A1/M2/M1/_0_  (.A1(\V2/s1 [9]),
    .A2(ground),
    .ZN(\V2/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M2/M1/_1_  (.A(\V2/s1 [9]),
    .B(ground),
    .Z(\V2/A2/A2/A1/M2/s1 ));
 AND2_X1 \V2/A2/A2/A1/M2/M2/_0_  (.A1(\V2/A2/A2/A1/M2/s1 ),
    .A2(\V2/A2/A2/A1/c1 ),
    .ZN(\V2/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M2/M2/_1_  (.A(\V2/A2/A2/A1/M2/s1 ),
    .B(\V2/A2/A2/A1/c1 ),
    .Z(\V2/s2 [9]));
 OR2_X1 \V2/A2/A2/A1/M2/_0_  (.A1(\V2/A2/A2/A1/M2/c1 ),
    .A2(\V2/A2/A2/A1/M2/c2 ),
    .ZN(\V2/A2/A2/A1/c2 ));
 AND2_X1 \V2/A2/A2/A1/M3/M1/_0_  (.A1(\V2/s1 [10]),
    .A2(ground),
    .ZN(\V2/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M3/M1/_1_  (.A(\V2/s1 [10]),
    .B(ground),
    .Z(\V2/A2/A2/A1/M3/s1 ));
 AND2_X1 \V2/A2/A2/A1/M3/M2/_0_  (.A1(\V2/A2/A2/A1/M3/s1 ),
    .A2(\V2/A2/A2/A1/c2 ),
    .ZN(\V2/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M3/M2/_1_  (.A(\V2/A2/A2/A1/M3/s1 ),
    .B(\V2/A2/A2/A1/c2 ),
    .Z(\V2/s2 [10]));
 OR2_X1 \V2/A2/A2/A1/M3/_0_  (.A1(\V2/A2/A2/A1/M3/c1 ),
    .A2(\V2/A2/A2/A1/M3/c2 ),
    .ZN(\V2/A2/A2/A1/c3 ));
 AND2_X1 \V2/A2/A2/A1/M4/M1/_0_  (.A1(\V2/s1 [11]),
    .A2(ground),
    .ZN(\V2/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M4/M1/_1_  (.A(\V2/s1 [11]),
    .B(ground),
    .Z(\V2/A2/A2/A1/M4/s1 ));
 AND2_X1 \V2/A2/A2/A1/M4/M2/_0_  (.A1(\V2/A2/A2/A1/M4/s1 ),
    .A2(\V2/A2/A2/A1/c3 ),
    .ZN(\V2/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M4/M2/_1_  (.A(\V2/A2/A2/A1/M4/s1 ),
    .B(\V2/A2/A2/A1/c3 ),
    .Z(\V2/s2 [11]));
 OR2_X1 \V2/A2/A2/A1/M4/_0_  (.A1(\V2/A2/A2/A1/M4/c1 ),
    .A2(\V2/A2/A2/A1/M4/c2 ),
    .ZN(\V2/A2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A2/M1/M1/_0_  (.A1(\V2/s1 [12]),
    .A2(ground),
    .ZN(\V2/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M1/M1/_1_  (.A(\V2/s1 [12]),
    .B(ground),
    .Z(\V2/A2/A2/A2/M1/s1 ));
 AND2_X1 \V2/A2/A2/A2/M1/M2/_0_  (.A1(\V2/A2/A2/A2/M1/s1 ),
    .A2(\V2/A2/A2/c1 ),
    .ZN(\V2/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M1/M2/_1_  (.A(\V2/A2/A2/A2/M1/s1 ),
    .B(\V2/A2/A2/c1 ),
    .Z(\V2/s2 [12]));
 OR2_X1 \V2/A2/A2/A2/M1/_0_  (.A1(\V2/A2/A2/A2/M1/c1 ),
    .A2(\V2/A2/A2/A2/M1/c2 ),
    .ZN(\V2/A2/A2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A2/M2/M1/_0_  (.A1(\V2/s1 [13]),
    .A2(ground),
    .ZN(\V2/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M2/M1/_1_  (.A(\V2/s1 [13]),
    .B(ground),
    .Z(\V2/A2/A2/A2/M2/s1 ));
 AND2_X1 \V2/A2/A2/A2/M2/M2/_0_  (.A1(\V2/A2/A2/A2/M2/s1 ),
    .A2(\V2/A2/A2/A2/c1 ),
    .ZN(\V2/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M2/M2/_1_  (.A(\V2/A2/A2/A2/M2/s1 ),
    .B(\V2/A2/A2/A2/c1 ),
    .Z(\V2/s2 [13]));
 OR2_X1 \V2/A2/A2/A2/M2/_0_  (.A1(\V2/A2/A2/A2/M2/c1 ),
    .A2(\V2/A2/A2/A2/M2/c2 ),
    .ZN(\V2/A2/A2/A2/c2 ));
 AND2_X1 \V2/A2/A2/A2/M3/M1/_0_  (.A1(\V2/s1 [14]),
    .A2(ground),
    .ZN(\V2/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M3/M1/_1_  (.A(\V2/s1 [14]),
    .B(ground),
    .Z(\V2/A2/A2/A2/M3/s1 ));
 AND2_X1 \V2/A2/A2/A2/M3/M2/_0_  (.A1(\V2/A2/A2/A2/M3/s1 ),
    .A2(\V2/A2/A2/A2/c2 ),
    .ZN(\V2/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M3/M2/_1_  (.A(\V2/A2/A2/A2/M3/s1 ),
    .B(\V2/A2/A2/A2/c2 ),
    .Z(\V2/s2 [14]));
 OR2_X1 \V2/A2/A2/A2/M3/_0_  (.A1(\V2/A2/A2/A2/M3/c1 ),
    .A2(\V2/A2/A2/A2/M3/c2 ),
    .ZN(\V2/A2/A2/A2/c3 ));
 AND2_X1 \V2/A2/A2/A2/M4/M1/_0_  (.A1(\V2/s1 [15]),
    .A2(ground),
    .ZN(\V2/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M4/M1/_1_  (.A(\V2/s1 [15]),
    .B(ground),
    .Z(\V2/A2/A2/A2/M4/s1 ));
 AND2_X1 \V2/A2/A2/A2/M4/M2/_0_  (.A1(\V2/A2/A2/A2/M4/s1 ),
    .A2(\V2/A2/A2/A2/c3 ),
    .ZN(\V2/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M4/M2/_1_  (.A(\V2/A2/A2/A2/M4/s1 ),
    .B(\V2/A2/A2/A2/c3 ),
    .Z(\V2/s2 [15]));
 OR2_X1 \V2/A2/A2/A2/M4/_0_  (.A1(\V2/A2/A2/A2/M4/c1 ),
    .A2(\V2/A2/A2/A2/M4/c2 ),
    .ZN(\V2/c2 ));
 AND2_X1 \V2/A3/A1/A1/M1/M1/_0_  (.A1(\V2/v4 [0]),
    .A2(\V2/s2 [8]),
    .ZN(\V2/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M1/M1/_1_  (.A(\V2/v4 [0]),
    .B(\V2/s2 [8]),
    .Z(\V2/A3/A1/A1/M1/s1 ));
 AND2_X1 \V2/A3/A1/A1/M1/M2/_0_  (.A1(\V2/A3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M1/M2/_1_  (.A(\V2/A3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v2[16]));
 OR2_X1 \V2/A3/A1/A1/M1/_0_  (.A1(\V2/A3/A1/A1/M1/c1 ),
    .A2(\V2/A3/A1/A1/M1/c2 ),
    .ZN(\V2/A3/A1/A1/c1 ));
 AND2_X1 \V2/A3/A1/A1/M2/M1/_0_  (.A1(\V2/v4 [1]),
    .A2(\V2/s2 [9]),
    .ZN(\V2/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M2/M1/_1_  (.A(\V2/v4 [1]),
    .B(\V2/s2 [9]),
    .Z(\V2/A3/A1/A1/M2/s1 ));
 AND2_X1 \V2/A3/A1/A1/M2/M2/_0_  (.A1(\V2/A3/A1/A1/M2/s1 ),
    .A2(\V2/A3/A1/A1/c1 ),
    .ZN(\V2/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M2/M2/_1_  (.A(\V2/A3/A1/A1/M2/s1 ),
    .B(\V2/A3/A1/A1/c1 ),
    .Z(v2[17]));
 OR2_X1 \V2/A3/A1/A1/M2/_0_  (.A1(\V2/A3/A1/A1/M2/c1 ),
    .A2(\V2/A3/A1/A1/M2/c2 ),
    .ZN(\V2/A3/A1/A1/c2 ));
 AND2_X1 \V2/A3/A1/A1/M3/M1/_0_  (.A1(\V2/v4 [2]),
    .A2(\V2/s2 [10]),
    .ZN(\V2/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M3/M1/_1_  (.A(\V2/v4 [2]),
    .B(\V2/s2 [10]),
    .Z(\V2/A3/A1/A1/M3/s1 ));
 AND2_X1 \V2/A3/A1/A1/M3/M2/_0_  (.A1(\V2/A3/A1/A1/M3/s1 ),
    .A2(\V2/A3/A1/A1/c2 ),
    .ZN(\V2/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M3/M2/_1_  (.A(\V2/A3/A1/A1/M3/s1 ),
    .B(\V2/A3/A1/A1/c2 ),
    .Z(v2[18]));
 OR2_X1 \V2/A3/A1/A1/M3/_0_  (.A1(\V2/A3/A1/A1/M3/c1 ),
    .A2(\V2/A3/A1/A1/M3/c2 ),
    .ZN(\V2/A3/A1/A1/c3 ));
 AND2_X1 \V2/A3/A1/A1/M4/M1/_0_  (.A1(\V2/v4 [3]),
    .A2(\V2/s2 [11]),
    .ZN(\V2/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M4/M1/_1_  (.A(\V2/v4 [3]),
    .B(\V2/s2 [11]),
    .Z(\V2/A3/A1/A1/M4/s1 ));
 AND2_X1 \V2/A3/A1/A1/M4/M2/_0_  (.A1(\V2/A3/A1/A1/M4/s1 ),
    .A2(\V2/A3/A1/A1/c3 ),
    .ZN(\V2/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M4/M2/_1_  (.A(\V2/A3/A1/A1/M4/s1 ),
    .B(\V2/A3/A1/A1/c3 ),
    .Z(v2[19]));
 OR2_X1 \V2/A3/A1/A1/M4/_0_  (.A1(\V2/A3/A1/A1/M4/c1 ),
    .A2(\V2/A3/A1/A1/M4/c2 ),
    .ZN(\V2/A3/A1/c1 ));
 AND2_X1 \V2/A3/A1/A2/M1/M1/_0_  (.A1(\V2/v4 [4]),
    .A2(\V2/s2 [12]),
    .ZN(\V2/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M1/M1/_1_  (.A(\V2/v4 [4]),
    .B(\V2/s2 [12]),
    .Z(\V2/A3/A1/A2/M1/s1 ));
 AND2_X1 \V2/A3/A1/A2/M1/M2/_0_  (.A1(\V2/A3/A1/A2/M1/s1 ),
    .A2(\V2/A3/A1/c1 ),
    .ZN(\V2/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M1/M2/_1_  (.A(\V2/A3/A1/A2/M1/s1 ),
    .B(\V2/A3/A1/c1 ),
    .Z(v2[20]));
 OR2_X1 \V2/A3/A1/A2/M1/_0_  (.A1(\V2/A3/A1/A2/M1/c1 ),
    .A2(\V2/A3/A1/A2/M1/c2 ),
    .ZN(\V2/A3/A1/A2/c1 ));
 AND2_X1 \V2/A3/A1/A2/M2/M1/_0_  (.A1(\V2/v4 [5]),
    .A2(\V2/s2 [13]),
    .ZN(\V2/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M2/M1/_1_  (.A(\V2/v4 [5]),
    .B(\V2/s2 [13]),
    .Z(\V2/A3/A1/A2/M2/s1 ));
 AND2_X1 \V2/A3/A1/A2/M2/M2/_0_  (.A1(\V2/A3/A1/A2/M2/s1 ),
    .A2(\V2/A3/A1/A2/c1 ),
    .ZN(\V2/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M2/M2/_1_  (.A(\V2/A3/A1/A2/M2/s1 ),
    .B(\V2/A3/A1/A2/c1 ),
    .Z(v2[21]));
 OR2_X1 \V2/A3/A1/A2/M2/_0_  (.A1(\V2/A3/A1/A2/M2/c1 ),
    .A2(\V2/A3/A1/A2/M2/c2 ),
    .ZN(\V2/A3/A1/A2/c2 ));
 AND2_X1 \V2/A3/A1/A2/M3/M1/_0_  (.A1(\V2/v4 [6]),
    .A2(\V2/s2 [14]),
    .ZN(\V2/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M3/M1/_1_  (.A(\V2/v4 [6]),
    .B(\V2/s2 [14]),
    .Z(\V2/A3/A1/A2/M3/s1 ));
 AND2_X1 \V2/A3/A1/A2/M3/M2/_0_  (.A1(\V2/A3/A1/A2/M3/s1 ),
    .A2(\V2/A3/A1/A2/c2 ),
    .ZN(\V2/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M3/M2/_1_  (.A(\V2/A3/A1/A2/M3/s1 ),
    .B(\V2/A3/A1/A2/c2 ),
    .Z(v2[22]));
 OR2_X1 \V2/A3/A1/A2/M3/_0_  (.A1(\V2/A3/A1/A2/M3/c1 ),
    .A2(\V2/A3/A1/A2/M3/c2 ),
    .ZN(\V2/A3/A1/A2/c3 ));
 AND2_X1 \V2/A3/A1/A2/M4/M1/_0_  (.A1(\V2/v4 [7]),
    .A2(\V2/s2 [15]),
    .ZN(\V2/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M4/M1/_1_  (.A(\V2/v4 [7]),
    .B(\V2/s2 [15]),
    .Z(\V2/A3/A1/A2/M4/s1 ));
 AND2_X1 \V2/A3/A1/A2/M4/M2/_0_  (.A1(\V2/A3/A1/A2/M4/s1 ),
    .A2(\V2/A3/A1/A2/c3 ),
    .ZN(\V2/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M4/M2/_1_  (.A(\V2/A3/A1/A2/M4/s1 ),
    .B(\V2/A3/A1/A2/c3 ),
    .Z(v2[23]));
 OR2_X1 \V2/A3/A1/A2/M4/_0_  (.A1(\V2/A3/A1/A2/M4/c1 ),
    .A2(\V2/A3/A1/A2/M4/c2 ),
    .ZN(\V2/A3/c1 ));
 AND2_X1 \V2/A3/A2/A1/M1/M1/_0_  (.A1(\V2/v4 [8]),
    .A2(\V2/c3 ),
    .ZN(\V2/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M1/M1/_1_  (.A(\V2/v4 [8]),
    .B(\V2/c3 ),
    .Z(\V2/A3/A2/A1/M1/s1 ));
 AND2_X1 \V2/A3/A2/A1/M1/M2/_0_  (.A1(\V2/A3/A2/A1/M1/s1 ),
    .A2(\V2/A3/c1 ),
    .ZN(\V2/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M1/M2/_1_  (.A(\V2/A3/A2/A1/M1/s1 ),
    .B(\V2/A3/c1 ),
    .Z(v2[24]));
 OR2_X1 \V2/A3/A2/A1/M1/_0_  (.A1(\V2/A3/A2/A1/M1/c1 ),
    .A2(\V2/A3/A2/A1/M1/c2 ),
    .ZN(\V2/A3/A2/A1/c1 ));
 AND2_X1 \V2/A3/A2/A1/M2/M1/_0_  (.A1(\V2/v4 [9]),
    .A2(ground),
    .ZN(\V2/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M2/M1/_1_  (.A(\V2/v4 [9]),
    .B(ground),
    .Z(\V2/A3/A2/A1/M2/s1 ));
 AND2_X1 \V2/A3/A2/A1/M2/M2/_0_  (.A1(\V2/A3/A2/A1/M2/s1 ),
    .A2(\V2/A3/A2/A1/c1 ),
    .ZN(\V2/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M2/M2/_1_  (.A(\V2/A3/A2/A1/M2/s1 ),
    .B(\V2/A3/A2/A1/c1 ),
    .Z(v2[25]));
 OR2_X1 \V2/A3/A2/A1/M2/_0_  (.A1(\V2/A3/A2/A1/M2/c1 ),
    .A2(\V2/A3/A2/A1/M2/c2 ),
    .ZN(\V2/A3/A2/A1/c2 ));
 AND2_X1 \V2/A3/A2/A1/M3/M1/_0_  (.A1(\V2/v4 [10]),
    .A2(ground),
    .ZN(\V2/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M3/M1/_1_  (.A(\V2/v4 [10]),
    .B(ground),
    .Z(\V2/A3/A2/A1/M3/s1 ));
 AND2_X1 \V2/A3/A2/A1/M3/M2/_0_  (.A1(\V2/A3/A2/A1/M3/s1 ),
    .A2(\V2/A3/A2/A1/c2 ),
    .ZN(\V2/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M3/M2/_1_  (.A(\V2/A3/A2/A1/M3/s1 ),
    .B(\V2/A3/A2/A1/c2 ),
    .Z(v2[26]));
 OR2_X1 \V2/A3/A2/A1/M3/_0_  (.A1(\V2/A3/A2/A1/M3/c1 ),
    .A2(\V2/A3/A2/A1/M3/c2 ),
    .ZN(\V2/A3/A2/A1/c3 ));
 AND2_X1 \V2/A3/A2/A1/M4/M1/_0_  (.A1(\V2/v4 [11]),
    .A2(ground),
    .ZN(\V2/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M4/M1/_1_  (.A(\V2/v4 [11]),
    .B(ground),
    .Z(\V2/A3/A2/A1/M4/s1 ));
 AND2_X1 \V2/A3/A2/A1/M4/M2/_0_  (.A1(\V2/A3/A2/A1/M4/s1 ),
    .A2(\V2/A3/A2/A1/c3 ),
    .ZN(\V2/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M4/M2/_1_  (.A(\V2/A3/A2/A1/M4/s1 ),
    .B(\V2/A3/A2/A1/c3 ),
    .Z(v2[27]));
 OR2_X1 \V2/A3/A2/A1/M4/_0_  (.A1(\V2/A3/A2/A1/M4/c1 ),
    .A2(\V2/A3/A2/A1/M4/c2 ),
    .ZN(\V2/A3/A2/c1 ));
 AND2_X1 \V2/A3/A2/A2/M1/M1/_0_  (.A1(\V2/v4 [12]),
    .A2(ground),
    .ZN(\V2/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M1/M1/_1_  (.A(\V2/v4 [12]),
    .B(ground),
    .Z(\V2/A3/A2/A2/M1/s1 ));
 AND2_X1 \V2/A3/A2/A2/M1/M2/_0_  (.A1(\V2/A3/A2/A2/M1/s1 ),
    .A2(\V2/A3/A2/c1 ),
    .ZN(\V2/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M1/M2/_1_  (.A(\V2/A3/A2/A2/M1/s1 ),
    .B(\V2/A3/A2/c1 ),
    .Z(v2[28]));
 OR2_X1 \V2/A3/A2/A2/M1/_0_  (.A1(\V2/A3/A2/A2/M1/c1 ),
    .A2(\V2/A3/A2/A2/M1/c2 ),
    .ZN(\V2/A3/A2/A2/c1 ));
 AND2_X1 \V2/A3/A2/A2/M2/M1/_0_  (.A1(\V2/v4 [13]),
    .A2(ground),
    .ZN(\V2/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M2/M1/_1_  (.A(\V2/v4 [13]),
    .B(ground),
    .Z(\V2/A3/A2/A2/M2/s1 ));
 AND2_X1 \V2/A3/A2/A2/M2/M2/_0_  (.A1(\V2/A3/A2/A2/M2/s1 ),
    .A2(\V2/A3/A2/A2/c1 ),
    .ZN(\V2/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M2/M2/_1_  (.A(\V2/A3/A2/A2/M2/s1 ),
    .B(\V2/A3/A2/A2/c1 ),
    .Z(v2[29]));
 OR2_X1 \V2/A3/A2/A2/M2/_0_  (.A1(\V2/A3/A2/A2/M2/c1 ),
    .A2(\V2/A3/A2/A2/M2/c2 ),
    .ZN(\V2/A3/A2/A2/c2 ));
 AND2_X1 \V2/A3/A2/A2/M3/M1/_0_  (.A1(\V2/v4 [14]),
    .A2(ground),
    .ZN(\V2/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M3/M1/_1_  (.A(\V2/v4 [14]),
    .B(ground),
    .Z(\V2/A3/A2/A2/M3/s1 ));
 AND2_X1 \V2/A3/A2/A2/M3/M2/_0_  (.A1(\V2/A3/A2/A2/M3/s1 ),
    .A2(\V2/A3/A2/A2/c2 ),
    .ZN(\V2/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M3/M2/_1_  (.A(\V2/A3/A2/A2/M3/s1 ),
    .B(\V2/A3/A2/A2/c2 ),
    .Z(v2[30]));
 OR2_X1 \V2/A3/A2/A2/M3/_0_  (.A1(\V2/A3/A2/A2/M3/c1 ),
    .A2(\V2/A3/A2/A2/M3/c2 ),
    .ZN(\V2/A3/A2/A2/c3 ));
 AND2_X1 \V2/A3/A2/A2/M4/M1/_0_  (.A1(\V2/v4 [15]),
    .A2(ground),
    .ZN(\V2/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M4/M1/_1_  (.A(\V2/v4 [15]),
    .B(ground),
    .Z(\V2/A3/A2/A2/M4/s1 ));
 AND2_X1 \V2/A3/A2/A2/M4/M2/_0_  (.A1(\V2/A3/A2/A2/M4/s1 ),
    .A2(\V2/A3/A2/A2/c3 ),
    .ZN(\V2/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M4/M2/_1_  (.A(\V2/A3/A2/A2/M4/s1 ),
    .B(\V2/A3/A2/A2/c3 ),
    .Z(v2[31]));
 OR2_X1 \V2/A3/A2/A2/M4/_0_  (.A1(\V2/A3/A2/A2/M4/c1 ),
    .A2(\V2/A3/A2/A2/M4/c2 ),
    .ZN(\V2/overflow ));
 AND2_X1 \V2/V1/A1/A1/M1/M1/_0_  (.A1(\V2/V1/v2 [0]),
    .A2(\V2/V1/v3 [0]),
    .ZN(\V2/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M1/M1/_1_  (.A(\V2/V1/v2 [0]),
    .B(\V2/V1/v3 [0]),
    .Z(\V2/V1/A1/A1/M1/s1 ));
 AND2_X1 \V2/V1/A1/A1/M1/M2/_0_  (.A1(\V2/V1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M1/M2/_1_  (.A(\V2/V1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/s1 [0]));
 OR2_X1 \V2/V1/A1/A1/M1/_0_  (.A1(\V2/V1/A1/A1/M1/c1 ),
    .A2(\V2/V1/A1/A1/M1/c2 ),
    .ZN(\V2/V1/A1/A1/c1 ));
 AND2_X1 \V2/V1/A1/A1/M2/M1/_0_  (.A1(\V2/V1/v2 [1]),
    .A2(\V2/V1/v3 [1]),
    .ZN(\V2/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M2/M1/_1_  (.A(\V2/V1/v2 [1]),
    .B(\V2/V1/v3 [1]),
    .Z(\V2/V1/A1/A1/M2/s1 ));
 AND2_X1 \V2/V1/A1/A1/M2/M2/_0_  (.A1(\V2/V1/A1/A1/M2/s1 ),
    .A2(\V2/V1/A1/A1/c1 ),
    .ZN(\V2/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M2/M2/_1_  (.A(\V2/V1/A1/A1/M2/s1 ),
    .B(\V2/V1/A1/A1/c1 ),
    .Z(\V2/V1/s1 [1]));
 OR2_X1 \V2/V1/A1/A1/M2/_0_  (.A1(\V2/V1/A1/A1/M2/c1 ),
    .A2(\V2/V1/A1/A1/M2/c2 ),
    .ZN(\V2/V1/A1/A1/c2 ));
 AND2_X1 \V2/V1/A1/A1/M3/M1/_0_  (.A1(\V2/V1/v2 [2]),
    .A2(\V2/V1/v3 [2]),
    .ZN(\V2/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M3/M1/_1_  (.A(\V2/V1/v2 [2]),
    .B(\V2/V1/v3 [2]),
    .Z(\V2/V1/A1/A1/M3/s1 ));
 AND2_X1 \V2/V1/A1/A1/M3/M2/_0_  (.A1(\V2/V1/A1/A1/M3/s1 ),
    .A2(\V2/V1/A1/A1/c2 ),
    .ZN(\V2/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M3/M2/_1_  (.A(\V2/V1/A1/A1/M3/s1 ),
    .B(\V2/V1/A1/A1/c2 ),
    .Z(\V2/V1/s1 [2]));
 OR2_X1 \V2/V1/A1/A1/M3/_0_  (.A1(\V2/V1/A1/A1/M3/c1 ),
    .A2(\V2/V1/A1/A1/M3/c2 ),
    .ZN(\V2/V1/A1/A1/c3 ));
 AND2_X1 \V2/V1/A1/A1/M4/M1/_0_  (.A1(\V2/V1/v2 [3]),
    .A2(\V2/V1/v3 [3]),
    .ZN(\V2/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M4/M1/_1_  (.A(\V2/V1/v2 [3]),
    .B(\V2/V1/v3 [3]),
    .Z(\V2/V1/A1/A1/M4/s1 ));
 AND2_X1 \V2/V1/A1/A1/M4/M2/_0_  (.A1(\V2/V1/A1/A1/M4/s1 ),
    .A2(\V2/V1/A1/A1/c3 ),
    .ZN(\V2/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M4/M2/_1_  (.A(\V2/V1/A1/A1/M4/s1 ),
    .B(\V2/V1/A1/A1/c3 ),
    .Z(\V2/V1/s1 [3]));
 OR2_X1 \V2/V1/A1/A1/M4/_0_  (.A1(\V2/V1/A1/A1/M4/c1 ),
    .A2(\V2/V1/A1/A1/M4/c2 ),
    .ZN(\V2/V1/A1/c1 ));
 AND2_X1 \V2/V1/A1/A2/M1/M1/_0_  (.A1(\V2/V1/v2 [4]),
    .A2(\V2/V1/v3 [4]),
    .ZN(\V2/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M1/M1/_1_  (.A(\V2/V1/v2 [4]),
    .B(\V2/V1/v3 [4]),
    .Z(\V2/V1/A1/A2/M1/s1 ));
 AND2_X1 \V2/V1/A1/A2/M1/M2/_0_  (.A1(\V2/V1/A1/A2/M1/s1 ),
    .A2(\V2/V1/A1/c1 ),
    .ZN(\V2/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M1/M2/_1_  (.A(\V2/V1/A1/A2/M1/s1 ),
    .B(\V2/V1/A1/c1 ),
    .Z(\V2/V1/s1 [4]));
 OR2_X1 \V2/V1/A1/A2/M1/_0_  (.A1(\V2/V1/A1/A2/M1/c1 ),
    .A2(\V2/V1/A1/A2/M1/c2 ),
    .ZN(\V2/V1/A1/A2/c1 ));
 AND2_X1 \V2/V1/A1/A2/M2/M1/_0_  (.A1(\V2/V1/v2 [5]),
    .A2(\V2/V1/v3 [5]),
    .ZN(\V2/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M2/M1/_1_  (.A(\V2/V1/v2 [5]),
    .B(\V2/V1/v3 [5]),
    .Z(\V2/V1/A1/A2/M2/s1 ));
 AND2_X1 \V2/V1/A1/A2/M2/M2/_0_  (.A1(\V2/V1/A1/A2/M2/s1 ),
    .A2(\V2/V1/A1/A2/c1 ),
    .ZN(\V2/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M2/M2/_1_  (.A(\V2/V1/A1/A2/M2/s1 ),
    .B(\V2/V1/A1/A2/c1 ),
    .Z(\V2/V1/s1 [5]));
 OR2_X1 \V2/V1/A1/A2/M2/_0_  (.A1(\V2/V1/A1/A2/M2/c1 ),
    .A2(\V2/V1/A1/A2/M2/c2 ),
    .ZN(\V2/V1/A1/A2/c2 ));
 AND2_X1 \V2/V1/A1/A2/M3/M1/_0_  (.A1(\V2/V1/v2 [6]),
    .A2(\V2/V1/v3 [6]),
    .ZN(\V2/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M3/M1/_1_  (.A(\V2/V1/v2 [6]),
    .B(\V2/V1/v3 [6]),
    .Z(\V2/V1/A1/A2/M3/s1 ));
 AND2_X1 \V2/V1/A1/A2/M3/M2/_0_  (.A1(\V2/V1/A1/A2/M3/s1 ),
    .A2(\V2/V1/A1/A2/c2 ),
    .ZN(\V2/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M3/M2/_1_  (.A(\V2/V1/A1/A2/M3/s1 ),
    .B(\V2/V1/A1/A2/c2 ),
    .Z(\V2/V1/s1 [6]));
 OR2_X1 \V2/V1/A1/A2/M3/_0_  (.A1(\V2/V1/A1/A2/M3/c1 ),
    .A2(\V2/V1/A1/A2/M3/c2 ),
    .ZN(\V2/V1/A1/A2/c3 ));
 AND2_X1 \V2/V1/A1/A2/M4/M1/_0_  (.A1(\V2/V1/v2 [7]),
    .A2(\V2/V1/v3 [7]),
    .ZN(\V2/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M4/M1/_1_  (.A(\V2/V1/v2 [7]),
    .B(\V2/V1/v3 [7]),
    .Z(\V2/V1/A1/A2/M4/s1 ));
 AND2_X1 \V2/V1/A1/A2/M4/M2/_0_  (.A1(\V2/V1/A1/A2/M4/s1 ),
    .A2(\V2/V1/A1/A2/c3 ),
    .ZN(\V2/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M4/M2/_1_  (.A(\V2/V1/A1/A2/M4/s1 ),
    .B(\V2/V1/A1/A2/c3 ),
    .Z(\V2/V1/s1 [7]));
 OR2_X1 \V2/V1/A1/A2/M4/_0_  (.A1(\V2/V1/A1/A2/M4/c1 ),
    .A2(\V2/V1/A1/A2/M4/c2 ),
    .ZN(\V2/V1/c1 ));
 AND2_X1 \V2/V1/A2/A1/M1/M1/_0_  (.A1(\V2/V1/s1 [0]),
    .A2(\V2/V1/v1 [4]),
    .ZN(\V2/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M1/M1/_1_  (.A(\V2/V1/s1 [0]),
    .B(\V2/V1/v1 [4]),
    .Z(\V2/V1/A2/A1/M1/s1 ));
 AND2_X1 \V2/V1/A2/A1/M1/M2/_0_  (.A1(\V2/V1/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M1/M2/_1_  (.A(\V2/V1/A2/A1/M1/s1 ),
    .B(ground),
    .Z(v2[4]));
 OR2_X1 \V2/V1/A2/A1/M1/_0_  (.A1(\V2/V1/A2/A1/M1/c1 ),
    .A2(\V2/V1/A2/A1/M1/c2 ),
    .ZN(\V2/V1/A2/A1/c1 ));
 AND2_X1 \V2/V1/A2/A1/M2/M1/_0_  (.A1(\V2/V1/s1 [1]),
    .A2(\V2/V1/v1 [5]),
    .ZN(\V2/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M2/M1/_1_  (.A(\V2/V1/s1 [1]),
    .B(\V2/V1/v1 [5]),
    .Z(\V2/V1/A2/A1/M2/s1 ));
 AND2_X1 \V2/V1/A2/A1/M2/M2/_0_  (.A1(\V2/V1/A2/A1/M2/s1 ),
    .A2(\V2/V1/A2/A1/c1 ),
    .ZN(\V2/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M2/M2/_1_  (.A(\V2/V1/A2/A1/M2/s1 ),
    .B(\V2/V1/A2/A1/c1 ),
    .Z(v2[5]));
 OR2_X1 \V2/V1/A2/A1/M2/_0_  (.A1(\V2/V1/A2/A1/M2/c1 ),
    .A2(\V2/V1/A2/A1/M2/c2 ),
    .ZN(\V2/V1/A2/A1/c2 ));
 AND2_X1 \V2/V1/A2/A1/M3/M1/_0_  (.A1(\V2/V1/s1 [2]),
    .A2(\V2/V1/v1 [6]),
    .ZN(\V2/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M3/M1/_1_  (.A(\V2/V1/s1 [2]),
    .B(\V2/V1/v1 [6]),
    .Z(\V2/V1/A2/A1/M3/s1 ));
 AND2_X1 \V2/V1/A2/A1/M3/M2/_0_  (.A1(\V2/V1/A2/A1/M3/s1 ),
    .A2(\V2/V1/A2/A1/c2 ),
    .ZN(\V2/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M3/M2/_1_  (.A(\V2/V1/A2/A1/M3/s1 ),
    .B(\V2/V1/A2/A1/c2 ),
    .Z(v2[6]));
 OR2_X1 \V2/V1/A2/A1/M3/_0_  (.A1(\V2/V1/A2/A1/M3/c1 ),
    .A2(\V2/V1/A2/A1/M3/c2 ),
    .ZN(\V2/V1/A2/A1/c3 ));
 AND2_X1 \V2/V1/A2/A1/M4/M1/_0_  (.A1(\V2/V1/s1 [3]),
    .A2(\V2/V1/v1 [7]),
    .ZN(\V2/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M4/M1/_1_  (.A(\V2/V1/s1 [3]),
    .B(\V2/V1/v1 [7]),
    .Z(\V2/V1/A2/A1/M4/s1 ));
 AND2_X1 \V2/V1/A2/A1/M4/M2/_0_  (.A1(\V2/V1/A2/A1/M4/s1 ),
    .A2(\V2/V1/A2/A1/c3 ),
    .ZN(\V2/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M4/M2/_1_  (.A(\V2/V1/A2/A1/M4/s1 ),
    .B(\V2/V1/A2/A1/c3 ),
    .Z(v2[7]));
 OR2_X1 \V2/V1/A2/A1/M4/_0_  (.A1(\V2/V1/A2/A1/M4/c1 ),
    .A2(\V2/V1/A2/A1/M4/c2 ),
    .ZN(\V2/V1/A2/c1 ));
 AND2_X1 \V2/V1/A2/A2/M1/M1/_0_  (.A1(\V2/V1/s1 [4]),
    .A2(ground),
    .ZN(\V2/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M1/M1/_1_  (.A(\V2/V1/s1 [4]),
    .B(ground),
    .Z(\V2/V1/A2/A2/M1/s1 ));
 AND2_X1 \V2/V1/A2/A2/M1/M2/_0_  (.A1(\V2/V1/A2/A2/M1/s1 ),
    .A2(\V2/V1/A2/c1 ),
    .ZN(\V2/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M1/M2/_1_  (.A(\V2/V1/A2/A2/M1/s1 ),
    .B(\V2/V1/A2/c1 ),
    .Z(\V2/V1/s2 [4]));
 OR2_X1 \V2/V1/A2/A2/M1/_0_  (.A1(\V2/V1/A2/A2/M1/c1 ),
    .A2(\V2/V1/A2/A2/M1/c2 ),
    .ZN(\V2/V1/A2/A2/c1 ));
 AND2_X1 \V2/V1/A2/A2/M2/M1/_0_  (.A1(\V2/V1/s1 [5]),
    .A2(ground),
    .ZN(\V2/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M2/M1/_1_  (.A(\V2/V1/s1 [5]),
    .B(ground),
    .Z(\V2/V1/A2/A2/M2/s1 ));
 AND2_X1 \V2/V1/A2/A2/M2/M2/_0_  (.A1(\V2/V1/A2/A2/M2/s1 ),
    .A2(\V2/V1/A2/A2/c1 ),
    .ZN(\V2/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M2/M2/_1_  (.A(\V2/V1/A2/A2/M2/s1 ),
    .B(\V2/V1/A2/A2/c1 ),
    .Z(\V2/V1/s2 [5]));
 OR2_X1 \V2/V1/A2/A2/M2/_0_  (.A1(\V2/V1/A2/A2/M2/c1 ),
    .A2(\V2/V1/A2/A2/M2/c2 ),
    .ZN(\V2/V1/A2/A2/c2 ));
 AND2_X1 \V2/V1/A2/A2/M3/M1/_0_  (.A1(\V2/V1/s1 [6]),
    .A2(ground),
    .ZN(\V2/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M3/M1/_1_  (.A(\V2/V1/s1 [6]),
    .B(ground),
    .Z(\V2/V1/A2/A2/M3/s1 ));
 AND2_X1 \V2/V1/A2/A2/M3/M2/_0_  (.A1(\V2/V1/A2/A2/M3/s1 ),
    .A2(\V2/V1/A2/A2/c2 ),
    .ZN(\V2/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M3/M2/_1_  (.A(\V2/V1/A2/A2/M3/s1 ),
    .B(\V2/V1/A2/A2/c2 ),
    .Z(\V2/V1/s2 [6]));
 OR2_X1 \V2/V1/A2/A2/M3/_0_  (.A1(\V2/V1/A2/A2/M3/c1 ),
    .A2(\V2/V1/A2/A2/M3/c2 ),
    .ZN(\V2/V1/A2/A2/c3 ));
 AND2_X1 \V2/V1/A2/A2/M4/M1/_0_  (.A1(\V2/V1/s1 [7]),
    .A2(ground),
    .ZN(\V2/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M4/M1/_1_  (.A(\V2/V1/s1 [7]),
    .B(ground),
    .Z(\V2/V1/A2/A2/M4/s1 ));
 AND2_X1 \V2/V1/A2/A2/M4/M2/_0_  (.A1(\V2/V1/A2/A2/M4/s1 ),
    .A2(\V2/V1/A2/A2/c3 ),
    .ZN(\V2/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M4/M2/_1_  (.A(\V2/V1/A2/A2/M4/s1 ),
    .B(\V2/V1/A2/A2/c3 ),
    .Z(\V2/V1/s2 [7]));
 OR2_X1 \V2/V1/A2/A2/M4/_0_  (.A1(\V2/V1/A2/A2/M4/c1 ),
    .A2(\V2/V1/A2/A2/M4/c2 ),
    .ZN(\V2/V1/c2 ));
 AND2_X1 \V2/V1/A3/A1/M1/M1/_0_  (.A1(\V2/V1/v4 [0]),
    .A2(\V2/V1/s2 [4]),
    .ZN(\V2/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M1/M1/_1_  (.A(\V2/V1/v4 [0]),
    .B(\V2/V1/s2 [4]),
    .Z(\V2/V1/A3/A1/M1/s1 ));
 AND2_X1 \V2/V1/A3/A1/M1/M2/_0_  (.A1(\V2/V1/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M1/M2/_1_  (.A(\V2/V1/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v1 [8]));
 OR2_X1 \V2/V1/A3/A1/M1/_0_  (.A1(\V2/V1/A3/A1/M1/c1 ),
    .A2(\V2/V1/A3/A1/M1/c2 ),
    .ZN(\V2/V1/A3/A1/c1 ));
 AND2_X1 \V2/V1/A3/A1/M2/M1/_0_  (.A1(\V2/V1/v4 [1]),
    .A2(\V2/V1/s2 [5]),
    .ZN(\V2/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M2/M1/_1_  (.A(\V2/V1/v4 [1]),
    .B(\V2/V1/s2 [5]),
    .Z(\V2/V1/A3/A1/M2/s1 ));
 AND2_X1 \V2/V1/A3/A1/M2/M2/_0_  (.A1(\V2/V1/A3/A1/M2/s1 ),
    .A2(\V2/V1/A3/A1/c1 ),
    .ZN(\V2/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M2/M2/_1_  (.A(\V2/V1/A3/A1/M2/s1 ),
    .B(\V2/V1/A3/A1/c1 ),
    .Z(\V2/v1 [9]));
 OR2_X1 \V2/V1/A3/A1/M2/_0_  (.A1(\V2/V1/A3/A1/M2/c1 ),
    .A2(\V2/V1/A3/A1/M2/c2 ),
    .ZN(\V2/V1/A3/A1/c2 ));
 AND2_X1 \V2/V1/A3/A1/M3/M1/_0_  (.A1(\V2/V1/v4 [2]),
    .A2(\V2/V1/s2 [6]),
    .ZN(\V2/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M3/M1/_1_  (.A(\V2/V1/v4 [2]),
    .B(\V2/V1/s2 [6]),
    .Z(\V2/V1/A3/A1/M3/s1 ));
 AND2_X1 \V2/V1/A3/A1/M3/M2/_0_  (.A1(\V2/V1/A3/A1/M3/s1 ),
    .A2(\V2/V1/A3/A1/c2 ),
    .ZN(\V2/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M3/M2/_1_  (.A(\V2/V1/A3/A1/M3/s1 ),
    .B(\V2/V1/A3/A1/c2 ),
    .Z(\V2/v1 [10]));
 OR2_X1 \V2/V1/A3/A1/M3/_0_  (.A1(\V2/V1/A3/A1/M3/c1 ),
    .A2(\V2/V1/A3/A1/M3/c2 ),
    .ZN(\V2/V1/A3/A1/c3 ));
 AND2_X1 \V2/V1/A3/A1/M4/M1/_0_  (.A1(\V2/V1/v4 [3]),
    .A2(\V2/V1/s2 [7]),
    .ZN(\V2/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M4/M1/_1_  (.A(\V2/V1/v4 [3]),
    .B(\V2/V1/s2 [7]),
    .Z(\V2/V1/A3/A1/M4/s1 ));
 AND2_X1 \V2/V1/A3/A1/M4/M2/_0_  (.A1(\V2/V1/A3/A1/M4/s1 ),
    .A2(\V2/V1/A3/A1/c3 ),
    .ZN(\V2/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M4/M2/_1_  (.A(\V2/V1/A3/A1/M4/s1 ),
    .B(\V2/V1/A3/A1/c3 ),
    .Z(\V2/v1 [11]));
 OR2_X1 \V2/V1/A3/A1/M4/_0_  (.A1(\V2/V1/A3/A1/M4/c1 ),
    .A2(\V2/V1/A3/A1/M4/c2 ),
    .ZN(\V2/V1/A3/c1 ));
 AND2_X1 \V2/V1/A3/A2/M1/M1/_0_  (.A1(\V2/V1/v4 [4]),
    .A2(\V2/V1/c3 ),
    .ZN(\V2/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M1/M1/_1_  (.A(\V2/V1/v4 [4]),
    .B(\V2/V1/c3 ),
    .Z(\V2/V1/A3/A2/M1/s1 ));
 AND2_X1 \V2/V1/A3/A2/M1/M2/_0_  (.A1(\V2/V1/A3/A2/M1/s1 ),
    .A2(\V2/V1/A3/c1 ),
    .ZN(\V2/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M1/M2/_1_  (.A(\V2/V1/A3/A2/M1/s1 ),
    .B(\V2/V1/A3/c1 ),
    .Z(\V2/v1 [12]));
 OR2_X1 \V2/V1/A3/A2/M1/_0_  (.A1(\V2/V1/A3/A2/M1/c1 ),
    .A2(\V2/V1/A3/A2/M1/c2 ),
    .ZN(\V2/V1/A3/A2/c1 ));
 AND2_X1 \V2/V1/A3/A2/M2/M1/_0_  (.A1(\V2/V1/v4 [5]),
    .A2(ground),
    .ZN(\V2/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M2/M1/_1_  (.A(\V2/V1/v4 [5]),
    .B(ground),
    .Z(\V2/V1/A3/A2/M2/s1 ));
 AND2_X1 \V2/V1/A3/A2/M2/M2/_0_  (.A1(\V2/V1/A3/A2/M2/s1 ),
    .A2(\V2/V1/A3/A2/c1 ),
    .ZN(\V2/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M2/M2/_1_  (.A(\V2/V1/A3/A2/M2/s1 ),
    .B(\V2/V1/A3/A2/c1 ),
    .Z(\V2/v1 [13]));
 OR2_X1 \V2/V1/A3/A2/M2/_0_  (.A1(\V2/V1/A3/A2/M2/c1 ),
    .A2(\V2/V1/A3/A2/M2/c2 ),
    .ZN(\V2/V1/A3/A2/c2 ));
 AND2_X1 \V2/V1/A3/A2/M3/M1/_0_  (.A1(\V2/V1/v4 [6]),
    .A2(ground),
    .ZN(\V2/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M3/M1/_1_  (.A(\V2/V1/v4 [6]),
    .B(ground),
    .Z(\V2/V1/A3/A2/M3/s1 ));
 AND2_X1 \V2/V1/A3/A2/M3/M2/_0_  (.A1(\V2/V1/A3/A2/M3/s1 ),
    .A2(\V2/V1/A3/A2/c2 ),
    .ZN(\V2/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M3/M2/_1_  (.A(\V2/V1/A3/A2/M3/s1 ),
    .B(\V2/V1/A3/A2/c2 ),
    .Z(\V2/v1 [14]));
 OR2_X1 \V2/V1/A3/A2/M3/_0_  (.A1(\V2/V1/A3/A2/M3/c1 ),
    .A2(\V2/V1/A3/A2/M3/c2 ),
    .ZN(\V2/V1/A3/A2/c3 ));
 AND2_X1 \V2/V1/A3/A2/M4/M1/_0_  (.A1(\V2/V1/v4 [7]),
    .A2(ground),
    .ZN(\V2/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M4/M1/_1_  (.A(\V2/V1/v4 [7]),
    .B(ground),
    .Z(\V2/V1/A3/A2/M4/s1 ));
 AND2_X1 \V2/V1/A3/A2/M4/M2/_0_  (.A1(\V2/V1/A3/A2/M4/s1 ),
    .A2(\V2/V1/A3/A2/c3 ),
    .ZN(\V2/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M4/M2/_1_  (.A(\V2/V1/A3/A2/M4/s1 ),
    .B(\V2/V1/A3/A2/c3 ),
    .Z(\V2/v1 [15]));
 OR2_X1 \V2/V1/A3/A2/M4/_0_  (.A1(\V2/V1/A3/A2/M4/c1 ),
    .A2(\V2/V1/A3/A2/M4/c2 ),
    .ZN(\V2/V1/overflow ));
 AND2_X1 \V2/V1/V1/A1/M1/M1/_0_  (.A1(\V2/V1/V1/v2 [0]),
    .A2(\V2/V1/V1/v3 [0]),
    .ZN(\V2/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M1/M1/_1_  (.A(\V2/V1/V1/v2 [0]),
    .B(\V2/V1/V1/v3 [0]),
    .Z(\V2/V1/V1/A1/M1/s1 ));
 AND2_X1 \V2/V1/V1/A1/M1/M2/_0_  (.A1(\V2/V1/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M1/M2/_1_  (.A(\V2/V1/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/V1/s1 [0]));
 OR2_X1 \V2/V1/V1/A1/M1/_0_  (.A1(\V2/V1/V1/A1/M1/c1 ),
    .A2(\V2/V1/V1/A1/M1/c2 ),
    .ZN(\V2/V1/V1/A1/c1 ));
 AND2_X1 \V2/V1/V1/A1/M2/M1/_0_  (.A1(\V2/V1/V1/v2 [1]),
    .A2(\V2/V1/V1/v3 [1]),
    .ZN(\V2/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M2/M1/_1_  (.A(\V2/V1/V1/v2 [1]),
    .B(\V2/V1/V1/v3 [1]),
    .Z(\V2/V1/V1/A1/M2/s1 ));
 AND2_X1 \V2/V1/V1/A1/M2/M2/_0_  (.A1(\V2/V1/V1/A1/M2/s1 ),
    .A2(\V2/V1/V1/A1/c1 ),
    .ZN(\V2/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M2/M2/_1_  (.A(\V2/V1/V1/A1/M2/s1 ),
    .B(\V2/V1/V1/A1/c1 ),
    .Z(\V2/V1/V1/s1 [1]));
 OR2_X1 \V2/V1/V1/A1/M2/_0_  (.A1(\V2/V1/V1/A1/M2/c1 ),
    .A2(\V2/V1/V1/A1/M2/c2 ),
    .ZN(\V2/V1/V1/A1/c2 ));
 AND2_X1 \V2/V1/V1/A1/M3/M1/_0_  (.A1(\V2/V1/V1/v2 [2]),
    .A2(\V2/V1/V1/v3 [2]),
    .ZN(\V2/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M3/M1/_1_  (.A(\V2/V1/V1/v2 [2]),
    .B(\V2/V1/V1/v3 [2]),
    .Z(\V2/V1/V1/A1/M3/s1 ));
 AND2_X1 \V2/V1/V1/A1/M3/M2/_0_  (.A1(\V2/V1/V1/A1/M3/s1 ),
    .A2(\V2/V1/V1/A1/c2 ),
    .ZN(\V2/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M3/M2/_1_  (.A(\V2/V1/V1/A1/M3/s1 ),
    .B(\V2/V1/V1/A1/c2 ),
    .Z(\V2/V1/V1/s1 [2]));
 OR2_X1 \V2/V1/V1/A1/M3/_0_  (.A1(\V2/V1/V1/A1/M3/c1 ),
    .A2(\V2/V1/V1/A1/M3/c2 ),
    .ZN(\V2/V1/V1/A1/c3 ));
 AND2_X1 \V2/V1/V1/A1/M4/M1/_0_  (.A1(\V2/V1/V1/v2 [3]),
    .A2(\V2/V1/V1/v3 [3]),
    .ZN(\V2/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M4/M1/_1_  (.A(\V2/V1/V1/v2 [3]),
    .B(\V2/V1/V1/v3 [3]),
    .Z(\V2/V1/V1/A1/M4/s1 ));
 AND2_X1 \V2/V1/V1/A1/M4/M2/_0_  (.A1(\V2/V1/V1/A1/M4/s1 ),
    .A2(\V2/V1/V1/A1/c3 ),
    .ZN(\V2/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M4/M2/_1_  (.A(\V2/V1/V1/A1/M4/s1 ),
    .B(\V2/V1/V1/A1/c3 ),
    .Z(\V2/V1/V1/s1 [3]));
 OR2_X1 \V2/V1/V1/A1/M4/_0_  (.A1(\V2/V1/V1/A1/M4/c1 ),
    .A2(\V2/V1/V1/A1/M4/c2 ),
    .ZN(\V2/V1/V1/c1 ));
 AND2_X1 \V2/V1/V1/A2/M1/M1/_0_  (.A1(\V2/V1/V1/s1 [0]),
    .A2(\V2/V1/V1/v1 [2]),
    .ZN(\V2/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M1/M1/_1_  (.A(\V2/V1/V1/s1 [0]),
    .B(\V2/V1/V1/v1 [2]),
    .Z(\V2/V1/V1/A2/M1/s1 ));
 AND2_X1 \V2/V1/V1/A2/M1/M2/_0_  (.A1(\V2/V1/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M1/M2/_1_  (.A(\V2/V1/V1/A2/M1/s1 ),
    .B(ground),
    .Z(v2[2]));
 OR2_X1 \V2/V1/V1/A2/M1/_0_  (.A1(\V2/V1/V1/A2/M1/c1 ),
    .A2(\V2/V1/V1/A2/M1/c2 ),
    .ZN(\V2/V1/V1/A2/c1 ));
 AND2_X1 \V2/V1/V1/A2/M2/M1/_0_  (.A1(\V2/V1/V1/s1 [1]),
    .A2(\V2/V1/V1/v1 [3]),
    .ZN(\V2/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M2/M1/_1_  (.A(\V2/V1/V1/s1 [1]),
    .B(\V2/V1/V1/v1 [3]),
    .Z(\V2/V1/V1/A2/M2/s1 ));
 AND2_X1 \V2/V1/V1/A2/M2/M2/_0_  (.A1(\V2/V1/V1/A2/M2/s1 ),
    .A2(\V2/V1/V1/A2/c1 ),
    .ZN(\V2/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M2/M2/_1_  (.A(\V2/V1/V1/A2/M2/s1 ),
    .B(\V2/V1/V1/A2/c1 ),
    .Z(v2[3]));
 OR2_X1 \V2/V1/V1/A2/M2/_0_  (.A1(\V2/V1/V1/A2/M2/c1 ),
    .A2(\V2/V1/V1/A2/M2/c2 ),
    .ZN(\V2/V1/V1/A2/c2 ));
 AND2_X1 \V2/V1/V1/A2/M3/M1/_0_  (.A1(\V2/V1/V1/s1 [2]),
    .A2(ground),
    .ZN(\V2/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M3/M1/_1_  (.A(\V2/V1/V1/s1 [2]),
    .B(ground),
    .Z(\V2/V1/V1/A2/M3/s1 ));
 AND2_X1 \V2/V1/V1/A2/M3/M2/_0_  (.A1(\V2/V1/V1/A2/M3/s1 ),
    .A2(\V2/V1/V1/A2/c2 ),
    .ZN(\V2/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M3/M2/_1_  (.A(\V2/V1/V1/A2/M3/s1 ),
    .B(\V2/V1/V1/A2/c2 ),
    .Z(\V2/V1/V1/s2 [2]));
 OR2_X1 \V2/V1/V1/A2/M3/_0_  (.A1(\V2/V1/V1/A2/M3/c1 ),
    .A2(\V2/V1/V1/A2/M3/c2 ),
    .ZN(\V2/V1/V1/A2/c3 ));
 AND2_X1 \V2/V1/V1/A2/M4/M1/_0_  (.A1(\V2/V1/V1/s1 [3]),
    .A2(ground),
    .ZN(\V2/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M4/M1/_1_  (.A(\V2/V1/V1/s1 [3]),
    .B(ground),
    .Z(\V2/V1/V1/A2/M4/s1 ));
 AND2_X1 \V2/V1/V1/A2/M4/M2/_0_  (.A1(\V2/V1/V1/A2/M4/s1 ),
    .A2(\V2/V1/V1/A2/c3 ),
    .ZN(\V2/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M4/M2/_1_  (.A(\V2/V1/V1/A2/M4/s1 ),
    .B(\V2/V1/V1/A2/c3 ),
    .Z(\V2/V1/V1/s2 [3]));
 OR2_X1 \V2/V1/V1/A2/M4/_0_  (.A1(\V2/V1/V1/A2/M4/c1 ),
    .A2(\V2/V1/V1/A2/M4/c2 ),
    .ZN(\V2/V1/V1/c2 ));
 AND2_X1 \V2/V1/V1/A3/M1/M1/_0_  (.A1(\V2/V1/V1/v4 [0]),
    .A2(\V2/V1/V1/s2 [2]),
    .ZN(\V2/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M1/M1/_1_  (.A(\V2/V1/V1/v4 [0]),
    .B(\V2/V1/V1/s2 [2]),
    .Z(\V2/V1/V1/A3/M1/s1 ));
 AND2_X1 \V2/V1/V1/A3/M1/M2/_0_  (.A1(\V2/V1/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M1/M2/_1_  (.A(\V2/V1/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v1 [4]));
 OR2_X1 \V2/V1/V1/A3/M1/_0_  (.A1(\V2/V1/V1/A3/M1/c1 ),
    .A2(\V2/V1/V1/A3/M1/c2 ),
    .ZN(\V2/V1/V1/A3/c1 ));
 AND2_X1 \V2/V1/V1/A3/M2/M1/_0_  (.A1(\V2/V1/V1/v4 [1]),
    .A2(\V2/V1/V1/s2 [3]),
    .ZN(\V2/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M2/M1/_1_  (.A(\V2/V1/V1/v4 [1]),
    .B(\V2/V1/V1/s2 [3]),
    .Z(\V2/V1/V1/A3/M2/s1 ));
 AND2_X1 \V2/V1/V1/A3/M2/M2/_0_  (.A1(\V2/V1/V1/A3/M2/s1 ),
    .A2(\V2/V1/V1/A3/c1 ),
    .ZN(\V2/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M2/M2/_1_  (.A(\V2/V1/V1/A3/M2/s1 ),
    .B(\V2/V1/V1/A3/c1 ),
    .Z(\V2/V1/v1 [5]));
 OR2_X1 \V2/V1/V1/A3/M2/_0_  (.A1(\V2/V1/V1/A3/M2/c1 ),
    .A2(\V2/V1/V1/A3/M2/c2 ),
    .ZN(\V2/V1/V1/A3/c2 ));
 AND2_X1 \V2/V1/V1/A3/M3/M1/_0_  (.A1(\V2/V1/V1/v4 [2]),
    .A2(\V2/V1/V1/c3 ),
    .ZN(\V2/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M3/M1/_1_  (.A(\V2/V1/V1/v4 [2]),
    .B(\V2/V1/V1/c3 ),
    .Z(\V2/V1/V1/A3/M3/s1 ));
 AND2_X1 \V2/V1/V1/A3/M3/M2/_0_  (.A1(\V2/V1/V1/A3/M3/s1 ),
    .A2(\V2/V1/V1/A3/c2 ),
    .ZN(\V2/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M3/M2/_1_  (.A(\V2/V1/V1/A3/M3/s1 ),
    .B(\V2/V1/V1/A3/c2 ),
    .Z(\V2/V1/v1 [6]));
 OR2_X1 \V2/V1/V1/A3/M3/_0_  (.A1(\V2/V1/V1/A3/M3/c1 ),
    .A2(\V2/V1/V1/A3/M3/c2 ),
    .ZN(\V2/V1/V1/A3/c3 ));
 AND2_X1 \V2/V1/V1/A3/M4/M1/_0_  (.A1(\V2/V1/V1/v4 [3]),
    .A2(ground),
    .ZN(\V2/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M4/M1/_1_  (.A(\V2/V1/V1/v4 [3]),
    .B(ground),
    .Z(\V2/V1/V1/A3/M4/s1 ));
 AND2_X1 \V2/V1/V1/A3/M4/M2/_0_  (.A1(\V2/V1/V1/A3/M4/s1 ),
    .A2(\V2/V1/V1/A3/c3 ),
    .ZN(\V2/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M4/M2/_1_  (.A(\V2/V1/V1/A3/M4/s1 ),
    .B(\V2/V1/V1/A3/c3 ),
    .Z(\V2/V1/v1 [7]));
 OR2_X1 \V2/V1/V1/A3/M4/_0_  (.A1(\V2/V1/V1/A3/M4/c1 ),
    .A2(\V2/V1/V1/A3/M4/c2 ),
    .ZN(\V2/V1/V1/overflow ));
 AND2_X1 \V2/V1/V1/V1/HA1/_0_  (.A1(\V2/V1/V1/V1/w2 ),
    .A2(\V2/V1/V1/V1/w1 ),
    .ZN(\V2/V1/V1/V1/w4 ));
 XOR2_X2 \V2/V1/V1/V1/HA1/_1_  (.A(\V2/V1/V1/V1/w2 ),
    .B(\V2/V1/V1/V1/w1 ),
    .Z(v2[1]));
 AND2_X1 \V2/V1/V1/V1/HA2/_0_  (.A1(\V2/V1/V1/V1/w4 ),
    .A2(\V2/V1/V1/V1/w3 ),
    .ZN(\V2/V1/V1/v1 [3]));
 XOR2_X2 \V2/V1/V1/V1/HA2/_1_  (.A(\V2/V1/V1/V1/w4 ),
    .B(\V2/V1/V1/V1/w3 ),
    .Z(\V2/V1/V1/v1 [2]));
 AND2_X1 \V2/V1/V1/V1/_0_  (.A1(A[16]),
    .A2(B[0]),
    .ZN(v2[0]));
 AND2_X1 \V2/V1/V1/V1/_1_  (.A1(A[16]),
    .A2(B[1]),
    .ZN(\V2/V1/V1/V1/w1 ));
 AND2_X1 \V2/V1/V1/V1/_2_  (.A1(B[0]),
    .A2(A[17]),
    .ZN(\V2/V1/V1/V1/w2 ));
 AND2_X1 \V2/V1/V1/V1/_3_  (.A1(B[1]),
    .A2(A[17]),
    .ZN(\V2/V1/V1/V1/w3 ));
 AND2_X1 \V2/V1/V1/V2/HA1/_0_  (.A1(\V2/V1/V1/V2/w2 ),
    .A2(\V2/V1/V1/V2/w1 ),
    .ZN(\V2/V1/V1/V2/w4 ));
 XOR2_X2 \V2/V1/V1/V2/HA1/_1_  (.A(\V2/V1/V1/V2/w2 ),
    .B(\V2/V1/V1/V2/w1 ),
    .Z(\V2/V1/V1/v2 [1]));
 AND2_X1 \V2/V1/V1/V2/HA2/_0_  (.A1(\V2/V1/V1/V2/w4 ),
    .A2(\V2/V1/V1/V2/w3 ),
    .ZN(\V2/V1/V1/v2 [3]));
 XOR2_X2 \V2/V1/V1/V2/HA2/_1_  (.A(\V2/V1/V1/V2/w4 ),
    .B(\V2/V1/V1/V2/w3 ),
    .Z(\V2/V1/V1/v2 [2]));
 AND2_X1 \V2/V1/V1/V2/_0_  (.A1(A[18]),
    .A2(B[0]),
    .ZN(\V2/V1/V1/v2 [0]));
 AND2_X1 \V2/V1/V1/V2/_1_  (.A1(A[18]),
    .A2(B[1]),
    .ZN(\V2/V1/V1/V2/w1 ));
 AND2_X1 \V2/V1/V1/V2/_2_  (.A1(B[0]),
    .A2(A[19]),
    .ZN(\V2/V1/V1/V2/w2 ));
 AND2_X1 \V2/V1/V1/V2/_3_  (.A1(B[1]),
    .A2(A[19]),
    .ZN(\V2/V1/V1/V2/w3 ));
 AND2_X1 \V2/V1/V1/V3/HA1/_0_  (.A1(\V2/V1/V1/V3/w2 ),
    .A2(\V2/V1/V1/V3/w1 ),
    .ZN(\V2/V1/V1/V3/w4 ));
 XOR2_X2 \V2/V1/V1/V3/HA1/_1_  (.A(\V2/V1/V1/V3/w2 ),
    .B(\V2/V1/V1/V3/w1 ),
    .Z(\V2/V1/V1/v3 [1]));
 AND2_X1 \V2/V1/V1/V3/HA2/_0_  (.A1(\V2/V1/V1/V3/w4 ),
    .A2(\V2/V1/V1/V3/w3 ),
    .ZN(\V2/V1/V1/v3 [3]));
 XOR2_X2 \V2/V1/V1/V3/HA2/_1_  (.A(\V2/V1/V1/V3/w4 ),
    .B(\V2/V1/V1/V3/w3 ),
    .Z(\V2/V1/V1/v3 [2]));
 AND2_X1 \V2/V1/V1/V3/_0_  (.A1(A[16]),
    .A2(B[2]),
    .ZN(\V2/V1/V1/v3 [0]));
 AND2_X1 \V2/V1/V1/V3/_1_  (.A1(A[16]),
    .A2(B[3]),
    .ZN(\V2/V1/V1/V3/w1 ));
 AND2_X1 \V2/V1/V1/V3/_2_  (.A1(B[2]),
    .A2(A[17]),
    .ZN(\V2/V1/V1/V3/w2 ));
 AND2_X1 \V2/V1/V1/V3/_3_  (.A1(B[3]),
    .A2(A[17]),
    .ZN(\V2/V1/V1/V3/w3 ));
 AND2_X1 \V2/V1/V1/V4/HA1/_0_  (.A1(\V2/V1/V1/V4/w2 ),
    .A2(\V2/V1/V1/V4/w1 ),
    .ZN(\V2/V1/V1/V4/w4 ));
 XOR2_X2 \V2/V1/V1/V4/HA1/_1_  (.A(\V2/V1/V1/V4/w2 ),
    .B(\V2/V1/V1/V4/w1 ),
    .Z(\V2/V1/V1/v4 [1]));
 AND2_X1 \V2/V1/V1/V4/HA2/_0_  (.A1(\V2/V1/V1/V4/w4 ),
    .A2(\V2/V1/V1/V4/w3 ),
    .ZN(\V2/V1/V1/v4 [3]));
 XOR2_X2 \V2/V1/V1/V4/HA2/_1_  (.A(\V2/V1/V1/V4/w4 ),
    .B(\V2/V1/V1/V4/w3 ),
    .Z(\V2/V1/V1/v4 [2]));
 AND2_X1 \V2/V1/V1/V4/_0_  (.A1(A[18]),
    .A2(B[2]),
    .ZN(\V2/V1/V1/v4 [0]));
 AND2_X1 \V2/V1/V1/V4/_1_  (.A1(A[18]),
    .A2(B[3]),
    .ZN(\V2/V1/V1/V4/w1 ));
 AND2_X1 \V2/V1/V1/V4/_2_  (.A1(B[2]),
    .A2(A[19]),
    .ZN(\V2/V1/V1/V4/w2 ));
 AND2_X1 \V2/V1/V1/V4/_3_  (.A1(B[3]),
    .A2(A[19]),
    .ZN(\V2/V1/V1/V4/w3 ));
 OR2_X1 \V2/V1/V1/_0_  (.A1(\V2/V1/V1/c1 ),
    .A2(\V2/V1/V1/c2 ),
    .ZN(\V2/V1/V1/c3 ));
 AND2_X1 \V2/V1/V2/A1/M1/M1/_0_  (.A1(\V2/V1/V2/v2 [0]),
    .A2(\V2/V1/V2/v3 [0]),
    .ZN(\V2/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M1/M1/_1_  (.A(\V2/V1/V2/v2 [0]),
    .B(\V2/V1/V2/v3 [0]),
    .Z(\V2/V1/V2/A1/M1/s1 ));
 AND2_X1 \V2/V1/V2/A1/M1/M2/_0_  (.A1(\V2/V1/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M1/M2/_1_  (.A(\V2/V1/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/V2/s1 [0]));
 OR2_X1 \V2/V1/V2/A1/M1/_0_  (.A1(\V2/V1/V2/A1/M1/c1 ),
    .A2(\V2/V1/V2/A1/M1/c2 ),
    .ZN(\V2/V1/V2/A1/c1 ));
 AND2_X1 \V2/V1/V2/A1/M2/M1/_0_  (.A1(\V2/V1/V2/v2 [1]),
    .A2(\V2/V1/V2/v3 [1]),
    .ZN(\V2/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M2/M1/_1_  (.A(\V2/V1/V2/v2 [1]),
    .B(\V2/V1/V2/v3 [1]),
    .Z(\V2/V1/V2/A1/M2/s1 ));
 AND2_X1 \V2/V1/V2/A1/M2/M2/_0_  (.A1(\V2/V1/V2/A1/M2/s1 ),
    .A2(\V2/V1/V2/A1/c1 ),
    .ZN(\V2/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M2/M2/_1_  (.A(\V2/V1/V2/A1/M2/s1 ),
    .B(\V2/V1/V2/A1/c1 ),
    .Z(\V2/V1/V2/s1 [1]));
 OR2_X1 \V2/V1/V2/A1/M2/_0_  (.A1(\V2/V1/V2/A1/M2/c1 ),
    .A2(\V2/V1/V2/A1/M2/c2 ),
    .ZN(\V2/V1/V2/A1/c2 ));
 AND2_X1 \V2/V1/V2/A1/M3/M1/_0_  (.A1(\V2/V1/V2/v2 [2]),
    .A2(\V2/V1/V2/v3 [2]),
    .ZN(\V2/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M3/M1/_1_  (.A(\V2/V1/V2/v2 [2]),
    .B(\V2/V1/V2/v3 [2]),
    .Z(\V2/V1/V2/A1/M3/s1 ));
 AND2_X1 \V2/V1/V2/A1/M3/M2/_0_  (.A1(\V2/V1/V2/A1/M3/s1 ),
    .A2(\V2/V1/V2/A1/c2 ),
    .ZN(\V2/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M3/M2/_1_  (.A(\V2/V1/V2/A1/M3/s1 ),
    .B(\V2/V1/V2/A1/c2 ),
    .Z(\V2/V1/V2/s1 [2]));
 OR2_X1 \V2/V1/V2/A1/M3/_0_  (.A1(\V2/V1/V2/A1/M3/c1 ),
    .A2(\V2/V1/V2/A1/M3/c2 ),
    .ZN(\V2/V1/V2/A1/c3 ));
 AND2_X1 \V2/V1/V2/A1/M4/M1/_0_  (.A1(\V2/V1/V2/v2 [3]),
    .A2(\V2/V1/V2/v3 [3]),
    .ZN(\V2/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M4/M1/_1_  (.A(\V2/V1/V2/v2 [3]),
    .B(\V2/V1/V2/v3 [3]),
    .Z(\V2/V1/V2/A1/M4/s1 ));
 AND2_X1 \V2/V1/V2/A1/M4/M2/_0_  (.A1(\V2/V1/V2/A1/M4/s1 ),
    .A2(\V2/V1/V2/A1/c3 ),
    .ZN(\V2/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M4/M2/_1_  (.A(\V2/V1/V2/A1/M4/s1 ),
    .B(\V2/V1/V2/A1/c3 ),
    .Z(\V2/V1/V2/s1 [3]));
 OR2_X1 \V2/V1/V2/A1/M4/_0_  (.A1(\V2/V1/V2/A1/M4/c1 ),
    .A2(\V2/V1/V2/A1/M4/c2 ),
    .ZN(\V2/V1/V2/c1 ));
 AND2_X1 \V2/V1/V2/A2/M1/M1/_0_  (.A1(\V2/V1/V2/s1 [0]),
    .A2(\V2/V1/V2/v1 [2]),
    .ZN(\V2/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M1/M1/_1_  (.A(\V2/V1/V2/s1 [0]),
    .B(\V2/V1/V2/v1 [2]),
    .Z(\V2/V1/V2/A2/M1/s1 ));
 AND2_X1 \V2/V1/V2/A2/M1/M2/_0_  (.A1(\V2/V1/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M1/M2/_1_  (.A(\V2/V1/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v2 [2]));
 OR2_X1 \V2/V1/V2/A2/M1/_0_  (.A1(\V2/V1/V2/A2/M1/c1 ),
    .A2(\V2/V1/V2/A2/M1/c2 ),
    .ZN(\V2/V1/V2/A2/c1 ));
 AND2_X1 \V2/V1/V2/A2/M2/M1/_0_  (.A1(\V2/V1/V2/s1 [1]),
    .A2(\V2/V1/V2/v1 [3]),
    .ZN(\V2/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M2/M1/_1_  (.A(\V2/V1/V2/s1 [1]),
    .B(\V2/V1/V2/v1 [3]),
    .Z(\V2/V1/V2/A2/M2/s1 ));
 AND2_X1 \V2/V1/V2/A2/M2/M2/_0_  (.A1(\V2/V1/V2/A2/M2/s1 ),
    .A2(\V2/V1/V2/A2/c1 ),
    .ZN(\V2/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M2/M2/_1_  (.A(\V2/V1/V2/A2/M2/s1 ),
    .B(\V2/V1/V2/A2/c1 ),
    .Z(\V2/V1/v2 [3]));
 OR2_X1 \V2/V1/V2/A2/M2/_0_  (.A1(\V2/V1/V2/A2/M2/c1 ),
    .A2(\V2/V1/V2/A2/M2/c2 ),
    .ZN(\V2/V1/V2/A2/c2 ));
 AND2_X1 \V2/V1/V2/A2/M3/M1/_0_  (.A1(\V2/V1/V2/s1 [2]),
    .A2(ground),
    .ZN(\V2/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M3/M1/_1_  (.A(\V2/V1/V2/s1 [2]),
    .B(ground),
    .Z(\V2/V1/V2/A2/M3/s1 ));
 AND2_X1 \V2/V1/V2/A2/M3/M2/_0_  (.A1(\V2/V1/V2/A2/M3/s1 ),
    .A2(\V2/V1/V2/A2/c2 ),
    .ZN(\V2/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M3/M2/_1_  (.A(\V2/V1/V2/A2/M3/s1 ),
    .B(\V2/V1/V2/A2/c2 ),
    .Z(\V2/V1/V2/s2 [2]));
 OR2_X1 \V2/V1/V2/A2/M3/_0_  (.A1(\V2/V1/V2/A2/M3/c1 ),
    .A2(\V2/V1/V2/A2/M3/c2 ),
    .ZN(\V2/V1/V2/A2/c3 ));
 AND2_X1 \V2/V1/V2/A2/M4/M1/_0_  (.A1(\V2/V1/V2/s1 [3]),
    .A2(ground),
    .ZN(\V2/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M4/M1/_1_  (.A(\V2/V1/V2/s1 [3]),
    .B(ground),
    .Z(\V2/V1/V2/A2/M4/s1 ));
 AND2_X1 \V2/V1/V2/A2/M4/M2/_0_  (.A1(\V2/V1/V2/A2/M4/s1 ),
    .A2(\V2/V1/V2/A2/c3 ),
    .ZN(\V2/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M4/M2/_1_  (.A(\V2/V1/V2/A2/M4/s1 ),
    .B(\V2/V1/V2/A2/c3 ),
    .Z(\V2/V1/V2/s2 [3]));
 OR2_X1 \V2/V1/V2/A2/M4/_0_  (.A1(\V2/V1/V2/A2/M4/c1 ),
    .A2(\V2/V1/V2/A2/M4/c2 ),
    .ZN(\V2/V1/V2/c2 ));
 AND2_X1 \V2/V1/V2/A3/M1/M1/_0_  (.A1(\V2/V1/V2/v4 [0]),
    .A2(\V2/V1/V2/s2 [2]),
    .ZN(\V2/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M1/M1/_1_  (.A(\V2/V1/V2/v4 [0]),
    .B(\V2/V1/V2/s2 [2]),
    .Z(\V2/V1/V2/A3/M1/s1 ));
 AND2_X1 \V2/V1/V2/A3/M1/M2/_0_  (.A1(\V2/V1/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M1/M2/_1_  (.A(\V2/V1/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v2 [4]));
 OR2_X1 \V2/V1/V2/A3/M1/_0_  (.A1(\V2/V1/V2/A3/M1/c1 ),
    .A2(\V2/V1/V2/A3/M1/c2 ),
    .ZN(\V2/V1/V2/A3/c1 ));
 AND2_X1 \V2/V1/V2/A3/M2/M1/_0_  (.A1(\V2/V1/V2/v4 [1]),
    .A2(\V2/V1/V2/s2 [3]),
    .ZN(\V2/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M2/M1/_1_  (.A(\V2/V1/V2/v4 [1]),
    .B(\V2/V1/V2/s2 [3]),
    .Z(\V2/V1/V2/A3/M2/s1 ));
 AND2_X1 \V2/V1/V2/A3/M2/M2/_0_  (.A1(\V2/V1/V2/A3/M2/s1 ),
    .A2(\V2/V1/V2/A3/c1 ),
    .ZN(\V2/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M2/M2/_1_  (.A(\V2/V1/V2/A3/M2/s1 ),
    .B(\V2/V1/V2/A3/c1 ),
    .Z(\V2/V1/v2 [5]));
 OR2_X1 \V2/V1/V2/A3/M2/_0_  (.A1(\V2/V1/V2/A3/M2/c1 ),
    .A2(\V2/V1/V2/A3/M2/c2 ),
    .ZN(\V2/V1/V2/A3/c2 ));
 AND2_X1 \V2/V1/V2/A3/M3/M1/_0_  (.A1(\V2/V1/V2/v4 [2]),
    .A2(\V2/V1/V2/c3 ),
    .ZN(\V2/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M3/M1/_1_  (.A(\V2/V1/V2/v4 [2]),
    .B(\V2/V1/V2/c3 ),
    .Z(\V2/V1/V2/A3/M3/s1 ));
 AND2_X1 \V2/V1/V2/A3/M3/M2/_0_  (.A1(\V2/V1/V2/A3/M3/s1 ),
    .A2(\V2/V1/V2/A3/c2 ),
    .ZN(\V2/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M3/M2/_1_  (.A(\V2/V1/V2/A3/M3/s1 ),
    .B(\V2/V1/V2/A3/c2 ),
    .Z(\V2/V1/v2 [6]));
 OR2_X1 \V2/V1/V2/A3/M3/_0_  (.A1(\V2/V1/V2/A3/M3/c1 ),
    .A2(\V2/V1/V2/A3/M3/c2 ),
    .ZN(\V2/V1/V2/A3/c3 ));
 AND2_X1 \V2/V1/V2/A3/M4/M1/_0_  (.A1(\V2/V1/V2/v4 [3]),
    .A2(ground),
    .ZN(\V2/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M4/M1/_1_  (.A(\V2/V1/V2/v4 [3]),
    .B(ground),
    .Z(\V2/V1/V2/A3/M4/s1 ));
 AND2_X1 \V2/V1/V2/A3/M4/M2/_0_  (.A1(\V2/V1/V2/A3/M4/s1 ),
    .A2(\V2/V1/V2/A3/c3 ),
    .ZN(\V2/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M4/M2/_1_  (.A(\V2/V1/V2/A3/M4/s1 ),
    .B(\V2/V1/V2/A3/c3 ),
    .Z(\V2/V1/v2 [7]));
 OR2_X1 \V2/V1/V2/A3/M4/_0_  (.A1(\V2/V1/V2/A3/M4/c1 ),
    .A2(\V2/V1/V2/A3/M4/c2 ),
    .ZN(\V2/V1/V2/overflow ));
 AND2_X1 \V2/V1/V2/V1/HA1/_0_  (.A1(\V2/V1/V2/V1/w2 ),
    .A2(\V2/V1/V2/V1/w1 ),
    .ZN(\V2/V1/V2/V1/w4 ));
 XOR2_X2 \V2/V1/V2/V1/HA1/_1_  (.A(\V2/V1/V2/V1/w2 ),
    .B(\V2/V1/V2/V1/w1 ),
    .Z(\V2/V1/v2 [1]));
 AND2_X1 \V2/V1/V2/V1/HA2/_0_  (.A1(\V2/V1/V2/V1/w4 ),
    .A2(\V2/V1/V2/V1/w3 ),
    .ZN(\V2/V1/V2/v1 [3]));
 XOR2_X2 \V2/V1/V2/V1/HA2/_1_  (.A(\V2/V1/V2/V1/w4 ),
    .B(\V2/V1/V2/V1/w3 ),
    .Z(\V2/V1/V2/v1 [2]));
 AND2_X1 \V2/V1/V2/V1/_0_  (.A1(A[20]),
    .A2(B[0]),
    .ZN(\V2/V1/v2 [0]));
 AND2_X1 \V2/V1/V2/V1/_1_  (.A1(A[20]),
    .A2(B[1]),
    .ZN(\V2/V1/V2/V1/w1 ));
 AND2_X1 \V2/V1/V2/V1/_2_  (.A1(B[0]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V1/w2 ));
 AND2_X1 \V2/V1/V2/V1/_3_  (.A1(B[1]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V1/w3 ));
 AND2_X1 \V2/V1/V2/V2/HA1/_0_  (.A1(\V2/V1/V2/V2/w2 ),
    .A2(\V2/V1/V2/V2/w1 ),
    .ZN(\V2/V1/V2/V2/w4 ));
 XOR2_X2 \V2/V1/V2/V2/HA1/_1_  (.A(\V2/V1/V2/V2/w2 ),
    .B(\V2/V1/V2/V2/w1 ),
    .Z(\V2/V1/V2/v2 [1]));
 AND2_X1 \V2/V1/V2/V2/HA2/_0_  (.A1(\V2/V1/V2/V2/w4 ),
    .A2(\V2/V1/V2/V2/w3 ),
    .ZN(\V2/V1/V2/v2 [3]));
 XOR2_X2 \V2/V1/V2/V2/HA2/_1_  (.A(\V2/V1/V2/V2/w4 ),
    .B(\V2/V1/V2/V2/w3 ),
    .Z(\V2/V1/V2/v2 [2]));
 AND2_X1 \V2/V1/V2/V2/_0_  (.A1(A[22]),
    .A2(B[0]),
    .ZN(\V2/V1/V2/v2 [0]));
 AND2_X1 \V2/V1/V2/V2/_1_  (.A1(A[22]),
    .A2(B[1]),
    .ZN(\V2/V1/V2/V2/w1 ));
 AND2_X1 \V2/V1/V2/V2/_2_  (.A1(B[0]),
    .A2(A[23]),
    .ZN(\V2/V1/V2/V2/w2 ));
 AND2_X1 \V2/V1/V2/V2/_3_  (.A1(B[1]),
    .A2(A[23]),
    .ZN(\V2/V1/V2/V2/w3 ));
 AND2_X1 \V2/V1/V2/V3/HA1/_0_  (.A1(\V2/V1/V2/V3/w2 ),
    .A2(\V2/V1/V2/V3/w1 ),
    .ZN(\V2/V1/V2/V3/w4 ));
 XOR2_X2 \V2/V1/V2/V3/HA1/_1_  (.A(\V2/V1/V2/V3/w2 ),
    .B(\V2/V1/V2/V3/w1 ),
    .Z(\V2/V1/V2/v3 [1]));
 AND2_X1 \V2/V1/V2/V3/HA2/_0_  (.A1(\V2/V1/V2/V3/w4 ),
    .A2(\V2/V1/V2/V3/w3 ),
    .ZN(\V2/V1/V2/v3 [3]));
 XOR2_X2 \V2/V1/V2/V3/HA2/_1_  (.A(\V2/V1/V2/V3/w4 ),
    .B(\V2/V1/V2/V3/w3 ),
    .Z(\V2/V1/V2/v3 [2]));
 AND2_X1 \V2/V1/V2/V3/_0_  (.A1(A[20]),
    .A2(B[2]),
    .ZN(\V2/V1/V2/v3 [0]));
 AND2_X1 \V2/V1/V2/V3/_1_  (.A1(A[20]),
    .A2(B[3]),
    .ZN(\V2/V1/V2/V3/w1 ));
 AND2_X1 \V2/V1/V2/V3/_2_  (.A1(B[2]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V3/w2 ));
 AND2_X1 \V2/V1/V2/V3/_3_  (.A1(B[3]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V3/w3 ));
 AND2_X1 \V2/V1/V2/V4/HA1/_0_  (.A1(\V2/V1/V2/V4/w2 ),
    .A2(\V2/V1/V2/V4/w1 ),
    .ZN(\V2/V1/V2/V4/w4 ));
 XOR2_X2 \V2/V1/V2/V4/HA1/_1_  (.A(\V2/V1/V2/V4/w2 ),
    .B(\V2/V1/V2/V4/w1 ),
    .Z(\V2/V1/V2/v4 [1]));
 AND2_X1 \V2/V1/V2/V4/HA2/_0_  (.A1(\V2/V1/V2/V4/w4 ),
    .A2(\V2/V1/V2/V4/w3 ),
    .ZN(\V2/V1/V2/v4 [3]));
 XOR2_X2 \V2/V1/V2/V4/HA2/_1_  (.A(\V2/V1/V2/V4/w4 ),
    .B(\V2/V1/V2/V4/w3 ),
    .Z(\V2/V1/V2/v4 [2]));
 AND2_X1 \V2/V1/V2/V4/_0_  (.A1(A[22]),
    .A2(B[2]),
    .ZN(\V2/V1/V2/v4 [0]));
 AND2_X1 \V2/V1/V2/V4/_1_  (.A1(A[22]),
    .A2(B[3]),
    .ZN(\V2/V1/V2/V4/w1 ));
 AND2_X1 \V2/V1/V2/V4/_2_  (.A1(B[2]),
    .A2(A[23]),
    .ZN(\V2/V1/V2/V4/w2 ));
 AND2_X1 \V2/V1/V2/V4/_3_  (.A1(B[3]),
    .A2(A[23]),
    .ZN(\V2/V1/V2/V4/w3 ));
 OR2_X1 \V2/V1/V2/_0_  (.A1(\V2/V1/V2/c1 ),
    .A2(\V2/V1/V2/c2 ),
    .ZN(\V2/V1/V2/c3 ));
 AND2_X1 \V2/V1/V3/A1/M1/M1/_0_  (.A1(\V2/V1/V3/v2 [0]),
    .A2(\V2/V1/V3/v3 [0]),
    .ZN(\V2/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M1/M1/_1_  (.A(\V2/V1/V3/v2 [0]),
    .B(\V2/V1/V3/v3 [0]),
    .Z(\V2/V1/V3/A1/M1/s1 ));
 AND2_X1 \V2/V1/V3/A1/M1/M2/_0_  (.A1(\V2/V1/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M1/M2/_1_  (.A(\V2/V1/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/V3/s1 [0]));
 OR2_X1 \V2/V1/V3/A1/M1/_0_  (.A1(\V2/V1/V3/A1/M1/c1 ),
    .A2(\V2/V1/V3/A1/M1/c2 ),
    .ZN(\V2/V1/V3/A1/c1 ));
 AND2_X1 \V2/V1/V3/A1/M2/M1/_0_  (.A1(\V2/V1/V3/v2 [1]),
    .A2(\V2/V1/V3/v3 [1]),
    .ZN(\V2/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M2/M1/_1_  (.A(\V2/V1/V3/v2 [1]),
    .B(\V2/V1/V3/v3 [1]),
    .Z(\V2/V1/V3/A1/M2/s1 ));
 AND2_X1 \V2/V1/V3/A1/M2/M2/_0_  (.A1(\V2/V1/V3/A1/M2/s1 ),
    .A2(\V2/V1/V3/A1/c1 ),
    .ZN(\V2/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M2/M2/_1_  (.A(\V2/V1/V3/A1/M2/s1 ),
    .B(\V2/V1/V3/A1/c1 ),
    .Z(\V2/V1/V3/s1 [1]));
 OR2_X1 \V2/V1/V3/A1/M2/_0_  (.A1(\V2/V1/V3/A1/M2/c1 ),
    .A2(\V2/V1/V3/A1/M2/c2 ),
    .ZN(\V2/V1/V3/A1/c2 ));
 AND2_X1 \V2/V1/V3/A1/M3/M1/_0_  (.A1(\V2/V1/V3/v2 [2]),
    .A2(\V2/V1/V3/v3 [2]),
    .ZN(\V2/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M3/M1/_1_  (.A(\V2/V1/V3/v2 [2]),
    .B(\V2/V1/V3/v3 [2]),
    .Z(\V2/V1/V3/A1/M3/s1 ));
 AND2_X1 \V2/V1/V3/A1/M3/M2/_0_  (.A1(\V2/V1/V3/A1/M3/s1 ),
    .A2(\V2/V1/V3/A1/c2 ),
    .ZN(\V2/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M3/M2/_1_  (.A(\V2/V1/V3/A1/M3/s1 ),
    .B(\V2/V1/V3/A1/c2 ),
    .Z(\V2/V1/V3/s1 [2]));
 OR2_X1 \V2/V1/V3/A1/M3/_0_  (.A1(\V2/V1/V3/A1/M3/c1 ),
    .A2(\V2/V1/V3/A1/M3/c2 ),
    .ZN(\V2/V1/V3/A1/c3 ));
 AND2_X1 \V2/V1/V3/A1/M4/M1/_0_  (.A1(\V2/V1/V3/v2 [3]),
    .A2(\V2/V1/V3/v3 [3]),
    .ZN(\V2/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M4/M1/_1_  (.A(\V2/V1/V3/v2 [3]),
    .B(\V2/V1/V3/v3 [3]),
    .Z(\V2/V1/V3/A1/M4/s1 ));
 AND2_X1 \V2/V1/V3/A1/M4/M2/_0_  (.A1(\V2/V1/V3/A1/M4/s1 ),
    .A2(\V2/V1/V3/A1/c3 ),
    .ZN(\V2/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M4/M2/_1_  (.A(\V2/V1/V3/A1/M4/s1 ),
    .B(\V2/V1/V3/A1/c3 ),
    .Z(\V2/V1/V3/s1 [3]));
 OR2_X1 \V2/V1/V3/A1/M4/_0_  (.A1(\V2/V1/V3/A1/M4/c1 ),
    .A2(\V2/V1/V3/A1/M4/c2 ),
    .ZN(\V2/V1/V3/c1 ));
 AND2_X1 \V2/V1/V3/A2/M1/M1/_0_  (.A1(\V2/V1/V3/s1 [0]),
    .A2(\V2/V1/V3/v1 [2]),
    .ZN(\V2/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M1/M1/_1_  (.A(\V2/V1/V3/s1 [0]),
    .B(\V2/V1/V3/v1 [2]),
    .Z(\V2/V1/V3/A2/M1/s1 ));
 AND2_X1 \V2/V1/V3/A2/M1/M2/_0_  (.A1(\V2/V1/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M1/M2/_1_  (.A(\V2/V1/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v3 [2]));
 OR2_X1 \V2/V1/V3/A2/M1/_0_  (.A1(\V2/V1/V3/A2/M1/c1 ),
    .A2(\V2/V1/V3/A2/M1/c2 ),
    .ZN(\V2/V1/V3/A2/c1 ));
 AND2_X1 \V2/V1/V3/A2/M2/M1/_0_  (.A1(\V2/V1/V3/s1 [1]),
    .A2(\V2/V1/V3/v1 [3]),
    .ZN(\V2/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M2/M1/_1_  (.A(\V2/V1/V3/s1 [1]),
    .B(\V2/V1/V3/v1 [3]),
    .Z(\V2/V1/V3/A2/M2/s1 ));
 AND2_X1 \V2/V1/V3/A2/M2/M2/_0_  (.A1(\V2/V1/V3/A2/M2/s1 ),
    .A2(\V2/V1/V3/A2/c1 ),
    .ZN(\V2/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M2/M2/_1_  (.A(\V2/V1/V3/A2/M2/s1 ),
    .B(\V2/V1/V3/A2/c1 ),
    .Z(\V2/V1/v3 [3]));
 OR2_X1 \V2/V1/V3/A2/M2/_0_  (.A1(\V2/V1/V3/A2/M2/c1 ),
    .A2(\V2/V1/V3/A2/M2/c2 ),
    .ZN(\V2/V1/V3/A2/c2 ));
 AND2_X1 \V2/V1/V3/A2/M3/M1/_0_  (.A1(\V2/V1/V3/s1 [2]),
    .A2(ground),
    .ZN(\V2/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M3/M1/_1_  (.A(\V2/V1/V3/s1 [2]),
    .B(ground),
    .Z(\V2/V1/V3/A2/M3/s1 ));
 AND2_X1 \V2/V1/V3/A2/M3/M2/_0_  (.A1(\V2/V1/V3/A2/M3/s1 ),
    .A2(\V2/V1/V3/A2/c2 ),
    .ZN(\V2/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M3/M2/_1_  (.A(\V2/V1/V3/A2/M3/s1 ),
    .B(\V2/V1/V3/A2/c2 ),
    .Z(\V2/V1/V3/s2 [2]));
 OR2_X1 \V2/V1/V3/A2/M3/_0_  (.A1(\V2/V1/V3/A2/M3/c1 ),
    .A2(\V2/V1/V3/A2/M3/c2 ),
    .ZN(\V2/V1/V3/A2/c3 ));
 AND2_X1 \V2/V1/V3/A2/M4/M1/_0_  (.A1(\V2/V1/V3/s1 [3]),
    .A2(ground),
    .ZN(\V2/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M4/M1/_1_  (.A(\V2/V1/V3/s1 [3]),
    .B(ground),
    .Z(\V2/V1/V3/A2/M4/s1 ));
 AND2_X1 \V2/V1/V3/A2/M4/M2/_0_  (.A1(\V2/V1/V3/A2/M4/s1 ),
    .A2(\V2/V1/V3/A2/c3 ),
    .ZN(\V2/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M4/M2/_1_  (.A(\V2/V1/V3/A2/M4/s1 ),
    .B(\V2/V1/V3/A2/c3 ),
    .Z(\V2/V1/V3/s2 [3]));
 OR2_X1 \V2/V1/V3/A2/M4/_0_  (.A1(\V2/V1/V3/A2/M4/c1 ),
    .A2(\V2/V1/V3/A2/M4/c2 ),
    .ZN(\V2/V1/V3/c2 ));
 AND2_X1 \V2/V1/V3/A3/M1/M1/_0_  (.A1(\V2/V1/V3/v4 [0]),
    .A2(\V2/V1/V3/s2 [2]),
    .ZN(\V2/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M1/M1/_1_  (.A(\V2/V1/V3/v4 [0]),
    .B(\V2/V1/V3/s2 [2]),
    .Z(\V2/V1/V3/A3/M1/s1 ));
 AND2_X1 \V2/V1/V3/A3/M1/M2/_0_  (.A1(\V2/V1/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M1/M2/_1_  (.A(\V2/V1/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v3 [4]));
 OR2_X1 \V2/V1/V3/A3/M1/_0_  (.A1(\V2/V1/V3/A3/M1/c1 ),
    .A2(\V2/V1/V3/A3/M1/c2 ),
    .ZN(\V2/V1/V3/A3/c1 ));
 AND2_X1 \V2/V1/V3/A3/M2/M1/_0_  (.A1(\V2/V1/V3/v4 [1]),
    .A2(\V2/V1/V3/s2 [3]),
    .ZN(\V2/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M2/M1/_1_  (.A(\V2/V1/V3/v4 [1]),
    .B(\V2/V1/V3/s2 [3]),
    .Z(\V2/V1/V3/A3/M2/s1 ));
 AND2_X1 \V2/V1/V3/A3/M2/M2/_0_  (.A1(\V2/V1/V3/A3/M2/s1 ),
    .A2(\V2/V1/V3/A3/c1 ),
    .ZN(\V2/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M2/M2/_1_  (.A(\V2/V1/V3/A3/M2/s1 ),
    .B(\V2/V1/V3/A3/c1 ),
    .Z(\V2/V1/v3 [5]));
 OR2_X1 \V2/V1/V3/A3/M2/_0_  (.A1(\V2/V1/V3/A3/M2/c1 ),
    .A2(\V2/V1/V3/A3/M2/c2 ),
    .ZN(\V2/V1/V3/A3/c2 ));
 AND2_X1 \V2/V1/V3/A3/M3/M1/_0_  (.A1(\V2/V1/V3/v4 [2]),
    .A2(\V2/V1/V3/c3 ),
    .ZN(\V2/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M3/M1/_1_  (.A(\V2/V1/V3/v4 [2]),
    .B(\V2/V1/V3/c3 ),
    .Z(\V2/V1/V3/A3/M3/s1 ));
 AND2_X1 \V2/V1/V3/A3/M3/M2/_0_  (.A1(\V2/V1/V3/A3/M3/s1 ),
    .A2(\V2/V1/V3/A3/c2 ),
    .ZN(\V2/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M3/M2/_1_  (.A(\V2/V1/V3/A3/M3/s1 ),
    .B(\V2/V1/V3/A3/c2 ),
    .Z(\V2/V1/v3 [6]));
 OR2_X1 \V2/V1/V3/A3/M3/_0_  (.A1(\V2/V1/V3/A3/M3/c1 ),
    .A2(\V2/V1/V3/A3/M3/c2 ),
    .ZN(\V2/V1/V3/A3/c3 ));
 AND2_X1 \V2/V1/V3/A3/M4/M1/_0_  (.A1(\V2/V1/V3/v4 [3]),
    .A2(ground),
    .ZN(\V2/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M4/M1/_1_  (.A(\V2/V1/V3/v4 [3]),
    .B(ground),
    .Z(\V2/V1/V3/A3/M4/s1 ));
 AND2_X1 \V2/V1/V3/A3/M4/M2/_0_  (.A1(\V2/V1/V3/A3/M4/s1 ),
    .A2(\V2/V1/V3/A3/c3 ),
    .ZN(\V2/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M4/M2/_1_  (.A(\V2/V1/V3/A3/M4/s1 ),
    .B(\V2/V1/V3/A3/c3 ),
    .Z(\V2/V1/v3 [7]));
 OR2_X1 \V2/V1/V3/A3/M4/_0_  (.A1(\V2/V1/V3/A3/M4/c1 ),
    .A2(\V2/V1/V3/A3/M4/c2 ),
    .ZN(\V2/V1/V3/overflow ));
 AND2_X1 \V2/V1/V3/V1/HA1/_0_  (.A1(\V2/V1/V3/V1/w2 ),
    .A2(\V2/V1/V3/V1/w1 ),
    .ZN(\V2/V1/V3/V1/w4 ));
 XOR2_X2 \V2/V1/V3/V1/HA1/_1_  (.A(\V2/V1/V3/V1/w2 ),
    .B(\V2/V1/V3/V1/w1 ),
    .Z(\V2/V1/v3 [1]));
 AND2_X1 \V2/V1/V3/V1/HA2/_0_  (.A1(\V2/V1/V3/V1/w4 ),
    .A2(\V2/V1/V3/V1/w3 ),
    .ZN(\V2/V1/V3/v1 [3]));
 XOR2_X2 \V2/V1/V3/V1/HA2/_1_  (.A(\V2/V1/V3/V1/w4 ),
    .B(\V2/V1/V3/V1/w3 ),
    .Z(\V2/V1/V3/v1 [2]));
 AND2_X1 \V2/V1/V3/V1/_0_  (.A1(A[16]),
    .A2(B[4]),
    .ZN(\V2/V1/v3 [0]));
 AND2_X1 \V2/V1/V3/V1/_1_  (.A1(A[16]),
    .A2(B[5]),
    .ZN(\V2/V1/V3/V1/w1 ));
 AND2_X1 \V2/V1/V3/V1/_2_  (.A1(B[4]),
    .A2(A[17]),
    .ZN(\V2/V1/V3/V1/w2 ));
 AND2_X1 \V2/V1/V3/V1/_3_  (.A1(B[5]),
    .A2(A[17]),
    .ZN(\V2/V1/V3/V1/w3 ));
 AND2_X1 \V2/V1/V3/V2/HA1/_0_  (.A1(\V2/V1/V3/V2/w2 ),
    .A2(\V2/V1/V3/V2/w1 ),
    .ZN(\V2/V1/V3/V2/w4 ));
 XOR2_X2 \V2/V1/V3/V2/HA1/_1_  (.A(\V2/V1/V3/V2/w2 ),
    .B(\V2/V1/V3/V2/w1 ),
    .Z(\V2/V1/V3/v2 [1]));
 AND2_X1 \V2/V1/V3/V2/HA2/_0_  (.A1(\V2/V1/V3/V2/w4 ),
    .A2(\V2/V1/V3/V2/w3 ),
    .ZN(\V2/V1/V3/v2 [3]));
 XOR2_X2 \V2/V1/V3/V2/HA2/_1_  (.A(\V2/V1/V3/V2/w4 ),
    .B(\V2/V1/V3/V2/w3 ),
    .Z(\V2/V1/V3/v2 [2]));
 AND2_X1 \V2/V1/V3/V2/_0_  (.A1(A[18]),
    .A2(B[4]),
    .ZN(\V2/V1/V3/v2 [0]));
 AND2_X1 \V2/V1/V3/V2/_1_  (.A1(A[18]),
    .A2(B[5]),
    .ZN(\V2/V1/V3/V2/w1 ));
 AND2_X1 \V2/V1/V3/V2/_2_  (.A1(B[4]),
    .A2(A[19]),
    .ZN(\V2/V1/V3/V2/w2 ));
 AND2_X1 \V2/V1/V3/V2/_3_  (.A1(B[5]),
    .A2(A[19]),
    .ZN(\V2/V1/V3/V2/w3 ));
 AND2_X1 \V2/V1/V3/V3/HA1/_0_  (.A1(\V2/V1/V3/V3/w2 ),
    .A2(\V2/V1/V3/V3/w1 ),
    .ZN(\V2/V1/V3/V3/w4 ));
 XOR2_X2 \V2/V1/V3/V3/HA1/_1_  (.A(\V2/V1/V3/V3/w2 ),
    .B(\V2/V1/V3/V3/w1 ),
    .Z(\V2/V1/V3/v3 [1]));
 AND2_X1 \V2/V1/V3/V3/HA2/_0_  (.A1(\V2/V1/V3/V3/w4 ),
    .A2(\V2/V1/V3/V3/w3 ),
    .ZN(\V2/V1/V3/v3 [3]));
 XOR2_X2 \V2/V1/V3/V3/HA2/_1_  (.A(\V2/V1/V3/V3/w4 ),
    .B(\V2/V1/V3/V3/w3 ),
    .Z(\V2/V1/V3/v3 [2]));
 AND2_X1 \V2/V1/V3/V3/_0_  (.A1(A[16]),
    .A2(B[6]),
    .ZN(\V2/V1/V3/v3 [0]));
 AND2_X1 \V2/V1/V3/V3/_1_  (.A1(A[16]),
    .A2(B[7]),
    .ZN(\V2/V1/V3/V3/w1 ));
 AND2_X1 \V2/V1/V3/V3/_2_  (.A1(B[6]),
    .A2(A[17]),
    .ZN(\V2/V1/V3/V3/w2 ));
 AND2_X1 \V2/V1/V3/V3/_3_  (.A1(B[7]),
    .A2(A[17]),
    .ZN(\V2/V1/V3/V3/w3 ));
 AND2_X1 \V2/V1/V3/V4/HA1/_0_  (.A1(\V2/V1/V3/V4/w2 ),
    .A2(\V2/V1/V3/V4/w1 ),
    .ZN(\V2/V1/V3/V4/w4 ));
 XOR2_X2 \V2/V1/V3/V4/HA1/_1_  (.A(\V2/V1/V3/V4/w2 ),
    .B(\V2/V1/V3/V4/w1 ),
    .Z(\V2/V1/V3/v4 [1]));
 AND2_X1 \V2/V1/V3/V4/HA2/_0_  (.A1(\V2/V1/V3/V4/w4 ),
    .A2(\V2/V1/V3/V4/w3 ),
    .ZN(\V2/V1/V3/v4 [3]));
 XOR2_X2 \V2/V1/V3/V4/HA2/_1_  (.A(\V2/V1/V3/V4/w4 ),
    .B(\V2/V1/V3/V4/w3 ),
    .Z(\V2/V1/V3/v4 [2]));
 AND2_X1 \V2/V1/V3/V4/_0_  (.A1(A[18]),
    .A2(B[6]),
    .ZN(\V2/V1/V3/v4 [0]));
 AND2_X1 \V2/V1/V3/V4/_1_  (.A1(A[18]),
    .A2(B[7]),
    .ZN(\V2/V1/V3/V4/w1 ));
 AND2_X1 \V2/V1/V3/V4/_2_  (.A1(B[6]),
    .A2(A[19]),
    .ZN(\V2/V1/V3/V4/w2 ));
 AND2_X1 \V2/V1/V3/V4/_3_  (.A1(B[7]),
    .A2(A[19]),
    .ZN(\V2/V1/V3/V4/w3 ));
 OR2_X1 \V2/V1/V3/_0_  (.A1(\V2/V1/V3/c1 ),
    .A2(\V2/V1/V3/c2 ),
    .ZN(\V2/V1/V3/c3 ));
 AND2_X1 \V2/V1/V4/A1/M1/M1/_0_  (.A1(\V2/V1/V4/v2 [0]),
    .A2(\V2/V1/V4/v3 [0]),
    .ZN(\V2/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M1/M1/_1_  (.A(\V2/V1/V4/v2 [0]),
    .B(\V2/V1/V4/v3 [0]),
    .Z(\V2/V1/V4/A1/M1/s1 ));
 AND2_X1 \V2/V1/V4/A1/M1/M2/_0_  (.A1(\V2/V1/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M1/M2/_1_  (.A(\V2/V1/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/V4/s1 [0]));
 OR2_X1 \V2/V1/V4/A1/M1/_0_  (.A1(\V2/V1/V4/A1/M1/c1 ),
    .A2(\V2/V1/V4/A1/M1/c2 ),
    .ZN(\V2/V1/V4/A1/c1 ));
 AND2_X1 \V2/V1/V4/A1/M2/M1/_0_  (.A1(\V2/V1/V4/v2 [1]),
    .A2(\V2/V1/V4/v3 [1]),
    .ZN(\V2/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M2/M1/_1_  (.A(\V2/V1/V4/v2 [1]),
    .B(\V2/V1/V4/v3 [1]),
    .Z(\V2/V1/V4/A1/M2/s1 ));
 AND2_X1 \V2/V1/V4/A1/M2/M2/_0_  (.A1(\V2/V1/V4/A1/M2/s1 ),
    .A2(\V2/V1/V4/A1/c1 ),
    .ZN(\V2/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M2/M2/_1_  (.A(\V2/V1/V4/A1/M2/s1 ),
    .B(\V2/V1/V4/A1/c1 ),
    .Z(\V2/V1/V4/s1 [1]));
 OR2_X1 \V2/V1/V4/A1/M2/_0_  (.A1(\V2/V1/V4/A1/M2/c1 ),
    .A2(\V2/V1/V4/A1/M2/c2 ),
    .ZN(\V2/V1/V4/A1/c2 ));
 AND2_X1 \V2/V1/V4/A1/M3/M1/_0_  (.A1(\V2/V1/V4/v2 [2]),
    .A2(\V2/V1/V4/v3 [2]),
    .ZN(\V2/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M3/M1/_1_  (.A(\V2/V1/V4/v2 [2]),
    .B(\V2/V1/V4/v3 [2]),
    .Z(\V2/V1/V4/A1/M3/s1 ));
 AND2_X1 \V2/V1/V4/A1/M3/M2/_0_  (.A1(\V2/V1/V4/A1/M3/s1 ),
    .A2(\V2/V1/V4/A1/c2 ),
    .ZN(\V2/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M3/M2/_1_  (.A(\V2/V1/V4/A1/M3/s1 ),
    .B(\V2/V1/V4/A1/c2 ),
    .Z(\V2/V1/V4/s1 [2]));
 OR2_X1 \V2/V1/V4/A1/M3/_0_  (.A1(\V2/V1/V4/A1/M3/c1 ),
    .A2(\V2/V1/V4/A1/M3/c2 ),
    .ZN(\V2/V1/V4/A1/c3 ));
 AND2_X1 \V2/V1/V4/A1/M4/M1/_0_  (.A1(\V2/V1/V4/v2 [3]),
    .A2(\V2/V1/V4/v3 [3]),
    .ZN(\V2/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M4/M1/_1_  (.A(\V2/V1/V4/v2 [3]),
    .B(\V2/V1/V4/v3 [3]),
    .Z(\V2/V1/V4/A1/M4/s1 ));
 AND2_X1 \V2/V1/V4/A1/M4/M2/_0_  (.A1(\V2/V1/V4/A1/M4/s1 ),
    .A2(\V2/V1/V4/A1/c3 ),
    .ZN(\V2/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M4/M2/_1_  (.A(\V2/V1/V4/A1/M4/s1 ),
    .B(\V2/V1/V4/A1/c3 ),
    .Z(\V2/V1/V4/s1 [3]));
 OR2_X1 \V2/V1/V4/A1/M4/_0_  (.A1(\V2/V1/V4/A1/M4/c1 ),
    .A2(\V2/V1/V4/A1/M4/c2 ),
    .ZN(\V2/V1/V4/c1 ));
 AND2_X1 \V2/V1/V4/A2/M1/M1/_0_  (.A1(\V2/V1/V4/s1 [0]),
    .A2(\V2/V1/V4/v1 [2]),
    .ZN(\V2/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M1/M1/_1_  (.A(\V2/V1/V4/s1 [0]),
    .B(\V2/V1/V4/v1 [2]),
    .Z(\V2/V1/V4/A2/M1/s1 ));
 AND2_X1 \V2/V1/V4/A2/M1/M2/_0_  (.A1(\V2/V1/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M1/M2/_1_  (.A(\V2/V1/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v4 [2]));
 OR2_X1 \V2/V1/V4/A2/M1/_0_  (.A1(\V2/V1/V4/A2/M1/c1 ),
    .A2(\V2/V1/V4/A2/M1/c2 ),
    .ZN(\V2/V1/V4/A2/c1 ));
 AND2_X1 \V2/V1/V4/A2/M2/M1/_0_  (.A1(\V2/V1/V4/s1 [1]),
    .A2(\V2/V1/V4/v1 [3]),
    .ZN(\V2/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M2/M1/_1_  (.A(\V2/V1/V4/s1 [1]),
    .B(\V2/V1/V4/v1 [3]),
    .Z(\V2/V1/V4/A2/M2/s1 ));
 AND2_X1 \V2/V1/V4/A2/M2/M2/_0_  (.A1(\V2/V1/V4/A2/M2/s1 ),
    .A2(\V2/V1/V4/A2/c1 ),
    .ZN(\V2/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M2/M2/_1_  (.A(\V2/V1/V4/A2/M2/s1 ),
    .B(\V2/V1/V4/A2/c1 ),
    .Z(\V2/V1/v4 [3]));
 OR2_X1 \V2/V1/V4/A2/M2/_0_  (.A1(\V2/V1/V4/A2/M2/c1 ),
    .A2(\V2/V1/V4/A2/M2/c2 ),
    .ZN(\V2/V1/V4/A2/c2 ));
 AND2_X1 \V2/V1/V4/A2/M3/M1/_0_  (.A1(\V2/V1/V4/s1 [2]),
    .A2(ground),
    .ZN(\V2/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M3/M1/_1_  (.A(\V2/V1/V4/s1 [2]),
    .B(ground),
    .Z(\V2/V1/V4/A2/M3/s1 ));
 AND2_X1 \V2/V1/V4/A2/M3/M2/_0_  (.A1(\V2/V1/V4/A2/M3/s1 ),
    .A2(\V2/V1/V4/A2/c2 ),
    .ZN(\V2/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M3/M2/_1_  (.A(\V2/V1/V4/A2/M3/s1 ),
    .B(\V2/V1/V4/A2/c2 ),
    .Z(\V2/V1/V4/s2 [2]));
 OR2_X1 \V2/V1/V4/A2/M3/_0_  (.A1(\V2/V1/V4/A2/M3/c1 ),
    .A2(\V2/V1/V4/A2/M3/c2 ),
    .ZN(\V2/V1/V4/A2/c3 ));
 AND2_X1 \V2/V1/V4/A2/M4/M1/_0_  (.A1(\V2/V1/V4/s1 [3]),
    .A2(ground),
    .ZN(\V2/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M4/M1/_1_  (.A(\V2/V1/V4/s1 [3]),
    .B(ground),
    .Z(\V2/V1/V4/A2/M4/s1 ));
 AND2_X1 \V2/V1/V4/A2/M4/M2/_0_  (.A1(\V2/V1/V4/A2/M4/s1 ),
    .A2(\V2/V1/V4/A2/c3 ),
    .ZN(\V2/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M4/M2/_1_  (.A(\V2/V1/V4/A2/M4/s1 ),
    .B(\V2/V1/V4/A2/c3 ),
    .Z(\V2/V1/V4/s2 [3]));
 OR2_X1 \V2/V1/V4/A2/M4/_0_  (.A1(\V2/V1/V4/A2/M4/c1 ),
    .A2(\V2/V1/V4/A2/M4/c2 ),
    .ZN(\V2/V1/V4/c2 ));
 AND2_X1 \V2/V1/V4/A3/M1/M1/_0_  (.A1(\V2/V1/V4/v4 [0]),
    .A2(\V2/V1/V4/s2 [2]),
    .ZN(\V2/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M1/M1/_1_  (.A(\V2/V1/V4/v4 [0]),
    .B(\V2/V1/V4/s2 [2]),
    .Z(\V2/V1/V4/A3/M1/s1 ));
 AND2_X1 \V2/V1/V4/A3/M1/M2/_0_  (.A1(\V2/V1/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M1/M2/_1_  (.A(\V2/V1/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V1/v4 [4]));
 OR2_X1 \V2/V1/V4/A3/M1/_0_  (.A1(\V2/V1/V4/A3/M1/c1 ),
    .A2(\V2/V1/V4/A3/M1/c2 ),
    .ZN(\V2/V1/V4/A3/c1 ));
 AND2_X1 \V2/V1/V4/A3/M2/M1/_0_  (.A1(\V2/V1/V4/v4 [1]),
    .A2(\V2/V1/V4/s2 [3]),
    .ZN(\V2/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M2/M1/_1_  (.A(\V2/V1/V4/v4 [1]),
    .B(\V2/V1/V4/s2 [3]),
    .Z(\V2/V1/V4/A3/M2/s1 ));
 AND2_X1 \V2/V1/V4/A3/M2/M2/_0_  (.A1(\V2/V1/V4/A3/M2/s1 ),
    .A2(\V2/V1/V4/A3/c1 ),
    .ZN(\V2/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M2/M2/_1_  (.A(\V2/V1/V4/A3/M2/s1 ),
    .B(\V2/V1/V4/A3/c1 ),
    .Z(\V2/V1/v4 [5]));
 OR2_X1 \V2/V1/V4/A3/M2/_0_  (.A1(\V2/V1/V4/A3/M2/c1 ),
    .A2(\V2/V1/V4/A3/M2/c2 ),
    .ZN(\V2/V1/V4/A3/c2 ));
 AND2_X1 \V2/V1/V4/A3/M3/M1/_0_  (.A1(\V2/V1/V4/v4 [2]),
    .A2(\V2/V1/V4/c3 ),
    .ZN(\V2/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M3/M1/_1_  (.A(\V2/V1/V4/v4 [2]),
    .B(\V2/V1/V4/c3 ),
    .Z(\V2/V1/V4/A3/M3/s1 ));
 AND2_X1 \V2/V1/V4/A3/M3/M2/_0_  (.A1(\V2/V1/V4/A3/M3/s1 ),
    .A2(\V2/V1/V4/A3/c2 ),
    .ZN(\V2/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M3/M2/_1_  (.A(\V2/V1/V4/A3/M3/s1 ),
    .B(\V2/V1/V4/A3/c2 ),
    .Z(\V2/V1/v4 [6]));
 OR2_X1 \V2/V1/V4/A3/M3/_0_  (.A1(\V2/V1/V4/A3/M3/c1 ),
    .A2(\V2/V1/V4/A3/M3/c2 ),
    .ZN(\V2/V1/V4/A3/c3 ));
 AND2_X1 \V2/V1/V4/A3/M4/M1/_0_  (.A1(\V2/V1/V4/v4 [3]),
    .A2(ground),
    .ZN(\V2/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M4/M1/_1_  (.A(\V2/V1/V4/v4 [3]),
    .B(ground),
    .Z(\V2/V1/V4/A3/M4/s1 ));
 AND2_X1 \V2/V1/V4/A3/M4/M2/_0_  (.A1(\V2/V1/V4/A3/M4/s1 ),
    .A2(\V2/V1/V4/A3/c3 ),
    .ZN(\V2/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M4/M2/_1_  (.A(\V2/V1/V4/A3/M4/s1 ),
    .B(\V2/V1/V4/A3/c3 ),
    .Z(\V2/V1/v4 [7]));
 OR2_X1 \V2/V1/V4/A3/M4/_0_  (.A1(\V2/V1/V4/A3/M4/c1 ),
    .A2(\V2/V1/V4/A3/M4/c2 ),
    .ZN(\V2/V1/V4/overflow ));
 AND2_X1 \V2/V1/V4/V1/HA1/_0_  (.A1(\V2/V1/V4/V1/w2 ),
    .A2(\V2/V1/V4/V1/w1 ),
    .ZN(\V2/V1/V4/V1/w4 ));
 XOR2_X2 \V2/V1/V4/V1/HA1/_1_  (.A(\V2/V1/V4/V1/w2 ),
    .B(\V2/V1/V4/V1/w1 ),
    .Z(\V2/V1/v4 [1]));
 AND2_X1 \V2/V1/V4/V1/HA2/_0_  (.A1(\V2/V1/V4/V1/w4 ),
    .A2(\V2/V1/V4/V1/w3 ),
    .ZN(\V2/V1/V4/v1 [3]));
 XOR2_X2 \V2/V1/V4/V1/HA2/_1_  (.A(\V2/V1/V4/V1/w4 ),
    .B(\V2/V1/V4/V1/w3 ),
    .Z(\V2/V1/V4/v1 [2]));
 AND2_X1 \V2/V1/V4/V1/_0_  (.A1(A[20]),
    .A2(B[4]),
    .ZN(\V2/V1/v4 [0]));
 AND2_X1 \V2/V1/V4/V1/_1_  (.A1(A[20]),
    .A2(B[5]),
    .ZN(\V2/V1/V4/V1/w1 ));
 AND2_X1 \V2/V1/V4/V1/_2_  (.A1(B[4]),
    .A2(A[21]),
    .ZN(\V2/V1/V4/V1/w2 ));
 AND2_X1 \V2/V1/V4/V1/_3_  (.A1(B[5]),
    .A2(A[21]),
    .ZN(\V2/V1/V4/V1/w3 ));
 AND2_X1 \V2/V1/V4/V2/HA1/_0_  (.A1(\V2/V1/V4/V2/w2 ),
    .A2(\V2/V1/V4/V2/w1 ),
    .ZN(\V2/V1/V4/V2/w4 ));
 XOR2_X2 \V2/V1/V4/V2/HA1/_1_  (.A(\V2/V1/V4/V2/w2 ),
    .B(\V2/V1/V4/V2/w1 ),
    .Z(\V2/V1/V4/v2 [1]));
 AND2_X1 \V2/V1/V4/V2/HA2/_0_  (.A1(\V2/V1/V4/V2/w4 ),
    .A2(\V2/V1/V4/V2/w3 ),
    .ZN(\V2/V1/V4/v2 [3]));
 XOR2_X2 \V2/V1/V4/V2/HA2/_1_  (.A(\V2/V1/V4/V2/w4 ),
    .B(\V2/V1/V4/V2/w3 ),
    .Z(\V2/V1/V4/v2 [2]));
 AND2_X1 \V2/V1/V4/V2/_0_  (.A1(A[22]),
    .A2(B[4]),
    .ZN(\V2/V1/V4/v2 [0]));
 AND2_X1 \V2/V1/V4/V2/_1_  (.A1(A[22]),
    .A2(B[5]),
    .ZN(\V2/V1/V4/V2/w1 ));
 AND2_X1 \V2/V1/V4/V2/_2_  (.A1(B[4]),
    .A2(A[23]),
    .ZN(\V2/V1/V4/V2/w2 ));
 AND2_X1 \V2/V1/V4/V2/_3_  (.A1(B[5]),
    .A2(A[23]),
    .ZN(\V2/V1/V4/V2/w3 ));
 AND2_X1 \V2/V1/V4/V3/HA1/_0_  (.A1(\V2/V1/V4/V3/w2 ),
    .A2(\V2/V1/V4/V3/w1 ),
    .ZN(\V2/V1/V4/V3/w4 ));
 XOR2_X2 \V2/V1/V4/V3/HA1/_1_  (.A(\V2/V1/V4/V3/w2 ),
    .B(\V2/V1/V4/V3/w1 ),
    .Z(\V2/V1/V4/v3 [1]));
 AND2_X1 \V2/V1/V4/V3/HA2/_0_  (.A1(\V2/V1/V4/V3/w4 ),
    .A2(\V2/V1/V4/V3/w3 ),
    .ZN(\V2/V1/V4/v3 [3]));
 XOR2_X2 \V2/V1/V4/V3/HA2/_1_  (.A(\V2/V1/V4/V3/w4 ),
    .B(\V2/V1/V4/V3/w3 ),
    .Z(\V2/V1/V4/v3 [2]));
 AND2_X1 \V2/V1/V4/V3/_0_  (.A1(A[20]),
    .A2(B[6]),
    .ZN(\V2/V1/V4/v3 [0]));
 AND2_X1 \V2/V1/V4/V3/_1_  (.A1(A[20]),
    .A2(B[7]),
    .ZN(\V2/V1/V4/V3/w1 ));
 AND2_X1 \V2/V1/V4/V3/_2_  (.A1(B[6]),
    .A2(A[21]),
    .ZN(\V2/V1/V4/V3/w2 ));
 AND2_X1 \V2/V1/V4/V3/_3_  (.A1(B[7]),
    .A2(A[21]),
    .ZN(\V2/V1/V4/V3/w3 ));
 AND2_X1 \V2/V1/V4/V4/HA1/_0_  (.A1(\V2/V1/V4/V4/w2 ),
    .A2(\V2/V1/V4/V4/w1 ),
    .ZN(\V2/V1/V4/V4/w4 ));
 XOR2_X2 \V2/V1/V4/V4/HA1/_1_  (.A(\V2/V1/V4/V4/w2 ),
    .B(\V2/V1/V4/V4/w1 ),
    .Z(\V2/V1/V4/v4 [1]));
 AND2_X1 \V2/V1/V4/V4/HA2/_0_  (.A1(\V2/V1/V4/V4/w4 ),
    .A2(\V2/V1/V4/V4/w3 ),
    .ZN(\V2/V1/V4/v4 [3]));
 XOR2_X2 \V2/V1/V4/V4/HA2/_1_  (.A(\V2/V1/V4/V4/w4 ),
    .B(\V2/V1/V4/V4/w3 ),
    .Z(\V2/V1/V4/v4 [2]));
 AND2_X1 \V2/V1/V4/V4/_0_  (.A1(A[22]),
    .A2(B[6]),
    .ZN(\V2/V1/V4/v4 [0]));
 AND2_X1 \V2/V1/V4/V4/_1_  (.A1(A[22]),
    .A2(B[7]),
    .ZN(\V2/V1/V4/V4/w1 ));
 AND2_X1 \V2/V1/V4/V4/_2_  (.A1(B[6]),
    .A2(A[23]),
    .ZN(\V2/V1/V4/V4/w2 ));
 AND2_X1 \V2/V1/V4/V4/_3_  (.A1(B[7]),
    .A2(A[23]),
    .ZN(\V2/V1/V4/V4/w3 ));
 OR2_X1 \V2/V1/V4/_0_  (.A1(\V2/V1/V4/c1 ),
    .A2(\V2/V1/V4/c2 ),
    .ZN(\V2/V1/V4/c3 ));
 OR2_X1 \V2/V1/_0_  (.A1(\V2/V1/c1 ),
    .A2(\V2/V1/c2 ),
    .ZN(\V2/V1/c3 ));
 AND2_X1 \V2/V2/A1/A1/M1/M1/_0_  (.A1(\V2/V2/v2 [0]),
    .A2(\V2/V2/v3 [0]),
    .ZN(\V2/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M1/M1/_1_  (.A(\V2/V2/v2 [0]),
    .B(\V2/V2/v3 [0]),
    .Z(\V2/V2/A1/A1/M1/s1 ));
 AND2_X1 \V2/V2/A1/A1/M1/M2/_0_  (.A1(\V2/V2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M1/M2/_1_  (.A(\V2/V2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/s1 [0]));
 OR2_X1 \V2/V2/A1/A1/M1/_0_  (.A1(\V2/V2/A1/A1/M1/c1 ),
    .A2(\V2/V2/A1/A1/M1/c2 ),
    .ZN(\V2/V2/A1/A1/c1 ));
 AND2_X1 \V2/V2/A1/A1/M2/M1/_0_  (.A1(\V2/V2/v2 [1]),
    .A2(\V2/V2/v3 [1]),
    .ZN(\V2/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M2/M1/_1_  (.A(\V2/V2/v2 [1]),
    .B(\V2/V2/v3 [1]),
    .Z(\V2/V2/A1/A1/M2/s1 ));
 AND2_X1 \V2/V2/A1/A1/M2/M2/_0_  (.A1(\V2/V2/A1/A1/M2/s1 ),
    .A2(\V2/V2/A1/A1/c1 ),
    .ZN(\V2/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M2/M2/_1_  (.A(\V2/V2/A1/A1/M2/s1 ),
    .B(\V2/V2/A1/A1/c1 ),
    .Z(\V2/V2/s1 [1]));
 OR2_X1 \V2/V2/A1/A1/M2/_0_  (.A1(\V2/V2/A1/A1/M2/c1 ),
    .A2(\V2/V2/A1/A1/M2/c2 ),
    .ZN(\V2/V2/A1/A1/c2 ));
 AND2_X1 \V2/V2/A1/A1/M3/M1/_0_  (.A1(\V2/V2/v2 [2]),
    .A2(\V2/V2/v3 [2]),
    .ZN(\V2/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M3/M1/_1_  (.A(\V2/V2/v2 [2]),
    .B(\V2/V2/v3 [2]),
    .Z(\V2/V2/A1/A1/M3/s1 ));
 AND2_X1 \V2/V2/A1/A1/M3/M2/_0_  (.A1(\V2/V2/A1/A1/M3/s1 ),
    .A2(\V2/V2/A1/A1/c2 ),
    .ZN(\V2/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M3/M2/_1_  (.A(\V2/V2/A1/A1/M3/s1 ),
    .B(\V2/V2/A1/A1/c2 ),
    .Z(\V2/V2/s1 [2]));
 OR2_X1 \V2/V2/A1/A1/M3/_0_  (.A1(\V2/V2/A1/A1/M3/c1 ),
    .A2(\V2/V2/A1/A1/M3/c2 ),
    .ZN(\V2/V2/A1/A1/c3 ));
 AND2_X1 \V2/V2/A1/A1/M4/M1/_0_  (.A1(\V2/V2/v2 [3]),
    .A2(\V2/V2/v3 [3]),
    .ZN(\V2/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M4/M1/_1_  (.A(\V2/V2/v2 [3]),
    .B(\V2/V2/v3 [3]),
    .Z(\V2/V2/A1/A1/M4/s1 ));
 AND2_X1 \V2/V2/A1/A1/M4/M2/_0_  (.A1(\V2/V2/A1/A1/M4/s1 ),
    .A2(\V2/V2/A1/A1/c3 ),
    .ZN(\V2/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M4/M2/_1_  (.A(\V2/V2/A1/A1/M4/s1 ),
    .B(\V2/V2/A1/A1/c3 ),
    .Z(\V2/V2/s1 [3]));
 OR2_X1 \V2/V2/A1/A1/M4/_0_  (.A1(\V2/V2/A1/A1/M4/c1 ),
    .A2(\V2/V2/A1/A1/M4/c2 ),
    .ZN(\V2/V2/A1/c1 ));
 AND2_X1 \V2/V2/A1/A2/M1/M1/_0_  (.A1(\V2/V2/v2 [4]),
    .A2(\V2/V2/v3 [4]),
    .ZN(\V2/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M1/M1/_1_  (.A(\V2/V2/v2 [4]),
    .B(\V2/V2/v3 [4]),
    .Z(\V2/V2/A1/A2/M1/s1 ));
 AND2_X1 \V2/V2/A1/A2/M1/M2/_0_  (.A1(\V2/V2/A1/A2/M1/s1 ),
    .A2(\V2/V2/A1/c1 ),
    .ZN(\V2/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M1/M2/_1_  (.A(\V2/V2/A1/A2/M1/s1 ),
    .B(\V2/V2/A1/c1 ),
    .Z(\V2/V2/s1 [4]));
 OR2_X1 \V2/V2/A1/A2/M1/_0_  (.A1(\V2/V2/A1/A2/M1/c1 ),
    .A2(\V2/V2/A1/A2/M1/c2 ),
    .ZN(\V2/V2/A1/A2/c1 ));
 AND2_X1 \V2/V2/A1/A2/M2/M1/_0_  (.A1(\V2/V2/v2 [5]),
    .A2(\V2/V2/v3 [5]),
    .ZN(\V2/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M2/M1/_1_  (.A(\V2/V2/v2 [5]),
    .B(\V2/V2/v3 [5]),
    .Z(\V2/V2/A1/A2/M2/s1 ));
 AND2_X1 \V2/V2/A1/A2/M2/M2/_0_  (.A1(\V2/V2/A1/A2/M2/s1 ),
    .A2(\V2/V2/A1/A2/c1 ),
    .ZN(\V2/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M2/M2/_1_  (.A(\V2/V2/A1/A2/M2/s1 ),
    .B(\V2/V2/A1/A2/c1 ),
    .Z(\V2/V2/s1 [5]));
 OR2_X1 \V2/V2/A1/A2/M2/_0_  (.A1(\V2/V2/A1/A2/M2/c1 ),
    .A2(\V2/V2/A1/A2/M2/c2 ),
    .ZN(\V2/V2/A1/A2/c2 ));
 AND2_X1 \V2/V2/A1/A2/M3/M1/_0_  (.A1(\V2/V2/v2 [6]),
    .A2(\V2/V2/v3 [6]),
    .ZN(\V2/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M3/M1/_1_  (.A(\V2/V2/v2 [6]),
    .B(\V2/V2/v3 [6]),
    .Z(\V2/V2/A1/A2/M3/s1 ));
 AND2_X1 \V2/V2/A1/A2/M3/M2/_0_  (.A1(\V2/V2/A1/A2/M3/s1 ),
    .A2(\V2/V2/A1/A2/c2 ),
    .ZN(\V2/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M3/M2/_1_  (.A(\V2/V2/A1/A2/M3/s1 ),
    .B(\V2/V2/A1/A2/c2 ),
    .Z(\V2/V2/s1 [6]));
 OR2_X1 \V2/V2/A1/A2/M3/_0_  (.A1(\V2/V2/A1/A2/M3/c1 ),
    .A2(\V2/V2/A1/A2/M3/c2 ),
    .ZN(\V2/V2/A1/A2/c3 ));
 AND2_X1 \V2/V2/A1/A2/M4/M1/_0_  (.A1(\V2/V2/v2 [7]),
    .A2(\V2/V2/v3 [7]),
    .ZN(\V2/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M4/M1/_1_  (.A(\V2/V2/v2 [7]),
    .B(\V2/V2/v3 [7]),
    .Z(\V2/V2/A1/A2/M4/s1 ));
 AND2_X1 \V2/V2/A1/A2/M4/M2/_0_  (.A1(\V2/V2/A1/A2/M4/s1 ),
    .A2(\V2/V2/A1/A2/c3 ),
    .ZN(\V2/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M4/M2/_1_  (.A(\V2/V2/A1/A2/M4/s1 ),
    .B(\V2/V2/A1/A2/c3 ),
    .Z(\V2/V2/s1 [7]));
 OR2_X1 \V2/V2/A1/A2/M4/_0_  (.A1(\V2/V2/A1/A2/M4/c1 ),
    .A2(\V2/V2/A1/A2/M4/c2 ),
    .ZN(\V2/V2/c1 ));
 AND2_X1 \V2/V2/A2/A1/M1/M1/_0_  (.A1(\V2/V2/s1 [0]),
    .A2(\V2/V2/v1 [4]),
    .ZN(\V2/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M1/M1/_1_  (.A(\V2/V2/s1 [0]),
    .B(\V2/V2/v1 [4]),
    .Z(\V2/V2/A2/A1/M1/s1 ));
 AND2_X1 \V2/V2/A2/A1/M1/M2/_0_  (.A1(\V2/V2/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M1/M2/_1_  (.A(\V2/V2/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v2 [4]));
 OR2_X1 \V2/V2/A2/A1/M1/_0_  (.A1(\V2/V2/A2/A1/M1/c1 ),
    .A2(\V2/V2/A2/A1/M1/c2 ),
    .ZN(\V2/V2/A2/A1/c1 ));
 AND2_X1 \V2/V2/A2/A1/M2/M1/_0_  (.A1(\V2/V2/s1 [1]),
    .A2(\V2/V2/v1 [5]),
    .ZN(\V2/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M2/M1/_1_  (.A(\V2/V2/s1 [1]),
    .B(\V2/V2/v1 [5]),
    .Z(\V2/V2/A2/A1/M2/s1 ));
 AND2_X1 \V2/V2/A2/A1/M2/M2/_0_  (.A1(\V2/V2/A2/A1/M2/s1 ),
    .A2(\V2/V2/A2/A1/c1 ),
    .ZN(\V2/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M2/M2/_1_  (.A(\V2/V2/A2/A1/M2/s1 ),
    .B(\V2/V2/A2/A1/c1 ),
    .Z(\V2/v2 [5]));
 OR2_X1 \V2/V2/A2/A1/M2/_0_  (.A1(\V2/V2/A2/A1/M2/c1 ),
    .A2(\V2/V2/A2/A1/M2/c2 ),
    .ZN(\V2/V2/A2/A1/c2 ));
 AND2_X1 \V2/V2/A2/A1/M3/M1/_0_  (.A1(\V2/V2/s1 [2]),
    .A2(\V2/V2/v1 [6]),
    .ZN(\V2/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M3/M1/_1_  (.A(\V2/V2/s1 [2]),
    .B(\V2/V2/v1 [6]),
    .Z(\V2/V2/A2/A1/M3/s1 ));
 AND2_X1 \V2/V2/A2/A1/M3/M2/_0_  (.A1(\V2/V2/A2/A1/M3/s1 ),
    .A2(\V2/V2/A2/A1/c2 ),
    .ZN(\V2/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M3/M2/_1_  (.A(\V2/V2/A2/A1/M3/s1 ),
    .B(\V2/V2/A2/A1/c2 ),
    .Z(\V2/v2 [6]));
 OR2_X1 \V2/V2/A2/A1/M3/_0_  (.A1(\V2/V2/A2/A1/M3/c1 ),
    .A2(\V2/V2/A2/A1/M3/c2 ),
    .ZN(\V2/V2/A2/A1/c3 ));
 AND2_X1 \V2/V2/A2/A1/M4/M1/_0_  (.A1(\V2/V2/s1 [3]),
    .A2(\V2/V2/v1 [7]),
    .ZN(\V2/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M4/M1/_1_  (.A(\V2/V2/s1 [3]),
    .B(\V2/V2/v1 [7]),
    .Z(\V2/V2/A2/A1/M4/s1 ));
 AND2_X1 \V2/V2/A2/A1/M4/M2/_0_  (.A1(\V2/V2/A2/A1/M4/s1 ),
    .A2(\V2/V2/A2/A1/c3 ),
    .ZN(\V2/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M4/M2/_1_  (.A(\V2/V2/A2/A1/M4/s1 ),
    .B(\V2/V2/A2/A1/c3 ),
    .Z(\V2/v2 [7]));
 OR2_X1 \V2/V2/A2/A1/M4/_0_  (.A1(\V2/V2/A2/A1/M4/c1 ),
    .A2(\V2/V2/A2/A1/M4/c2 ),
    .ZN(\V2/V2/A2/c1 ));
 AND2_X1 \V2/V2/A2/A2/M1/M1/_0_  (.A1(\V2/V2/s1 [4]),
    .A2(ground),
    .ZN(\V2/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M1/M1/_1_  (.A(\V2/V2/s1 [4]),
    .B(ground),
    .Z(\V2/V2/A2/A2/M1/s1 ));
 AND2_X1 \V2/V2/A2/A2/M1/M2/_0_  (.A1(\V2/V2/A2/A2/M1/s1 ),
    .A2(\V2/V2/A2/c1 ),
    .ZN(\V2/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M1/M2/_1_  (.A(\V2/V2/A2/A2/M1/s1 ),
    .B(\V2/V2/A2/c1 ),
    .Z(\V2/V2/s2 [4]));
 OR2_X1 \V2/V2/A2/A2/M1/_0_  (.A1(\V2/V2/A2/A2/M1/c1 ),
    .A2(\V2/V2/A2/A2/M1/c2 ),
    .ZN(\V2/V2/A2/A2/c1 ));
 AND2_X1 \V2/V2/A2/A2/M2/M1/_0_  (.A1(\V2/V2/s1 [5]),
    .A2(ground),
    .ZN(\V2/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M2/M1/_1_  (.A(\V2/V2/s1 [5]),
    .B(ground),
    .Z(\V2/V2/A2/A2/M2/s1 ));
 AND2_X1 \V2/V2/A2/A2/M2/M2/_0_  (.A1(\V2/V2/A2/A2/M2/s1 ),
    .A2(\V2/V2/A2/A2/c1 ),
    .ZN(\V2/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M2/M2/_1_  (.A(\V2/V2/A2/A2/M2/s1 ),
    .B(\V2/V2/A2/A2/c1 ),
    .Z(\V2/V2/s2 [5]));
 OR2_X1 \V2/V2/A2/A2/M2/_0_  (.A1(\V2/V2/A2/A2/M2/c1 ),
    .A2(\V2/V2/A2/A2/M2/c2 ),
    .ZN(\V2/V2/A2/A2/c2 ));
 AND2_X1 \V2/V2/A2/A2/M3/M1/_0_  (.A1(\V2/V2/s1 [6]),
    .A2(ground),
    .ZN(\V2/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M3/M1/_1_  (.A(\V2/V2/s1 [6]),
    .B(ground),
    .Z(\V2/V2/A2/A2/M3/s1 ));
 AND2_X1 \V2/V2/A2/A2/M3/M2/_0_  (.A1(\V2/V2/A2/A2/M3/s1 ),
    .A2(\V2/V2/A2/A2/c2 ),
    .ZN(\V2/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M3/M2/_1_  (.A(\V2/V2/A2/A2/M3/s1 ),
    .B(\V2/V2/A2/A2/c2 ),
    .Z(\V2/V2/s2 [6]));
 OR2_X1 \V2/V2/A2/A2/M3/_0_  (.A1(\V2/V2/A2/A2/M3/c1 ),
    .A2(\V2/V2/A2/A2/M3/c2 ),
    .ZN(\V2/V2/A2/A2/c3 ));
 AND2_X1 \V2/V2/A2/A2/M4/M1/_0_  (.A1(\V2/V2/s1 [7]),
    .A2(ground),
    .ZN(\V2/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M4/M1/_1_  (.A(\V2/V2/s1 [7]),
    .B(ground),
    .Z(\V2/V2/A2/A2/M4/s1 ));
 AND2_X1 \V2/V2/A2/A2/M4/M2/_0_  (.A1(\V2/V2/A2/A2/M4/s1 ),
    .A2(\V2/V2/A2/A2/c3 ),
    .ZN(\V2/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M4/M2/_1_  (.A(\V2/V2/A2/A2/M4/s1 ),
    .B(\V2/V2/A2/A2/c3 ),
    .Z(\V2/V2/s2 [7]));
 OR2_X1 \V2/V2/A2/A2/M4/_0_  (.A1(\V2/V2/A2/A2/M4/c1 ),
    .A2(\V2/V2/A2/A2/M4/c2 ),
    .ZN(\V2/V2/c2 ));
 AND2_X1 \V2/V2/A3/A1/M1/M1/_0_  (.A1(\V2/V2/v4 [0]),
    .A2(\V2/V2/s2 [4]),
    .ZN(\V2/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M1/M1/_1_  (.A(\V2/V2/v4 [0]),
    .B(\V2/V2/s2 [4]),
    .Z(\V2/V2/A3/A1/M1/s1 ));
 AND2_X1 \V2/V2/A3/A1/M1/M2/_0_  (.A1(\V2/V2/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M1/M2/_1_  (.A(\V2/V2/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v2 [8]));
 OR2_X1 \V2/V2/A3/A1/M1/_0_  (.A1(\V2/V2/A3/A1/M1/c1 ),
    .A2(\V2/V2/A3/A1/M1/c2 ),
    .ZN(\V2/V2/A3/A1/c1 ));
 AND2_X1 \V2/V2/A3/A1/M2/M1/_0_  (.A1(\V2/V2/v4 [1]),
    .A2(\V2/V2/s2 [5]),
    .ZN(\V2/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M2/M1/_1_  (.A(\V2/V2/v4 [1]),
    .B(\V2/V2/s2 [5]),
    .Z(\V2/V2/A3/A1/M2/s1 ));
 AND2_X1 \V2/V2/A3/A1/M2/M2/_0_  (.A1(\V2/V2/A3/A1/M2/s1 ),
    .A2(\V2/V2/A3/A1/c1 ),
    .ZN(\V2/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M2/M2/_1_  (.A(\V2/V2/A3/A1/M2/s1 ),
    .B(\V2/V2/A3/A1/c1 ),
    .Z(\V2/v2 [9]));
 OR2_X1 \V2/V2/A3/A1/M2/_0_  (.A1(\V2/V2/A3/A1/M2/c1 ),
    .A2(\V2/V2/A3/A1/M2/c2 ),
    .ZN(\V2/V2/A3/A1/c2 ));
 AND2_X1 \V2/V2/A3/A1/M3/M1/_0_  (.A1(\V2/V2/v4 [2]),
    .A2(\V2/V2/s2 [6]),
    .ZN(\V2/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M3/M1/_1_  (.A(\V2/V2/v4 [2]),
    .B(\V2/V2/s2 [6]),
    .Z(\V2/V2/A3/A1/M3/s1 ));
 AND2_X1 \V2/V2/A3/A1/M3/M2/_0_  (.A1(\V2/V2/A3/A1/M3/s1 ),
    .A2(\V2/V2/A3/A1/c2 ),
    .ZN(\V2/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M3/M2/_1_  (.A(\V2/V2/A3/A1/M3/s1 ),
    .B(\V2/V2/A3/A1/c2 ),
    .Z(\V2/v2 [10]));
 OR2_X1 \V2/V2/A3/A1/M3/_0_  (.A1(\V2/V2/A3/A1/M3/c1 ),
    .A2(\V2/V2/A3/A1/M3/c2 ),
    .ZN(\V2/V2/A3/A1/c3 ));
 AND2_X1 \V2/V2/A3/A1/M4/M1/_0_  (.A1(\V2/V2/v4 [3]),
    .A2(\V2/V2/s2 [7]),
    .ZN(\V2/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M4/M1/_1_  (.A(\V2/V2/v4 [3]),
    .B(\V2/V2/s2 [7]),
    .Z(\V2/V2/A3/A1/M4/s1 ));
 AND2_X1 \V2/V2/A3/A1/M4/M2/_0_  (.A1(\V2/V2/A3/A1/M4/s1 ),
    .A2(\V2/V2/A3/A1/c3 ),
    .ZN(\V2/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M4/M2/_1_  (.A(\V2/V2/A3/A1/M4/s1 ),
    .B(\V2/V2/A3/A1/c3 ),
    .Z(\V2/v2 [11]));
 OR2_X1 \V2/V2/A3/A1/M4/_0_  (.A1(\V2/V2/A3/A1/M4/c1 ),
    .A2(\V2/V2/A3/A1/M4/c2 ),
    .ZN(\V2/V2/A3/c1 ));
 AND2_X1 \V2/V2/A3/A2/M1/M1/_0_  (.A1(\V2/V2/v4 [4]),
    .A2(\V2/V2/c3 ),
    .ZN(\V2/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M1/M1/_1_  (.A(\V2/V2/v4 [4]),
    .B(\V2/V2/c3 ),
    .Z(\V2/V2/A3/A2/M1/s1 ));
 AND2_X1 \V2/V2/A3/A2/M1/M2/_0_  (.A1(\V2/V2/A3/A2/M1/s1 ),
    .A2(\V2/V2/A3/c1 ),
    .ZN(\V2/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M1/M2/_1_  (.A(\V2/V2/A3/A2/M1/s1 ),
    .B(\V2/V2/A3/c1 ),
    .Z(\V2/v2 [12]));
 OR2_X1 \V2/V2/A3/A2/M1/_0_  (.A1(\V2/V2/A3/A2/M1/c1 ),
    .A2(\V2/V2/A3/A2/M1/c2 ),
    .ZN(\V2/V2/A3/A2/c1 ));
 AND2_X1 \V2/V2/A3/A2/M2/M1/_0_  (.A1(\V2/V2/v4 [5]),
    .A2(ground),
    .ZN(\V2/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M2/M1/_1_  (.A(\V2/V2/v4 [5]),
    .B(ground),
    .Z(\V2/V2/A3/A2/M2/s1 ));
 AND2_X1 \V2/V2/A3/A2/M2/M2/_0_  (.A1(\V2/V2/A3/A2/M2/s1 ),
    .A2(\V2/V2/A3/A2/c1 ),
    .ZN(\V2/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M2/M2/_1_  (.A(\V2/V2/A3/A2/M2/s1 ),
    .B(\V2/V2/A3/A2/c1 ),
    .Z(\V2/v2 [13]));
 OR2_X1 \V2/V2/A3/A2/M2/_0_  (.A1(\V2/V2/A3/A2/M2/c1 ),
    .A2(\V2/V2/A3/A2/M2/c2 ),
    .ZN(\V2/V2/A3/A2/c2 ));
 AND2_X1 \V2/V2/A3/A2/M3/M1/_0_  (.A1(\V2/V2/v4 [6]),
    .A2(ground),
    .ZN(\V2/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M3/M1/_1_  (.A(\V2/V2/v4 [6]),
    .B(ground),
    .Z(\V2/V2/A3/A2/M3/s1 ));
 AND2_X1 \V2/V2/A3/A2/M3/M2/_0_  (.A1(\V2/V2/A3/A2/M3/s1 ),
    .A2(\V2/V2/A3/A2/c2 ),
    .ZN(\V2/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M3/M2/_1_  (.A(\V2/V2/A3/A2/M3/s1 ),
    .B(\V2/V2/A3/A2/c2 ),
    .Z(\V2/v2 [14]));
 OR2_X1 \V2/V2/A3/A2/M3/_0_  (.A1(\V2/V2/A3/A2/M3/c1 ),
    .A2(\V2/V2/A3/A2/M3/c2 ),
    .ZN(\V2/V2/A3/A2/c3 ));
 AND2_X1 \V2/V2/A3/A2/M4/M1/_0_  (.A1(\V2/V2/v4 [7]),
    .A2(ground),
    .ZN(\V2/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M4/M1/_1_  (.A(\V2/V2/v4 [7]),
    .B(ground),
    .Z(\V2/V2/A3/A2/M4/s1 ));
 AND2_X1 \V2/V2/A3/A2/M4/M2/_0_  (.A1(\V2/V2/A3/A2/M4/s1 ),
    .A2(\V2/V2/A3/A2/c3 ),
    .ZN(\V2/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M4/M2/_1_  (.A(\V2/V2/A3/A2/M4/s1 ),
    .B(\V2/V2/A3/A2/c3 ),
    .Z(\V2/v2 [15]));
 OR2_X1 \V2/V2/A3/A2/M4/_0_  (.A1(\V2/V2/A3/A2/M4/c1 ),
    .A2(\V2/V2/A3/A2/M4/c2 ),
    .ZN(\V2/V2/overflow ));
 AND2_X1 \V2/V2/V1/A1/M1/M1/_0_  (.A1(\V2/V2/V1/v2 [0]),
    .A2(\V2/V2/V1/v3 [0]),
    .ZN(\V2/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M1/M1/_1_  (.A(\V2/V2/V1/v2 [0]),
    .B(\V2/V2/V1/v3 [0]),
    .Z(\V2/V2/V1/A1/M1/s1 ));
 AND2_X1 \V2/V2/V1/A1/M1/M2/_0_  (.A1(\V2/V2/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M1/M2/_1_  (.A(\V2/V2/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/V1/s1 [0]));
 OR2_X1 \V2/V2/V1/A1/M1/_0_  (.A1(\V2/V2/V1/A1/M1/c1 ),
    .A2(\V2/V2/V1/A1/M1/c2 ),
    .ZN(\V2/V2/V1/A1/c1 ));
 AND2_X1 \V2/V2/V1/A1/M2/M1/_0_  (.A1(\V2/V2/V1/v2 [1]),
    .A2(\V2/V2/V1/v3 [1]),
    .ZN(\V2/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M2/M1/_1_  (.A(\V2/V2/V1/v2 [1]),
    .B(\V2/V2/V1/v3 [1]),
    .Z(\V2/V2/V1/A1/M2/s1 ));
 AND2_X1 \V2/V2/V1/A1/M2/M2/_0_  (.A1(\V2/V2/V1/A1/M2/s1 ),
    .A2(\V2/V2/V1/A1/c1 ),
    .ZN(\V2/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M2/M2/_1_  (.A(\V2/V2/V1/A1/M2/s1 ),
    .B(\V2/V2/V1/A1/c1 ),
    .Z(\V2/V2/V1/s1 [1]));
 OR2_X1 \V2/V2/V1/A1/M2/_0_  (.A1(\V2/V2/V1/A1/M2/c1 ),
    .A2(\V2/V2/V1/A1/M2/c2 ),
    .ZN(\V2/V2/V1/A1/c2 ));
 AND2_X1 \V2/V2/V1/A1/M3/M1/_0_  (.A1(\V2/V2/V1/v2 [2]),
    .A2(\V2/V2/V1/v3 [2]),
    .ZN(\V2/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M3/M1/_1_  (.A(\V2/V2/V1/v2 [2]),
    .B(\V2/V2/V1/v3 [2]),
    .Z(\V2/V2/V1/A1/M3/s1 ));
 AND2_X1 \V2/V2/V1/A1/M3/M2/_0_  (.A1(\V2/V2/V1/A1/M3/s1 ),
    .A2(\V2/V2/V1/A1/c2 ),
    .ZN(\V2/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M3/M2/_1_  (.A(\V2/V2/V1/A1/M3/s1 ),
    .B(\V2/V2/V1/A1/c2 ),
    .Z(\V2/V2/V1/s1 [2]));
 OR2_X1 \V2/V2/V1/A1/M3/_0_  (.A1(\V2/V2/V1/A1/M3/c1 ),
    .A2(\V2/V2/V1/A1/M3/c2 ),
    .ZN(\V2/V2/V1/A1/c3 ));
 AND2_X1 \V2/V2/V1/A1/M4/M1/_0_  (.A1(\V2/V2/V1/v2 [3]),
    .A2(\V2/V2/V1/v3 [3]),
    .ZN(\V2/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M4/M1/_1_  (.A(\V2/V2/V1/v2 [3]),
    .B(\V2/V2/V1/v3 [3]),
    .Z(\V2/V2/V1/A1/M4/s1 ));
 AND2_X1 \V2/V2/V1/A1/M4/M2/_0_  (.A1(\V2/V2/V1/A1/M4/s1 ),
    .A2(\V2/V2/V1/A1/c3 ),
    .ZN(\V2/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M4/M2/_1_  (.A(\V2/V2/V1/A1/M4/s1 ),
    .B(\V2/V2/V1/A1/c3 ),
    .Z(\V2/V2/V1/s1 [3]));
 OR2_X1 \V2/V2/V1/A1/M4/_0_  (.A1(\V2/V2/V1/A1/M4/c1 ),
    .A2(\V2/V2/V1/A1/M4/c2 ),
    .ZN(\V2/V2/V1/c1 ));
 AND2_X1 \V2/V2/V1/A2/M1/M1/_0_  (.A1(\V2/V2/V1/s1 [0]),
    .A2(\V2/V2/V1/v1 [2]),
    .ZN(\V2/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M1/M1/_1_  (.A(\V2/V2/V1/s1 [0]),
    .B(\V2/V2/V1/v1 [2]),
    .Z(\V2/V2/V1/A2/M1/s1 ));
 AND2_X1 \V2/V2/V1/A2/M1/M2/_0_  (.A1(\V2/V2/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M1/M2/_1_  (.A(\V2/V2/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/v2 [2]));
 OR2_X1 \V2/V2/V1/A2/M1/_0_  (.A1(\V2/V2/V1/A2/M1/c1 ),
    .A2(\V2/V2/V1/A2/M1/c2 ),
    .ZN(\V2/V2/V1/A2/c1 ));
 AND2_X1 \V2/V2/V1/A2/M2/M1/_0_  (.A1(\V2/V2/V1/s1 [1]),
    .A2(\V2/V2/V1/v1 [3]),
    .ZN(\V2/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M2/M1/_1_  (.A(\V2/V2/V1/s1 [1]),
    .B(\V2/V2/V1/v1 [3]),
    .Z(\V2/V2/V1/A2/M2/s1 ));
 AND2_X1 \V2/V2/V1/A2/M2/M2/_0_  (.A1(\V2/V2/V1/A2/M2/s1 ),
    .A2(\V2/V2/V1/A2/c1 ),
    .ZN(\V2/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M2/M2/_1_  (.A(\V2/V2/V1/A2/M2/s1 ),
    .B(\V2/V2/V1/A2/c1 ),
    .Z(\V2/v2 [3]));
 OR2_X1 \V2/V2/V1/A2/M2/_0_  (.A1(\V2/V2/V1/A2/M2/c1 ),
    .A2(\V2/V2/V1/A2/M2/c2 ),
    .ZN(\V2/V2/V1/A2/c2 ));
 AND2_X1 \V2/V2/V1/A2/M3/M1/_0_  (.A1(\V2/V2/V1/s1 [2]),
    .A2(ground),
    .ZN(\V2/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M3/M1/_1_  (.A(\V2/V2/V1/s1 [2]),
    .B(ground),
    .Z(\V2/V2/V1/A2/M3/s1 ));
 AND2_X1 \V2/V2/V1/A2/M3/M2/_0_  (.A1(\V2/V2/V1/A2/M3/s1 ),
    .A2(\V2/V2/V1/A2/c2 ),
    .ZN(\V2/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M3/M2/_1_  (.A(\V2/V2/V1/A2/M3/s1 ),
    .B(\V2/V2/V1/A2/c2 ),
    .Z(\V2/V2/V1/s2 [2]));
 OR2_X1 \V2/V2/V1/A2/M3/_0_  (.A1(\V2/V2/V1/A2/M3/c1 ),
    .A2(\V2/V2/V1/A2/M3/c2 ),
    .ZN(\V2/V2/V1/A2/c3 ));
 AND2_X1 \V2/V2/V1/A2/M4/M1/_0_  (.A1(\V2/V2/V1/s1 [3]),
    .A2(ground),
    .ZN(\V2/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M4/M1/_1_  (.A(\V2/V2/V1/s1 [3]),
    .B(ground),
    .Z(\V2/V2/V1/A2/M4/s1 ));
 AND2_X1 \V2/V2/V1/A2/M4/M2/_0_  (.A1(\V2/V2/V1/A2/M4/s1 ),
    .A2(\V2/V2/V1/A2/c3 ),
    .ZN(\V2/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M4/M2/_1_  (.A(\V2/V2/V1/A2/M4/s1 ),
    .B(\V2/V2/V1/A2/c3 ),
    .Z(\V2/V2/V1/s2 [3]));
 OR2_X1 \V2/V2/V1/A2/M4/_0_  (.A1(\V2/V2/V1/A2/M4/c1 ),
    .A2(\V2/V2/V1/A2/M4/c2 ),
    .ZN(\V2/V2/V1/c2 ));
 AND2_X1 \V2/V2/V1/A3/M1/M1/_0_  (.A1(\V2/V2/V1/v4 [0]),
    .A2(\V2/V2/V1/s2 [2]),
    .ZN(\V2/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M1/M1/_1_  (.A(\V2/V2/V1/v4 [0]),
    .B(\V2/V2/V1/s2 [2]),
    .Z(\V2/V2/V1/A3/M1/s1 ));
 AND2_X1 \V2/V2/V1/A3/M1/M2/_0_  (.A1(\V2/V2/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M1/M2/_1_  (.A(\V2/V2/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v1 [4]));
 OR2_X1 \V2/V2/V1/A3/M1/_0_  (.A1(\V2/V2/V1/A3/M1/c1 ),
    .A2(\V2/V2/V1/A3/M1/c2 ),
    .ZN(\V2/V2/V1/A3/c1 ));
 AND2_X1 \V2/V2/V1/A3/M2/M1/_0_  (.A1(\V2/V2/V1/v4 [1]),
    .A2(\V2/V2/V1/s2 [3]),
    .ZN(\V2/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M2/M1/_1_  (.A(\V2/V2/V1/v4 [1]),
    .B(\V2/V2/V1/s2 [3]),
    .Z(\V2/V2/V1/A3/M2/s1 ));
 AND2_X1 \V2/V2/V1/A3/M2/M2/_0_  (.A1(\V2/V2/V1/A3/M2/s1 ),
    .A2(\V2/V2/V1/A3/c1 ),
    .ZN(\V2/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M2/M2/_1_  (.A(\V2/V2/V1/A3/M2/s1 ),
    .B(\V2/V2/V1/A3/c1 ),
    .Z(\V2/V2/v1 [5]));
 OR2_X1 \V2/V2/V1/A3/M2/_0_  (.A1(\V2/V2/V1/A3/M2/c1 ),
    .A2(\V2/V2/V1/A3/M2/c2 ),
    .ZN(\V2/V2/V1/A3/c2 ));
 AND2_X1 \V2/V2/V1/A3/M3/M1/_0_  (.A1(\V2/V2/V1/v4 [2]),
    .A2(\V2/V2/V1/c3 ),
    .ZN(\V2/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M3/M1/_1_  (.A(\V2/V2/V1/v4 [2]),
    .B(\V2/V2/V1/c3 ),
    .Z(\V2/V2/V1/A3/M3/s1 ));
 AND2_X1 \V2/V2/V1/A3/M3/M2/_0_  (.A1(\V2/V2/V1/A3/M3/s1 ),
    .A2(\V2/V2/V1/A3/c2 ),
    .ZN(\V2/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M3/M2/_1_  (.A(\V2/V2/V1/A3/M3/s1 ),
    .B(\V2/V2/V1/A3/c2 ),
    .Z(\V2/V2/v1 [6]));
 OR2_X1 \V2/V2/V1/A3/M3/_0_  (.A1(\V2/V2/V1/A3/M3/c1 ),
    .A2(\V2/V2/V1/A3/M3/c2 ),
    .ZN(\V2/V2/V1/A3/c3 ));
 AND2_X1 \V2/V2/V1/A3/M4/M1/_0_  (.A1(\V2/V2/V1/v4 [3]),
    .A2(ground),
    .ZN(\V2/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M4/M1/_1_  (.A(\V2/V2/V1/v4 [3]),
    .B(ground),
    .Z(\V2/V2/V1/A3/M4/s1 ));
 AND2_X1 \V2/V2/V1/A3/M4/M2/_0_  (.A1(\V2/V2/V1/A3/M4/s1 ),
    .A2(\V2/V2/V1/A3/c3 ),
    .ZN(\V2/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M4/M2/_1_  (.A(\V2/V2/V1/A3/M4/s1 ),
    .B(\V2/V2/V1/A3/c3 ),
    .Z(\V2/V2/v1 [7]));
 OR2_X1 \V2/V2/V1/A3/M4/_0_  (.A1(\V2/V2/V1/A3/M4/c1 ),
    .A2(\V2/V2/V1/A3/M4/c2 ),
    .ZN(\V2/V2/V1/overflow ));
 AND2_X1 \V2/V2/V1/V1/HA1/_0_  (.A1(\V2/V2/V1/V1/w2 ),
    .A2(\V2/V2/V1/V1/w1 ),
    .ZN(\V2/V2/V1/V1/w4 ));
 XOR2_X2 \V2/V2/V1/V1/HA1/_1_  (.A(\V2/V2/V1/V1/w2 ),
    .B(\V2/V2/V1/V1/w1 ),
    .Z(\V2/v2 [1]));
 AND2_X1 \V2/V2/V1/V1/HA2/_0_  (.A1(\V2/V2/V1/V1/w4 ),
    .A2(\V2/V2/V1/V1/w3 ),
    .ZN(\V2/V2/V1/v1 [3]));
 XOR2_X2 \V2/V2/V1/V1/HA2/_1_  (.A(\V2/V2/V1/V1/w4 ),
    .B(\V2/V2/V1/V1/w3 ),
    .Z(\V2/V2/V1/v1 [2]));
 AND2_X1 \V2/V2/V1/V1/_0_  (.A1(A[24]),
    .A2(B[0]),
    .ZN(\V2/v2 [0]));
 AND2_X1 \V2/V2/V1/V1/_1_  (.A1(A[24]),
    .A2(B[1]),
    .ZN(\V2/V2/V1/V1/w1 ));
 AND2_X1 \V2/V2/V1/V1/_2_  (.A1(B[0]),
    .A2(A[25]),
    .ZN(\V2/V2/V1/V1/w2 ));
 AND2_X1 \V2/V2/V1/V1/_3_  (.A1(B[1]),
    .A2(A[25]),
    .ZN(\V2/V2/V1/V1/w3 ));
 AND2_X1 \V2/V2/V1/V2/HA1/_0_  (.A1(\V2/V2/V1/V2/w2 ),
    .A2(\V2/V2/V1/V2/w1 ),
    .ZN(\V2/V2/V1/V2/w4 ));
 XOR2_X2 \V2/V2/V1/V2/HA1/_1_  (.A(\V2/V2/V1/V2/w2 ),
    .B(\V2/V2/V1/V2/w1 ),
    .Z(\V2/V2/V1/v2 [1]));
 AND2_X1 \V2/V2/V1/V2/HA2/_0_  (.A1(\V2/V2/V1/V2/w4 ),
    .A2(\V2/V2/V1/V2/w3 ),
    .ZN(\V2/V2/V1/v2 [3]));
 XOR2_X2 \V2/V2/V1/V2/HA2/_1_  (.A(\V2/V2/V1/V2/w4 ),
    .B(\V2/V2/V1/V2/w3 ),
    .Z(\V2/V2/V1/v2 [2]));
 AND2_X1 \V2/V2/V1/V2/_0_  (.A1(A[26]),
    .A2(B[0]),
    .ZN(\V2/V2/V1/v2 [0]));
 AND2_X1 \V2/V2/V1/V2/_1_  (.A1(A[26]),
    .A2(B[1]),
    .ZN(\V2/V2/V1/V2/w1 ));
 AND2_X1 \V2/V2/V1/V2/_2_  (.A1(B[0]),
    .A2(A[27]),
    .ZN(\V2/V2/V1/V2/w2 ));
 AND2_X1 \V2/V2/V1/V2/_3_  (.A1(B[1]),
    .A2(A[27]),
    .ZN(\V2/V2/V1/V2/w3 ));
 AND2_X1 \V2/V2/V1/V3/HA1/_0_  (.A1(\V2/V2/V1/V3/w2 ),
    .A2(\V2/V2/V1/V3/w1 ),
    .ZN(\V2/V2/V1/V3/w4 ));
 XOR2_X2 \V2/V2/V1/V3/HA1/_1_  (.A(\V2/V2/V1/V3/w2 ),
    .B(\V2/V2/V1/V3/w1 ),
    .Z(\V2/V2/V1/v3 [1]));
 AND2_X1 \V2/V2/V1/V3/HA2/_0_  (.A1(\V2/V2/V1/V3/w4 ),
    .A2(\V2/V2/V1/V3/w3 ),
    .ZN(\V2/V2/V1/v3 [3]));
 XOR2_X2 \V2/V2/V1/V3/HA2/_1_  (.A(\V2/V2/V1/V3/w4 ),
    .B(\V2/V2/V1/V3/w3 ),
    .Z(\V2/V2/V1/v3 [2]));
 AND2_X1 \V2/V2/V1/V3/_0_  (.A1(A[24]),
    .A2(B[2]),
    .ZN(\V2/V2/V1/v3 [0]));
 AND2_X1 \V2/V2/V1/V3/_1_  (.A1(A[24]),
    .A2(B[3]),
    .ZN(\V2/V2/V1/V3/w1 ));
 AND2_X1 \V2/V2/V1/V3/_2_  (.A1(B[2]),
    .A2(A[25]),
    .ZN(\V2/V2/V1/V3/w2 ));
 AND2_X1 \V2/V2/V1/V3/_3_  (.A1(B[3]),
    .A2(A[25]),
    .ZN(\V2/V2/V1/V3/w3 ));
 AND2_X1 \V2/V2/V1/V4/HA1/_0_  (.A1(\V2/V2/V1/V4/w2 ),
    .A2(\V2/V2/V1/V4/w1 ),
    .ZN(\V2/V2/V1/V4/w4 ));
 XOR2_X2 \V2/V2/V1/V4/HA1/_1_  (.A(\V2/V2/V1/V4/w2 ),
    .B(\V2/V2/V1/V4/w1 ),
    .Z(\V2/V2/V1/v4 [1]));
 AND2_X1 \V2/V2/V1/V4/HA2/_0_  (.A1(\V2/V2/V1/V4/w4 ),
    .A2(\V2/V2/V1/V4/w3 ),
    .ZN(\V2/V2/V1/v4 [3]));
 XOR2_X2 \V2/V2/V1/V4/HA2/_1_  (.A(\V2/V2/V1/V4/w4 ),
    .B(\V2/V2/V1/V4/w3 ),
    .Z(\V2/V2/V1/v4 [2]));
 AND2_X1 \V2/V2/V1/V4/_0_  (.A1(A[26]),
    .A2(B[2]),
    .ZN(\V2/V2/V1/v4 [0]));
 AND2_X1 \V2/V2/V1/V4/_1_  (.A1(A[26]),
    .A2(B[3]),
    .ZN(\V2/V2/V1/V4/w1 ));
 AND2_X1 \V2/V2/V1/V4/_2_  (.A1(B[2]),
    .A2(A[27]),
    .ZN(\V2/V2/V1/V4/w2 ));
 AND2_X1 \V2/V2/V1/V4/_3_  (.A1(B[3]),
    .A2(A[27]),
    .ZN(\V2/V2/V1/V4/w3 ));
 OR2_X1 \V2/V2/V1/_0_  (.A1(\V2/V2/V1/c1 ),
    .A2(\V2/V2/V1/c2 ),
    .ZN(\V2/V2/V1/c3 ));
 AND2_X1 \V2/V2/V2/A1/M1/M1/_0_  (.A1(\V2/V2/V2/v2 [0]),
    .A2(\V2/V2/V2/v3 [0]),
    .ZN(\V2/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M1/M1/_1_  (.A(\V2/V2/V2/v2 [0]),
    .B(\V2/V2/V2/v3 [0]),
    .Z(\V2/V2/V2/A1/M1/s1 ));
 AND2_X1 \V2/V2/V2/A1/M1/M2/_0_  (.A1(\V2/V2/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M1/M2/_1_  (.A(\V2/V2/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/V2/s1 [0]));
 OR2_X1 \V2/V2/V2/A1/M1/_0_  (.A1(\V2/V2/V2/A1/M1/c1 ),
    .A2(\V2/V2/V2/A1/M1/c2 ),
    .ZN(\V2/V2/V2/A1/c1 ));
 AND2_X1 \V2/V2/V2/A1/M2/M1/_0_  (.A1(\V2/V2/V2/v2 [1]),
    .A2(\V2/V2/V2/v3 [1]),
    .ZN(\V2/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M2/M1/_1_  (.A(\V2/V2/V2/v2 [1]),
    .B(\V2/V2/V2/v3 [1]),
    .Z(\V2/V2/V2/A1/M2/s1 ));
 AND2_X1 \V2/V2/V2/A1/M2/M2/_0_  (.A1(\V2/V2/V2/A1/M2/s1 ),
    .A2(\V2/V2/V2/A1/c1 ),
    .ZN(\V2/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M2/M2/_1_  (.A(\V2/V2/V2/A1/M2/s1 ),
    .B(\V2/V2/V2/A1/c1 ),
    .Z(\V2/V2/V2/s1 [1]));
 OR2_X1 \V2/V2/V2/A1/M2/_0_  (.A1(\V2/V2/V2/A1/M2/c1 ),
    .A2(\V2/V2/V2/A1/M2/c2 ),
    .ZN(\V2/V2/V2/A1/c2 ));
 AND2_X1 \V2/V2/V2/A1/M3/M1/_0_  (.A1(\V2/V2/V2/v2 [2]),
    .A2(\V2/V2/V2/v3 [2]),
    .ZN(\V2/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M3/M1/_1_  (.A(\V2/V2/V2/v2 [2]),
    .B(\V2/V2/V2/v3 [2]),
    .Z(\V2/V2/V2/A1/M3/s1 ));
 AND2_X1 \V2/V2/V2/A1/M3/M2/_0_  (.A1(\V2/V2/V2/A1/M3/s1 ),
    .A2(\V2/V2/V2/A1/c2 ),
    .ZN(\V2/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M3/M2/_1_  (.A(\V2/V2/V2/A1/M3/s1 ),
    .B(\V2/V2/V2/A1/c2 ),
    .Z(\V2/V2/V2/s1 [2]));
 OR2_X1 \V2/V2/V2/A1/M3/_0_  (.A1(\V2/V2/V2/A1/M3/c1 ),
    .A2(\V2/V2/V2/A1/M3/c2 ),
    .ZN(\V2/V2/V2/A1/c3 ));
 AND2_X1 \V2/V2/V2/A1/M4/M1/_0_  (.A1(\V2/V2/V2/v2 [3]),
    .A2(\V2/V2/V2/v3 [3]),
    .ZN(\V2/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M4/M1/_1_  (.A(\V2/V2/V2/v2 [3]),
    .B(\V2/V2/V2/v3 [3]),
    .Z(\V2/V2/V2/A1/M4/s1 ));
 AND2_X1 \V2/V2/V2/A1/M4/M2/_0_  (.A1(\V2/V2/V2/A1/M4/s1 ),
    .A2(\V2/V2/V2/A1/c3 ),
    .ZN(\V2/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M4/M2/_1_  (.A(\V2/V2/V2/A1/M4/s1 ),
    .B(\V2/V2/V2/A1/c3 ),
    .Z(\V2/V2/V2/s1 [3]));
 OR2_X1 \V2/V2/V2/A1/M4/_0_  (.A1(\V2/V2/V2/A1/M4/c1 ),
    .A2(\V2/V2/V2/A1/M4/c2 ),
    .ZN(\V2/V2/V2/c1 ));
 AND2_X1 \V2/V2/V2/A2/M1/M1/_0_  (.A1(\V2/V2/V2/s1 [0]),
    .A2(\V2/V2/V2/v1 [2]),
    .ZN(\V2/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M1/M1/_1_  (.A(\V2/V2/V2/s1 [0]),
    .B(\V2/V2/V2/v1 [2]),
    .Z(\V2/V2/V2/A2/M1/s1 ));
 AND2_X1 \V2/V2/V2/A2/M1/M2/_0_  (.A1(\V2/V2/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M1/M2/_1_  (.A(\V2/V2/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v2 [2]));
 OR2_X1 \V2/V2/V2/A2/M1/_0_  (.A1(\V2/V2/V2/A2/M1/c1 ),
    .A2(\V2/V2/V2/A2/M1/c2 ),
    .ZN(\V2/V2/V2/A2/c1 ));
 AND2_X1 \V2/V2/V2/A2/M2/M1/_0_  (.A1(\V2/V2/V2/s1 [1]),
    .A2(\V2/V2/V2/v1 [3]),
    .ZN(\V2/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M2/M1/_1_  (.A(\V2/V2/V2/s1 [1]),
    .B(\V2/V2/V2/v1 [3]),
    .Z(\V2/V2/V2/A2/M2/s1 ));
 AND2_X1 \V2/V2/V2/A2/M2/M2/_0_  (.A1(\V2/V2/V2/A2/M2/s1 ),
    .A2(\V2/V2/V2/A2/c1 ),
    .ZN(\V2/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M2/M2/_1_  (.A(\V2/V2/V2/A2/M2/s1 ),
    .B(\V2/V2/V2/A2/c1 ),
    .Z(\V2/V2/v2 [3]));
 OR2_X1 \V2/V2/V2/A2/M2/_0_  (.A1(\V2/V2/V2/A2/M2/c1 ),
    .A2(\V2/V2/V2/A2/M2/c2 ),
    .ZN(\V2/V2/V2/A2/c2 ));
 AND2_X1 \V2/V2/V2/A2/M3/M1/_0_  (.A1(\V2/V2/V2/s1 [2]),
    .A2(ground),
    .ZN(\V2/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M3/M1/_1_  (.A(\V2/V2/V2/s1 [2]),
    .B(ground),
    .Z(\V2/V2/V2/A2/M3/s1 ));
 AND2_X1 \V2/V2/V2/A2/M3/M2/_0_  (.A1(\V2/V2/V2/A2/M3/s1 ),
    .A2(\V2/V2/V2/A2/c2 ),
    .ZN(\V2/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M3/M2/_1_  (.A(\V2/V2/V2/A2/M3/s1 ),
    .B(\V2/V2/V2/A2/c2 ),
    .Z(\V2/V2/V2/s2 [2]));
 OR2_X1 \V2/V2/V2/A2/M3/_0_  (.A1(\V2/V2/V2/A2/M3/c1 ),
    .A2(\V2/V2/V2/A2/M3/c2 ),
    .ZN(\V2/V2/V2/A2/c3 ));
 AND2_X1 \V2/V2/V2/A2/M4/M1/_0_  (.A1(\V2/V2/V2/s1 [3]),
    .A2(ground),
    .ZN(\V2/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M4/M1/_1_  (.A(\V2/V2/V2/s1 [3]),
    .B(ground),
    .Z(\V2/V2/V2/A2/M4/s1 ));
 AND2_X1 \V2/V2/V2/A2/M4/M2/_0_  (.A1(\V2/V2/V2/A2/M4/s1 ),
    .A2(\V2/V2/V2/A2/c3 ),
    .ZN(\V2/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M4/M2/_1_  (.A(\V2/V2/V2/A2/M4/s1 ),
    .B(\V2/V2/V2/A2/c3 ),
    .Z(\V2/V2/V2/s2 [3]));
 OR2_X1 \V2/V2/V2/A2/M4/_0_  (.A1(\V2/V2/V2/A2/M4/c1 ),
    .A2(\V2/V2/V2/A2/M4/c2 ),
    .ZN(\V2/V2/V2/c2 ));
 AND2_X1 \V2/V2/V2/A3/M1/M1/_0_  (.A1(\V2/V2/V2/v4 [0]),
    .A2(\V2/V2/V2/s2 [2]),
    .ZN(\V2/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M1/M1/_1_  (.A(\V2/V2/V2/v4 [0]),
    .B(\V2/V2/V2/s2 [2]),
    .Z(\V2/V2/V2/A3/M1/s1 ));
 AND2_X1 \V2/V2/V2/A3/M1/M2/_0_  (.A1(\V2/V2/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M1/M2/_1_  (.A(\V2/V2/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v2 [4]));
 OR2_X1 \V2/V2/V2/A3/M1/_0_  (.A1(\V2/V2/V2/A3/M1/c1 ),
    .A2(\V2/V2/V2/A3/M1/c2 ),
    .ZN(\V2/V2/V2/A3/c1 ));
 AND2_X1 \V2/V2/V2/A3/M2/M1/_0_  (.A1(\V2/V2/V2/v4 [1]),
    .A2(\V2/V2/V2/s2 [3]),
    .ZN(\V2/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M2/M1/_1_  (.A(\V2/V2/V2/v4 [1]),
    .B(\V2/V2/V2/s2 [3]),
    .Z(\V2/V2/V2/A3/M2/s1 ));
 AND2_X1 \V2/V2/V2/A3/M2/M2/_0_  (.A1(\V2/V2/V2/A3/M2/s1 ),
    .A2(\V2/V2/V2/A3/c1 ),
    .ZN(\V2/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M2/M2/_1_  (.A(\V2/V2/V2/A3/M2/s1 ),
    .B(\V2/V2/V2/A3/c1 ),
    .Z(\V2/V2/v2 [5]));
 OR2_X1 \V2/V2/V2/A3/M2/_0_  (.A1(\V2/V2/V2/A3/M2/c1 ),
    .A2(\V2/V2/V2/A3/M2/c2 ),
    .ZN(\V2/V2/V2/A3/c2 ));
 AND2_X1 \V2/V2/V2/A3/M3/M1/_0_  (.A1(\V2/V2/V2/v4 [2]),
    .A2(\V2/V2/V2/c3 ),
    .ZN(\V2/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M3/M1/_1_  (.A(\V2/V2/V2/v4 [2]),
    .B(\V2/V2/V2/c3 ),
    .Z(\V2/V2/V2/A3/M3/s1 ));
 AND2_X1 \V2/V2/V2/A3/M3/M2/_0_  (.A1(\V2/V2/V2/A3/M3/s1 ),
    .A2(\V2/V2/V2/A3/c2 ),
    .ZN(\V2/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M3/M2/_1_  (.A(\V2/V2/V2/A3/M3/s1 ),
    .B(\V2/V2/V2/A3/c2 ),
    .Z(\V2/V2/v2 [6]));
 OR2_X1 \V2/V2/V2/A3/M3/_0_  (.A1(\V2/V2/V2/A3/M3/c1 ),
    .A2(\V2/V2/V2/A3/M3/c2 ),
    .ZN(\V2/V2/V2/A3/c3 ));
 AND2_X1 \V2/V2/V2/A3/M4/M1/_0_  (.A1(\V2/V2/V2/v4 [3]),
    .A2(ground),
    .ZN(\V2/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M4/M1/_1_  (.A(\V2/V2/V2/v4 [3]),
    .B(ground),
    .Z(\V2/V2/V2/A3/M4/s1 ));
 AND2_X1 \V2/V2/V2/A3/M4/M2/_0_  (.A1(\V2/V2/V2/A3/M4/s1 ),
    .A2(\V2/V2/V2/A3/c3 ),
    .ZN(\V2/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M4/M2/_1_  (.A(\V2/V2/V2/A3/M4/s1 ),
    .B(\V2/V2/V2/A3/c3 ),
    .Z(\V2/V2/v2 [7]));
 OR2_X1 \V2/V2/V2/A3/M4/_0_  (.A1(\V2/V2/V2/A3/M4/c1 ),
    .A2(\V2/V2/V2/A3/M4/c2 ),
    .ZN(\V2/V2/V2/overflow ));
 AND2_X1 \V2/V2/V2/V1/HA1/_0_  (.A1(\V2/V2/V2/V1/w2 ),
    .A2(\V2/V2/V2/V1/w1 ),
    .ZN(\V2/V2/V2/V1/w4 ));
 XOR2_X2 \V2/V2/V2/V1/HA1/_1_  (.A(\V2/V2/V2/V1/w2 ),
    .B(\V2/V2/V2/V1/w1 ),
    .Z(\V2/V2/v2 [1]));
 AND2_X1 \V2/V2/V2/V1/HA2/_0_  (.A1(\V2/V2/V2/V1/w4 ),
    .A2(\V2/V2/V2/V1/w3 ),
    .ZN(\V2/V2/V2/v1 [3]));
 XOR2_X2 \V2/V2/V2/V1/HA2/_1_  (.A(\V2/V2/V2/V1/w4 ),
    .B(\V2/V2/V2/V1/w3 ),
    .Z(\V2/V2/V2/v1 [2]));
 AND2_X1 \V2/V2/V2/V1/_0_  (.A1(A[28]),
    .A2(B[0]),
    .ZN(\V2/V2/v2 [0]));
 AND2_X1 \V2/V2/V2/V1/_1_  (.A1(A[28]),
    .A2(B[1]),
    .ZN(\V2/V2/V2/V1/w1 ));
 AND2_X1 \V2/V2/V2/V1/_2_  (.A1(B[0]),
    .A2(A[29]),
    .ZN(\V2/V2/V2/V1/w2 ));
 AND2_X1 \V2/V2/V2/V1/_3_  (.A1(B[1]),
    .A2(A[29]),
    .ZN(\V2/V2/V2/V1/w3 ));
 AND2_X1 \V2/V2/V2/V2/HA1/_0_  (.A1(\V2/V2/V2/V2/w2 ),
    .A2(\V2/V2/V2/V2/w1 ),
    .ZN(\V2/V2/V2/V2/w4 ));
 XOR2_X2 \V2/V2/V2/V2/HA1/_1_  (.A(\V2/V2/V2/V2/w2 ),
    .B(\V2/V2/V2/V2/w1 ),
    .Z(\V2/V2/V2/v2 [1]));
 AND2_X1 \V2/V2/V2/V2/HA2/_0_  (.A1(\V2/V2/V2/V2/w4 ),
    .A2(\V2/V2/V2/V2/w3 ),
    .ZN(\V2/V2/V2/v2 [3]));
 XOR2_X2 \V2/V2/V2/V2/HA2/_1_  (.A(\V2/V2/V2/V2/w4 ),
    .B(\V2/V2/V2/V2/w3 ),
    .Z(\V2/V2/V2/v2 [2]));
 AND2_X1 \V2/V2/V2/V2/_0_  (.A1(A[30]),
    .A2(B[0]),
    .ZN(\V2/V2/V2/v2 [0]));
 AND2_X1 \V2/V2/V2/V2/_1_  (.A1(A[30]),
    .A2(B[1]),
    .ZN(\V2/V2/V2/V2/w1 ));
 AND2_X1 \V2/V2/V2/V2/_2_  (.A1(B[0]),
    .A2(A[31]),
    .ZN(\V2/V2/V2/V2/w2 ));
 AND2_X1 \V2/V2/V2/V2/_3_  (.A1(B[1]),
    .A2(A[31]),
    .ZN(\V2/V2/V2/V2/w3 ));
 AND2_X1 \V2/V2/V2/V3/HA1/_0_  (.A1(\V2/V2/V2/V3/w2 ),
    .A2(\V2/V2/V2/V3/w1 ),
    .ZN(\V2/V2/V2/V3/w4 ));
 XOR2_X2 \V2/V2/V2/V3/HA1/_1_  (.A(\V2/V2/V2/V3/w2 ),
    .B(\V2/V2/V2/V3/w1 ),
    .Z(\V2/V2/V2/v3 [1]));
 AND2_X1 \V2/V2/V2/V3/HA2/_0_  (.A1(\V2/V2/V2/V3/w4 ),
    .A2(\V2/V2/V2/V3/w3 ),
    .ZN(\V2/V2/V2/v3 [3]));
 XOR2_X2 \V2/V2/V2/V3/HA2/_1_  (.A(\V2/V2/V2/V3/w4 ),
    .B(\V2/V2/V2/V3/w3 ),
    .Z(\V2/V2/V2/v3 [2]));
 AND2_X1 \V2/V2/V2/V3/_0_  (.A1(A[28]),
    .A2(B[2]),
    .ZN(\V2/V2/V2/v3 [0]));
 AND2_X1 \V2/V2/V2/V3/_1_  (.A1(A[28]),
    .A2(B[3]),
    .ZN(\V2/V2/V2/V3/w1 ));
 AND2_X1 \V2/V2/V2/V3/_2_  (.A1(B[2]),
    .A2(A[29]),
    .ZN(\V2/V2/V2/V3/w2 ));
 AND2_X1 \V2/V2/V2/V3/_3_  (.A1(B[3]),
    .A2(A[29]),
    .ZN(\V2/V2/V2/V3/w3 ));
 AND2_X1 \V2/V2/V2/V4/HA1/_0_  (.A1(\V2/V2/V2/V4/w2 ),
    .A2(\V2/V2/V2/V4/w1 ),
    .ZN(\V2/V2/V2/V4/w4 ));
 XOR2_X2 \V2/V2/V2/V4/HA1/_1_  (.A(\V2/V2/V2/V4/w2 ),
    .B(\V2/V2/V2/V4/w1 ),
    .Z(\V2/V2/V2/v4 [1]));
 AND2_X1 \V2/V2/V2/V4/HA2/_0_  (.A1(\V2/V2/V2/V4/w4 ),
    .A2(\V2/V2/V2/V4/w3 ),
    .ZN(\V2/V2/V2/v4 [3]));
 XOR2_X2 \V2/V2/V2/V4/HA2/_1_  (.A(\V2/V2/V2/V4/w4 ),
    .B(\V2/V2/V2/V4/w3 ),
    .Z(\V2/V2/V2/v4 [2]));
 AND2_X1 \V2/V2/V2/V4/_0_  (.A1(A[30]),
    .A2(B[2]),
    .ZN(\V2/V2/V2/v4 [0]));
 AND2_X1 \V2/V2/V2/V4/_1_  (.A1(A[30]),
    .A2(B[3]),
    .ZN(\V2/V2/V2/V4/w1 ));
 AND2_X1 \V2/V2/V2/V4/_2_  (.A1(B[2]),
    .A2(A[31]),
    .ZN(\V2/V2/V2/V4/w2 ));
 AND2_X1 \V2/V2/V2/V4/_3_  (.A1(B[3]),
    .A2(A[31]),
    .ZN(\V2/V2/V2/V4/w3 ));
 OR2_X1 \V2/V2/V2/_0_  (.A1(\V2/V2/V2/c1 ),
    .A2(\V2/V2/V2/c2 ),
    .ZN(\V2/V2/V2/c3 ));
 AND2_X1 \V2/V2/V3/A1/M1/M1/_0_  (.A1(\V2/V2/V3/v2 [0]),
    .A2(\V2/V2/V3/v3 [0]),
    .ZN(\V2/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M1/M1/_1_  (.A(\V2/V2/V3/v2 [0]),
    .B(\V2/V2/V3/v3 [0]),
    .Z(\V2/V2/V3/A1/M1/s1 ));
 AND2_X1 \V2/V2/V3/A1/M1/M2/_0_  (.A1(\V2/V2/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M1/M2/_1_  (.A(\V2/V2/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/V3/s1 [0]));
 OR2_X1 \V2/V2/V3/A1/M1/_0_  (.A1(\V2/V2/V3/A1/M1/c1 ),
    .A2(\V2/V2/V3/A1/M1/c2 ),
    .ZN(\V2/V2/V3/A1/c1 ));
 AND2_X1 \V2/V2/V3/A1/M2/M1/_0_  (.A1(\V2/V2/V3/v2 [1]),
    .A2(\V2/V2/V3/v3 [1]),
    .ZN(\V2/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M2/M1/_1_  (.A(\V2/V2/V3/v2 [1]),
    .B(\V2/V2/V3/v3 [1]),
    .Z(\V2/V2/V3/A1/M2/s1 ));
 AND2_X1 \V2/V2/V3/A1/M2/M2/_0_  (.A1(\V2/V2/V3/A1/M2/s1 ),
    .A2(\V2/V2/V3/A1/c1 ),
    .ZN(\V2/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M2/M2/_1_  (.A(\V2/V2/V3/A1/M2/s1 ),
    .B(\V2/V2/V3/A1/c1 ),
    .Z(\V2/V2/V3/s1 [1]));
 OR2_X1 \V2/V2/V3/A1/M2/_0_  (.A1(\V2/V2/V3/A1/M2/c1 ),
    .A2(\V2/V2/V3/A1/M2/c2 ),
    .ZN(\V2/V2/V3/A1/c2 ));
 AND2_X1 \V2/V2/V3/A1/M3/M1/_0_  (.A1(\V2/V2/V3/v2 [2]),
    .A2(\V2/V2/V3/v3 [2]),
    .ZN(\V2/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M3/M1/_1_  (.A(\V2/V2/V3/v2 [2]),
    .B(\V2/V2/V3/v3 [2]),
    .Z(\V2/V2/V3/A1/M3/s1 ));
 AND2_X1 \V2/V2/V3/A1/M3/M2/_0_  (.A1(\V2/V2/V3/A1/M3/s1 ),
    .A2(\V2/V2/V3/A1/c2 ),
    .ZN(\V2/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M3/M2/_1_  (.A(\V2/V2/V3/A1/M3/s1 ),
    .B(\V2/V2/V3/A1/c2 ),
    .Z(\V2/V2/V3/s1 [2]));
 OR2_X1 \V2/V2/V3/A1/M3/_0_  (.A1(\V2/V2/V3/A1/M3/c1 ),
    .A2(\V2/V2/V3/A1/M3/c2 ),
    .ZN(\V2/V2/V3/A1/c3 ));
 AND2_X1 \V2/V2/V3/A1/M4/M1/_0_  (.A1(\V2/V2/V3/v2 [3]),
    .A2(\V2/V2/V3/v3 [3]),
    .ZN(\V2/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M4/M1/_1_  (.A(\V2/V2/V3/v2 [3]),
    .B(\V2/V2/V3/v3 [3]),
    .Z(\V2/V2/V3/A1/M4/s1 ));
 AND2_X1 \V2/V2/V3/A1/M4/M2/_0_  (.A1(\V2/V2/V3/A1/M4/s1 ),
    .A2(\V2/V2/V3/A1/c3 ),
    .ZN(\V2/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M4/M2/_1_  (.A(\V2/V2/V3/A1/M4/s1 ),
    .B(\V2/V2/V3/A1/c3 ),
    .Z(\V2/V2/V3/s1 [3]));
 OR2_X1 \V2/V2/V3/A1/M4/_0_  (.A1(\V2/V2/V3/A1/M4/c1 ),
    .A2(\V2/V2/V3/A1/M4/c2 ),
    .ZN(\V2/V2/V3/c1 ));
 AND2_X1 \V2/V2/V3/A2/M1/M1/_0_  (.A1(\V2/V2/V3/s1 [0]),
    .A2(\V2/V2/V3/v1 [2]),
    .ZN(\V2/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M1/M1/_1_  (.A(\V2/V2/V3/s1 [0]),
    .B(\V2/V2/V3/v1 [2]),
    .Z(\V2/V2/V3/A2/M1/s1 ));
 AND2_X1 \V2/V2/V3/A2/M1/M2/_0_  (.A1(\V2/V2/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M1/M2/_1_  (.A(\V2/V2/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v3 [2]));
 OR2_X1 \V2/V2/V3/A2/M1/_0_  (.A1(\V2/V2/V3/A2/M1/c1 ),
    .A2(\V2/V2/V3/A2/M1/c2 ),
    .ZN(\V2/V2/V3/A2/c1 ));
 AND2_X1 \V2/V2/V3/A2/M2/M1/_0_  (.A1(\V2/V2/V3/s1 [1]),
    .A2(\V2/V2/V3/v1 [3]),
    .ZN(\V2/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M2/M1/_1_  (.A(\V2/V2/V3/s1 [1]),
    .B(\V2/V2/V3/v1 [3]),
    .Z(\V2/V2/V3/A2/M2/s1 ));
 AND2_X1 \V2/V2/V3/A2/M2/M2/_0_  (.A1(\V2/V2/V3/A2/M2/s1 ),
    .A2(\V2/V2/V3/A2/c1 ),
    .ZN(\V2/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M2/M2/_1_  (.A(\V2/V2/V3/A2/M2/s1 ),
    .B(\V2/V2/V3/A2/c1 ),
    .Z(\V2/V2/v3 [3]));
 OR2_X1 \V2/V2/V3/A2/M2/_0_  (.A1(\V2/V2/V3/A2/M2/c1 ),
    .A2(\V2/V2/V3/A2/M2/c2 ),
    .ZN(\V2/V2/V3/A2/c2 ));
 AND2_X1 \V2/V2/V3/A2/M3/M1/_0_  (.A1(\V2/V2/V3/s1 [2]),
    .A2(ground),
    .ZN(\V2/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M3/M1/_1_  (.A(\V2/V2/V3/s1 [2]),
    .B(ground),
    .Z(\V2/V2/V3/A2/M3/s1 ));
 AND2_X1 \V2/V2/V3/A2/M3/M2/_0_  (.A1(\V2/V2/V3/A2/M3/s1 ),
    .A2(\V2/V2/V3/A2/c2 ),
    .ZN(\V2/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M3/M2/_1_  (.A(\V2/V2/V3/A2/M3/s1 ),
    .B(\V2/V2/V3/A2/c2 ),
    .Z(\V2/V2/V3/s2 [2]));
 OR2_X1 \V2/V2/V3/A2/M3/_0_  (.A1(\V2/V2/V3/A2/M3/c1 ),
    .A2(\V2/V2/V3/A2/M3/c2 ),
    .ZN(\V2/V2/V3/A2/c3 ));
 AND2_X1 \V2/V2/V3/A2/M4/M1/_0_  (.A1(\V2/V2/V3/s1 [3]),
    .A2(ground),
    .ZN(\V2/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M4/M1/_1_  (.A(\V2/V2/V3/s1 [3]),
    .B(ground),
    .Z(\V2/V2/V3/A2/M4/s1 ));
 AND2_X1 \V2/V2/V3/A2/M4/M2/_0_  (.A1(\V2/V2/V3/A2/M4/s1 ),
    .A2(\V2/V2/V3/A2/c3 ),
    .ZN(\V2/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M4/M2/_1_  (.A(\V2/V2/V3/A2/M4/s1 ),
    .B(\V2/V2/V3/A2/c3 ),
    .Z(\V2/V2/V3/s2 [3]));
 OR2_X1 \V2/V2/V3/A2/M4/_0_  (.A1(\V2/V2/V3/A2/M4/c1 ),
    .A2(\V2/V2/V3/A2/M4/c2 ),
    .ZN(\V2/V2/V3/c2 ));
 AND2_X1 \V2/V2/V3/A3/M1/M1/_0_  (.A1(\V2/V2/V3/v4 [0]),
    .A2(\V2/V2/V3/s2 [2]),
    .ZN(\V2/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M1/M1/_1_  (.A(\V2/V2/V3/v4 [0]),
    .B(\V2/V2/V3/s2 [2]),
    .Z(\V2/V2/V3/A3/M1/s1 ));
 AND2_X1 \V2/V2/V3/A3/M1/M2/_0_  (.A1(\V2/V2/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M1/M2/_1_  (.A(\V2/V2/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v3 [4]));
 OR2_X1 \V2/V2/V3/A3/M1/_0_  (.A1(\V2/V2/V3/A3/M1/c1 ),
    .A2(\V2/V2/V3/A3/M1/c2 ),
    .ZN(\V2/V2/V3/A3/c1 ));
 AND2_X1 \V2/V2/V3/A3/M2/M1/_0_  (.A1(\V2/V2/V3/v4 [1]),
    .A2(\V2/V2/V3/s2 [3]),
    .ZN(\V2/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M2/M1/_1_  (.A(\V2/V2/V3/v4 [1]),
    .B(\V2/V2/V3/s2 [3]),
    .Z(\V2/V2/V3/A3/M2/s1 ));
 AND2_X1 \V2/V2/V3/A3/M2/M2/_0_  (.A1(\V2/V2/V3/A3/M2/s1 ),
    .A2(\V2/V2/V3/A3/c1 ),
    .ZN(\V2/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M2/M2/_1_  (.A(\V2/V2/V3/A3/M2/s1 ),
    .B(\V2/V2/V3/A3/c1 ),
    .Z(\V2/V2/v3 [5]));
 OR2_X1 \V2/V2/V3/A3/M2/_0_  (.A1(\V2/V2/V3/A3/M2/c1 ),
    .A2(\V2/V2/V3/A3/M2/c2 ),
    .ZN(\V2/V2/V3/A3/c2 ));
 AND2_X1 \V2/V2/V3/A3/M3/M1/_0_  (.A1(\V2/V2/V3/v4 [2]),
    .A2(\V2/V2/V3/c3 ),
    .ZN(\V2/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M3/M1/_1_  (.A(\V2/V2/V3/v4 [2]),
    .B(\V2/V2/V3/c3 ),
    .Z(\V2/V2/V3/A3/M3/s1 ));
 AND2_X1 \V2/V2/V3/A3/M3/M2/_0_  (.A1(\V2/V2/V3/A3/M3/s1 ),
    .A2(\V2/V2/V3/A3/c2 ),
    .ZN(\V2/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M3/M2/_1_  (.A(\V2/V2/V3/A3/M3/s1 ),
    .B(\V2/V2/V3/A3/c2 ),
    .Z(\V2/V2/v3 [6]));
 OR2_X1 \V2/V2/V3/A3/M3/_0_  (.A1(\V2/V2/V3/A3/M3/c1 ),
    .A2(\V2/V2/V3/A3/M3/c2 ),
    .ZN(\V2/V2/V3/A3/c3 ));
 AND2_X1 \V2/V2/V3/A3/M4/M1/_0_  (.A1(\V2/V2/V3/v4 [3]),
    .A2(ground),
    .ZN(\V2/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M4/M1/_1_  (.A(\V2/V2/V3/v4 [3]),
    .B(ground),
    .Z(\V2/V2/V3/A3/M4/s1 ));
 AND2_X1 \V2/V2/V3/A3/M4/M2/_0_  (.A1(\V2/V2/V3/A3/M4/s1 ),
    .A2(\V2/V2/V3/A3/c3 ),
    .ZN(\V2/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M4/M2/_1_  (.A(\V2/V2/V3/A3/M4/s1 ),
    .B(\V2/V2/V3/A3/c3 ),
    .Z(\V2/V2/v3 [7]));
 OR2_X1 \V2/V2/V3/A3/M4/_0_  (.A1(\V2/V2/V3/A3/M4/c1 ),
    .A2(\V2/V2/V3/A3/M4/c2 ),
    .ZN(\V2/V2/V3/overflow ));
 AND2_X1 \V2/V2/V3/V1/HA1/_0_  (.A1(\V2/V2/V3/V1/w2 ),
    .A2(\V2/V2/V3/V1/w1 ),
    .ZN(\V2/V2/V3/V1/w4 ));
 XOR2_X2 \V2/V2/V3/V1/HA1/_1_  (.A(\V2/V2/V3/V1/w2 ),
    .B(\V2/V2/V3/V1/w1 ),
    .Z(\V2/V2/v3 [1]));
 AND2_X1 \V2/V2/V3/V1/HA2/_0_  (.A1(\V2/V2/V3/V1/w4 ),
    .A2(\V2/V2/V3/V1/w3 ),
    .ZN(\V2/V2/V3/v1 [3]));
 XOR2_X2 \V2/V2/V3/V1/HA2/_1_  (.A(\V2/V2/V3/V1/w4 ),
    .B(\V2/V2/V3/V1/w3 ),
    .Z(\V2/V2/V3/v1 [2]));
 AND2_X1 \V2/V2/V3/V1/_0_  (.A1(A[24]),
    .A2(B[4]),
    .ZN(\V2/V2/v3 [0]));
 AND2_X1 \V2/V2/V3/V1/_1_  (.A1(A[24]),
    .A2(B[5]),
    .ZN(\V2/V2/V3/V1/w1 ));
 AND2_X1 \V2/V2/V3/V1/_2_  (.A1(B[4]),
    .A2(A[25]),
    .ZN(\V2/V2/V3/V1/w2 ));
 AND2_X1 \V2/V2/V3/V1/_3_  (.A1(B[5]),
    .A2(A[25]),
    .ZN(\V2/V2/V3/V1/w3 ));
 AND2_X1 \V2/V2/V3/V2/HA1/_0_  (.A1(\V2/V2/V3/V2/w2 ),
    .A2(\V2/V2/V3/V2/w1 ),
    .ZN(\V2/V2/V3/V2/w4 ));
 XOR2_X2 \V2/V2/V3/V2/HA1/_1_  (.A(\V2/V2/V3/V2/w2 ),
    .B(\V2/V2/V3/V2/w1 ),
    .Z(\V2/V2/V3/v2 [1]));
 AND2_X1 \V2/V2/V3/V2/HA2/_0_  (.A1(\V2/V2/V3/V2/w4 ),
    .A2(\V2/V2/V3/V2/w3 ),
    .ZN(\V2/V2/V3/v2 [3]));
 XOR2_X2 \V2/V2/V3/V2/HA2/_1_  (.A(\V2/V2/V3/V2/w4 ),
    .B(\V2/V2/V3/V2/w3 ),
    .Z(\V2/V2/V3/v2 [2]));
 AND2_X1 \V2/V2/V3/V2/_0_  (.A1(A[26]),
    .A2(B[4]),
    .ZN(\V2/V2/V3/v2 [0]));
 AND2_X1 \V2/V2/V3/V2/_1_  (.A1(A[26]),
    .A2(B[5]),
    .ZN(\V2/V2/V3/V2/w1 ));
 AND2_X1 \V2/V2/V3/V2/_2_  (.A1(B[4]),
    .A2(A[27]),
    .ZN(\V2/V2/V3/V2/w2 ));
 AND2_X1 \V2/V2/V3/V2/_3_  (.A1(B[5]),
    .A2(A[27]),
    .ZN(\V2/V2/V3/V2/w3 ));
 AND2_X1 \V2/V2/V3/V3/HA1/_0_  (.A1(\V2/V2/V3/V3/w2 ),
    .A2(\V2/V2/V3/V3/w1 ),
    .ZN(\V2/V2/V3/V3/w4 ));
 XOR2_X2 \V2/V2/V3/V3/HA1/_1_  (.A(\V2/V2/V3/V3/w2 ),
    .B(\V2/V2/V3/V3/w1 ),
    .Z(\V2/V2/V3/v3 [1]));
 AND2_X1 \V2/V2/V3/V3/HA2/_0_  (.A1(\V2/V2/V3/V3/w4 ),
    .A2(\V2/V2/V3/V3/w3 ),
    .ZN(\V2/V2/V3/v3 [3]));
 XOR2_X2 \V2/V2/V3/V3/HA2/_1_  (.A(\V2/V2/V3/V3/w4 ),
    .B(\V2/V2/V3/V3/w3 ),
    .Z(\V2/V2/V3/v3 [2]));
 AND2_X1 \V2/V2/V3/V3/_0_  (.A1(A[24]),
    .A2(B[6]),
    .ZN(\V2/V2/V3/v3 [0]));
 AND2_X1 \V2/V2/V3/V3/_1_  (.A1(A[24]),
    .A2(B[7]),
    .ZN(\V2/V2/V3/V3/w1 ));
 AND2_X1 \V2/V2/V3/V3/_2_  (.A1(B[6]),
    .A2(A[25]),
    .ZN(\V2/V2/V3/V3/w2 ));
 AND2_X1 \V2/V2/V3/V3/_3_  (.A1(B[7]),
    .A2(A[25]),
    .ZN(\V2/V2/V3/V3/w3 ));
 AND2_X1 \V2/V2/V3/V4/HA1/_0_  (.A1(\V2/V2/V3/V4/w2 ),
    .A2(\V2/V2/V3/V4/w1 ),
    .ZN(\V2/V2/V3/V4/w4 ));
 XOR2_X2 \V2/V2/V3/V4/HA1/_1_  (.A(\V2/V2/V3/V4/w2 ),
    .B(\V2/V2/V3/V4/w1 ),
    .Z(\V2/V2/V3/v4 [1]));
 AND2_X1 \V2/V2/V3/V4/HA2/_0_  (.A1(\V2/V2/V3/V4/w4 ),
    .A2(\V2/V2/V3/V4/w3 ),
    .ZN(\V2/V2/V3/v4 [3]));
 XOR2_X2 \V2/V2/V3/V4/HA2/_1_  (.A(\V2/V2/V3/V4/w4 ),
    .B(\V2/V2/V3/V4/w3 ),
    .Z(\V2/V2/V3/v4 [2]));
 AND2_X1 \V2/V2/V3/V4/_0_  (.A1(A[26]),
    .A2(B[6]),
    .ZN(\V2/V2/V3/v4 [0]));
 AND2_X1 \V2/V2/V3/V4/_1_  (.A1(A[26]),
    .A2(B[7]),
    .ZN(\V2/V2/V3/V4/w1 ));
 AND2_X1 \V2/V2/V3/V4/_2_  (.A1(B[6]),
    .A2(A[27]),
    .ZN(\V2/V2/V3/V4/w2 ));
 AND2_X1 \V2/V2/V3/V4/_3_  (.A1(B[7]),
    .A2(A[27]),
    .ZN(\V2/V2/V3/V4/w3 ));
 OR2_X1 \V2/V2/V3/_0_  (.A1(\V2/V2/V3/c1 ),
    .A2(\V2/V2/V3/c2 ),
    .ZN(\V2/V2/V3/c3 ));
 AND2_X1 \V2/V2/V4/A1/M1/M1/_0_  (.A1(\V2/V2/V4/v2 [0]),
    .A2(\V2/V2/V4/v3 [0]),
    .ZN(\V2/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M1/M1/_1_  (.A(\V2/V2/V4/v2 [0]),
    .B(\V2/V2/V4/v3 [0]),
    .Z(\V2/V2/V4/A1/M1/s1 ));
 AND2_X1 \V2/V2/V4/A1/M1/M2/_0_  (.A1(\V2/V2/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M1/M2/_1_  (.A(\V2/V2/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/V4/s1 [0]));
 OR2_X1 \V2/V2/V4/A1/M1/_0_  (.A1(\V2/V2/V4/A1/M1/c1 ),
    .A2(\V2/V2/V4/A1/M1/c2 ),
    .ZN(\V2/V2/V4/A1/c1 ));
 AND2_X1 \V2/V2/V4/A1/M2/M1/_0_  (.A1(\V2/V2/V4/v2 [1]),
    .A2(\V2/V2/V4/v3 [1]),
    .ZN(\V2/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M2/M1/_1_  (.A(\V2/V2/V4/v2 [1]),
    .B(\V2/V2/V4/v3 [1]),
    .Z(\V2/V2/V4/A1/M2/s1 ));
 AND2_X1 \V2/V2/V4/A1/M2/M2/_0_  (.A1(\V2/V2/V4/A1/M2/s1 ),
    .A2(\V2/V2/V4/A1/c1 ),
    .ZN(\V2/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M2/M2/_1_  (.A(\V2/V2/V4/A1/M2/s1 ),
    .B(\V2/V2/V4/A1/c1 ),
    .Z(\V2/V2/V4/s1 [1]));
 OR2_X1 \V2/V2/V4/A1/M2/_0_  (.A1(\V2/V2/V4/A1/M2/c1 ),
    .A2(\V2/V2/V4/A1/M2/c2 ),
    .ZN(\V2/V2/V4/A1/c2 ));
 AND2_X1 \V2/V2/V4/A1/M3/M1/_0_  (.A1(\V2/V2/V4/v2 [2]),
    .A2(\V2/V2/V4/v3 [2]),
    .ZN(\V2/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M3/M1/_1_  (.A(\V2/V2/V4/v2 [2]),
    .B(\V2/V2/V4/v3 [2]),
    .Z(\V2/V2/V4/A1/M3/s1 ));
 AND2_X1 \V2/V2/V4/A1/M3/M2/_0_  (.A1(\V2/V2/V4/A1/M3/s1 ),
    .A2(\V2/V2/V4/A1/c2 ),
    .ZN(\V2/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M3/M2/_1_  (.A(\V2/V2/V4/A1/M3/s1 ),
    .B(\V2/V2/V4/A1/c2 ),
    .Z(\V2/V2/V4/s1 [2]));
 OR2_X1 \V2/V2/V4/A1/M3/_0_  (.A1(\V2/V2/V4/A1/M3/c1 ),
    .A2(\V2/V2/V4/A1/M3/c2 ),
    .ZN(\V2/V2/V4/A1/c3 ));
 AND2_X1 \V2/V2/V4/A1/M4/M1/_0_  (.A1(\V2/V2/V4/v2 [3]),
    .A2(\V2/V2/V4/v3 [3]),
    .ZN(\V2/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M4/M1/_1_  (.A(\V2/V2/V4/v2 [3]),
    .B(\V2/V2/V4/v3 [3]),
    .Z(\V2/V2/V4/A1/M4/s1 ));
 AND2_X1 \V2/V2/V4/A1/M4/M2/_0_  (.A1(\V2/V2/V4/A1/M4/s1 ),
    .A2(\V2/V2/V4/A1/c3 ),
    .ZN(\V2/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M4/M2/_1_  (.A(\V2/V2/V4/A1/M4/s1 ),
    .B(\V2/V2/V4/A1/c3 ),
    .Z(\V2/V2/V4/s1 [3]));
 OR2_X1 \V2/V2/V4/A1/M4/_0_  (.A1(\V2/V2/V4/A1/M4/c1 ),
    .A2(\V2/V2/V4/A1/M4/c2 ),
    .ZN(\V2/V2/V4/c1 ));
 AND2_X1 \V2/V2/V4/A2/M1/M1/_0_  (.A1(\V2/V2/V4/s1 [0]),
    .A2(\V2/V2/V4/v1 [2]),
    .ZN(\V2/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M1/M1/_1_  (.A(\V2/V2/V4/s1 [0]),
    .B(\V2/V2/V4/v1 [2]),
    .Z(\V2/V2/V4/A2/M1/s1 ));
 AND2_X1 \V2/V2/V4/A2/M1/M2/_0_  (.A1(\V2/V2/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M1/M2/_1_  (.A(\V2/V2/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v4 [2]));
 OR2_X1 \V2/V2/V4/A2/M1/_0_  (.A1(\V2/V2/V4/A2/M1/c1 ),
    .A2(\V2/V2/V4/A2/M1/c2 ),
    .ZN(\V2/V2/V4/A2/c1 ));
 AND2_X1 \V2/V2/V4/A2/M2/M1/_0_  (.A1(\V2/V2/V4/s1 [1]),
    .A2(\V2/V2/V4/v1 [3]),
    .ZN(\V2/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M2/M1/_1_  (.A(\V2/V2/V4/s1 [1]),
    .B(\V2/V2/V4/v1 [3]),
    .Z(\V2/V2/V4/A2/M2/s1 ));
 AND2_X1 \V2/V2/V4/A2/M2/M2/_0_  (.A1(\V2/V2/V4/A2/M2/s1 ),
    .A2(\V2/V2/V4/A2/c1 ),
    .ZN(\V2/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M2/M2/_1_  (.A(\V2/V2/V4/A2/M2/s1 ),
    .B(\V2/V2/V4/A2/c1 ),
    .Z(\V2/V2/v4 [3]));
 OR2_X1 \V2/V2/V4/A2/M2/_0_  (.A1(\V2/V2/V4/A2/M2/c1 ),
    .A2(\V2/V2/V4/A2/M2/c2 ),
    .ZN(\V2/V2/V4/A2/c2 ));
 AND2_X1 \V2/V2/V4/A2/M3/M1/_0_  (.A1(\V2/V2/V4/s1 [2]),
    .A2(ground),
    .ZN(\V2/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M3/M1/_1_  (.A(\V2/V2/V4/s1 [2]),
    .B(ground),
    .Z(\V2/V2/V4/A2/M3/s1 ));
 AND2_X1 \V2/V2/V4/A2/M3/M2/_0_  (.A1(\V2/V2/V4/A2/M3/s1 ),
    .A2(\V2/V2/V4/A2/c2 ),
    .ZN(\V2/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M3/M2/_1_  (.A(\V2/V2/V4/A2/M3/s1 ),
    .B(\V2/V2/V4/A2/c2 ),
    .Z(\V2/V2/V4/s2 [2]));
 OR2_X1 \V2/V2/V4/A2/M3/_0_  (.A1(\V2/V2/V4/A2/M3/c1 ),
    .A2(\V2/V2/V4/A2/M3/c2 ),
    .ZN(\V2/V2/V4/A2/c3 ));
 AND2_X1 \V2/V2/V4/A2/M4/M1/_0_  (.A1(\V2/V2/V4/s1 [3]),
    .A2(ground),
    .ZN(\V2/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M4/M1/_1_  (.A(\V2/V2/V4/s1 [3]),
    .B(ground),
    .Z(\V2/V2/V4/A2/M4/s1 ));
 AND2_X1 \V2/V2/V4/A2/M4/M2/_0_  (.A1(\V2/V2/V4/A2/M4/s1 ),
    .A2(\V2/V2/V4/A2/c3 ),
    .ZN(\V2/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M4/M2/_1_  (.A(\V2/V2/V4/A2/M4/s1 ),
    .B(\V2/V2/V4/A2/c3 ),
    .Z(\V2/V2/V4/s2 [3]));
 OR2_X1 \V2/V2/V4/A2/M4/_0_  (.A1(\V2/V2/V4/A2/M4/c1 ),
    .A2(\V2/V2/V4/A2/M4/c2 ),
    .ZN(\V2/V2/V4/c2 ));
 AND2_X1 \V2/V2/V4/A3/M1/M1/_0_  (.A1(\V2/V2/V4/v4 [0]),
    .A2(\V2/V2/V4/s2 [2]),
    .ZN(\V2/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M1/M1/_1_  (.A(\V2/V2/V4/v4 [0]),
    .B(\V2/V2/V4/s2 [2]),
    .Z(\V2/V2/V4/A3/M1/s1 ));
 AND2_X1 \V2/V2/V4/A3/M1/M2/_0_  (.A1(\V2/V2/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M1/M2/_1_  (.A(\V2/V2/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V2/v4 [4]));
 OR2_X1 \V2/V2/V4/A3/M1/_0_  (.A1(\V2/V2/V4/A3/M1/c1 ),
    .A2(\V2/V2/V4/A3/M1/c2 ),
    .ZN(\V2/V2/V4/A3/c1 ));
 AND2_X1 \V2/V2/V4/A3/M2/M1/_0_  (.A1(\V2/V2/V4/v4 [1]),
    .A2(\V2/V2/V4/s2 [3]),
    .ZN(\V2/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M2/M1/_1_  (.A(\V2/V2/V4/v4 [1]),
    .B(\V2/V2/V4/s2 [3]),
    .Z(\V2/V2/V4/A3/M2/s1 ));
 AND2_X1 \V2/V2/V4/A3/M2/M2/_0_  (.A1(\V2/V2/V4/A3/M2/s1 ),
    .A2(\V2/V2/V4/A3/c1 ),
    .ZN(\V2/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M2/M2/_1_  (.A(\V2/V2/V4/A3/M2/s1 ),
    .B(\V2/V2/V4/A3/c1 ),
    .Z(\V2/V2/v4 [5]));
 OR2_X1 \V2/V2/V4/A3/M2/_0_  (.A1(\V2/V2/V4/A3/M2/c1 ),
    .A2(\V2/V2/V4/A3/M2/c2 ),
    .ZN(\V2/V2/V4/A3/c2 ));
 AND2_X1 \V2/V2/V4/A3/M3/M1/_0_  (.A1(\V2/V2/V4/v4 [2]),
    .A2(\V2/V2/V4/c3 ),
    .ZN(\V2/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M3/M1/_1_  (.A(\V2/V2/V4/v4 [2]),
    .B(\V2/V2/V4/c3 ),
    .Z(\V2/V2/V4/A3/M3/s1 ));
 AND2_X1 \V2/V2/V4/A3/M3/M2/_0_  (.A1(\V2/V2/V4/A3/M3/s1 ),
    .A2(\V2/V2/V4/A3/c2 ),
    .ZN(\V2/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M3/M2/_1_  (.A(\V2/V2/V4/A3/M3/s1 ),
    .B(\V2/V2/V4/A3/c2 ),
    .Z(\V2/V2/v4 [6]));
 OR2_X1 \V2/V2/V4/A3/M3/_0_  (.A1(\V2/V2/V4/A3/M3/c1 ),
    .A2(\V2/V2/V4/A3/M3/c2 ),
    .ZN(\V2/V2/V4/A3/c3 ));
 AND2_X1 \V2/V2/V4/A3/M4/M1/_0_  (.A1(\V2/V2/V4/v4 [3]),
    .A2(ground),
    .ZN(\V2/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M4/M1/_1_  (.A(\V2/V2/V4/v4 [3]),
    .B(ground),
    .Z(\V2/V2/V4/A3/M4/s1 ));
 AND2_X1 \V2/V2/V4/A3/M4/M2/_0_  (.A1(\V2/V2/V4/A3/M4/s1 ),
    .A2(\V2/V2/V4/A3/c3 ),
    .ZN(\V2/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M4/M2/_1_  (.A(\V2/V2/V4/A3/M4/s1 ),
    .B(\V2/V2/V4/A3/c3 ),
    .Z(\V2/V2/v4 [7]));
 OR2_X1 \V2/V2/V4/A3/M4/_0_  (.A1(\V2/V2/V4/A3/M4/c1 ),
    .A2(\V2/V2/V4/A3/M4/c2 ),
    .ZN(\V2/V2/V4/overflow ));
 AND2_X1 \V2/V2/V4/V1/HA1/_0_  (.A1(\V2/V2/V4/V1/w2 ),
    .A2(\V2/V2/V4/V1/w1 ),
    .ZN(\V2/V2/V4/V1/w4 ));
 XOR2_X2 \V2/V2/V4/V1/HA1/_1_  (.A(\V2/V2/V4/V1/w2 ),
    .B(\V2/V2/V4/V1/w1 ),
    .Z(\V2/V2/v4 [1]));
 AND2_X1 \V2/V2/V4/V1/HA2/_0_  (.A1(\V2/V2/V4/V1/w4 ),
    .A2(\V2/V2/V4/V1/w3 ),
    .ZN(\V2/V2/V4/v1 [3]));
 XOR2_X2 \V2/V2/V4/V1/HA2/_1_  (.A(\V2/V2/V4/V1/w4 ),
    .B(\V2/V2/V4/V1/w3 ),
    .Z(\V2/V2/V4/v1 [2]));
 AND2_X1 \V2/V2/V4/V1/_0_  (.A1(A[28]),
    .A2(B[4]),
    .ZN(\V2/V2/v4 [0]));
 AND2_X1 \V2/V2/V4/V1/_1_  (.A1(A[28]),
    .A2(B[5]),
    .ZN(\V2/V2/V4/V1/w1 ));
 AND2_X1 \V2/V2/V4/V1/_2_  (.A1(B[4]),
    .A2(A[29]),
    .ZN(\V2/V2/V4/V1/w2 ));
 AND2_X1 \V2/V2/V4/V1/_3_  (.A1(B[5]),
    .A2(A[29]),
    .ZN(\V2/V2/V4/V1/w3 ));
 AND2_X1 \V2/V2/V4/V2/HA1/_0_  (.A1(\V2/V2/V4/V2/w2 ),
    .A2(\V2/V2/V4/V2/w1 ),
    .ZN(\V2/V2/V4/V2/w4 ));
 XOR2_X2 \V2/V2/V4/V2/HA1/_1_  (.A(\V2/V2/V4/V2/w2 ),
    .B(\V2/V2/V4/V2/w1 ),
    .Z(\V2/V2/V4/v2 [1]));
 AND2_X1 \V2/V2/V4/V2/HA2/_0_  (.A1(\V2/V2/V4/V2/w4 ),
    .A2(\V2/V2/V4/V2/w3 ),
    .ZN(\V2/V2/V4/v2 [3]));
 XOR2_X2 \V2/V2/V4/V2/HA2/_1_  (.A(\V2/V2/V4/V2/w4 ),
    .B(\V2/V2/V4/V2/w3 ),
    .Z(\V2/V2/V4/v2 [2]));
 AND2_X1 \V2/V2/V4/V2/_0_  (.A1(A[30]),
    .A2(B[4]),
    .ZN(\V2/V2/V4/v2 [0]));
 AND2_X1 \V2/V2/V4/V2/_1_  (.A1(A[30]),
    .A2(B[5]),
    .ZN(\V2/V2/V4/V2/w1 ));
 AND2_X1 \V2/V2/V4/V2/_2_  (.A1(B[4]),
    .A2(A[31]),
    .ZN(\V2/V2/V4/V2/w2 ));
 AND2_X1 \V2/V2/V4/V2/_3_  (.A1(B[5]),
    .A2(A[31]),
    .ZN(\V2/V2/V4/V2/w3 ));
 AND2_X1 \V2/V2/V4/V3/HA1/_0_  (.A1(\V2/V2/V4/V3/w2 ),
    .A2(\V2/V2/V4/V3/w1 ),
    .ZN(\V2/V2/V4/V3/w4 ));
 XOR2_X2 \V2/V2/V4/V3/HA1/_1_  (.A(\V2/V2/V4/V3/w2 ),
    .B(\V2/V2/V4/V3/w1 ),
    .Z(\V2/V2/V4/v3 [1]));
 AND2_X1 \V2/V2/V4/V3/HA2/_0_  (.A1(\V2/V2/V4/V3/w4 ),
    .A2(\V2/V2/V4/V3/w3 ),
    .ZN(\V2/V2/V4/v3 [3]));
 XOR2_X2 \V2/V2/V4/V3/HA2/_1_  (.A(\V2/V2/V4/V3/w4 ),
    .B(\V2/V2/V4/V3/w3 ),
    .Z(\V2/V2/V4/v3 [2]));
 AND2_X1 \V2/V2/V4/V3/_0_  (.A1(A[28]),
    .A2(B[6]),
    .ZN(\V2/V2/V4/v3 [0]));
 AND2_X1 \V2/V2/V4/V3/_1_  (.A1(A[28]),
    .A2(B[7]),
    .ZN(\V2/V2/V4/V3/w1 ));
 AND2_X1 \V2/V2/V4/V3/_2_  (.A1(B[6]),
    .A2(A[29]),
    .ZN(\V2/V2/V4/V3/w2 ));
 AND2_X1 \V2/V2/V4/V3/_3_  (.A1(B[7]),
    .A2(A[29]),
    .ZN(\V2/V2/V4/V3/w3 ));
 AND2_X1 \V2/V2/V4/V4/HA1/_0_  (.A1(\V2/V2/V4/V4/w2 ),
    .A2(\V2/V2/V4/V4/w1 ),
    .ZN(\V2/V2/V4/V4/w4 ));
 XOR2_X2 \V2/V2/V4/V4/HA1/_1_  (.A(\V2/V2/V4/V4/w2 ),
    .B(\V2/V2/V4/V4/w1 ),
    .Z(\V2/V2/V4/v4 [1]));
 AND2_X1 \V2/V2/V4/V4/HA2/_0_  (.A1(\V2/V2/V4/V4/w4 ),
    .A2(\V2/V2/V4/V4/w3 ),
    .ZN(\V2/V2/V4/v4 [3]));
 XOR2_X2 \V2/V2/V4/V4/HA2/_1_  (.A(\V2/V2/V4/V4/w4 ),
    .B(\V2/V2/V4/V4/w3 ),
    .Z(\V2/V2/V4/v4 [2]));
 AND2_X1 \V2/V2/V4/V4/_0_  (.A1(A[30]),
    .A2(B[6]),
    .ZN(\V2/V2/V4/v4 [0]));
 AND2_X1 \V2/V2/V4/V4/_1_  (.A1(A[30]),
    .A2(B[7]),
    .ZN(\V2/V2/V4/V4/w1 ));
 AND2_X1 \V2/V2/V4/V4/_2_  (.A1(B[6]),
    .A2(A[31]),
    .ZN(\V2/V2/V4/V4/w2 ));
 AND2_X1 \V2/V2/V4/V4/_3_  (.A1(B[7]),
    .A2(A[31]),
    .ZN(\V2/V2/V4/V4/w3 ));
 OR2_X1 \V2/V2/V4/_0_  (.A1(\V2/V2/V4/c1 ),
    .A2(\V2/V2/V4/c2 ),
    .ZN(\V2/V2/V4/c3 ));
 OR2_X1 \V2/V2/_0_  (.A1(\V2/V2/c1 ),
    .A2(\V2/V2/c2 ),
    .ZN(\V2/V2/c3 ));
 AND2_X1 \V2/V3/A1/A1/M1/M1/_0_  (.A1(\V2/V3/v2 [0]),
    .A2(\V2/V3/v3 [0]),
    .ZN(\V2/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M1/M1/_1_  (.A(\V2/V3/v2 [0]),
    .B(\V2/V3/v3 [0]),
    .Z(\V2/V3/A1/A1/M1/s1 ));
 AND2_X1 \V2/V3/A1/A1/M1/M2/_0_  (.A1(\V2/V3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M1/M2/_1_  (.A(\V2/V3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/s1 [0]));
 OR2_X1 \V2/V3/A1/A1/M1/_0_  (.A1(\V2/V3/A1/A1/M1/c1 ),
    .A2(\V2/V3/A1/A1/M1/c2 ),
    .ZN(\V2/V3/A1/A1/c1 ));
 AND2_X1 \V2/V3/A1/A1/M2/M1/_0_  (.A1(\V2/V3/v2 [1]),
    .A2(\V2/V3/v3 [1]),
    .ZN(\V2/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M2/M1/_1_  (.A(\V2/V3/v2 [1]),
    .B(\V2/V3/v3 [1]),
    .Z(\V2/V3/A1/A1/M2/s1 ));
 AND2_X1 \V2/V3/A1/A1/M2/M2/_0_  (.A1(\V2/V3/A1/A1/M2/s1 ),
    .A2(\V2/V3/A1/A1/c1 ),
    .ZN(\V2/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M2/M2/_1_  (.A(\V2/V3/A1/A1/M2/s1 ),
    .B(\V2/V3/A1/A1/c1 ),
    .Z(\V2/V3/s1 [1]));
 OR2_X1 \V2/V3/A1/A1/M2/_0_  (.A1(\V2/V3/A1/A1/M2/c1 ),
    .A2(\V2/V3/A1/A1/M2/c2 ),
    .ZN(\V2/V3/A1/A1/c2 ));
 AND2_X1 \V2/V3/A1/A1/M3/M1/_0_  (.A1(\V2/V3/v2 [2]),
    .A2(\V2/V3/v3 [2]),
    .ZN(\V2/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M3/M1/_1_  (.A(\V2/V3/v2 [2]),
    .B(\V2/V3/v3 [2]),
    .Z(\V2/V3/A1/A1/M3/s1 ));
 AND2_X1 \V2/V3/A1/A1/M3/M2/_0_  (.A1(\V2/V3/A1/A1/M3/s1 ),
    .A2(\V2/V3/A1/A1/c2 ),
    .ZN(\V2/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M3/M2/_1_  (.A(\V2/V3/A1/A1/M3/s1 ),
    .B(\V2/V3/A1/A1/c2 ),
    .Z(\V2/V3/s1 [2]));
 OR2_X1 \V2/V3/A1/A1/M3/_0_  (.A1(\V2/V3/A1/A1/M3/c1 ),
    .A2(\V2/V3/A1/A1/M3/c2 ),
    .ZN(\V2/V3/A1/A1/c3 ));
 AND2_X1 \V2/V3/A1/A1/M4/M1/_0_  (.A1(\V2/V3/v2 [3]),
    .A2(\V2/V3/v3 [3]),
    .ZN(\V2/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M4/M1/_1_  (.A(\V2/V3/v2 [3]),
    .B(\V2/V3/v3 [3]),
    .Z(\V2/V3/A1/A1/M4/s1 ));
 AND2_X1 \V2/V3/A1/A1/M4/M2/_0_  (.A1(\V2/V3/A1/A1/M4/s1 ),
    .A2(\V2/V3/A1/A1/c3 ),
    .ZN(\V2/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M4/M2/_1_  (.A(\V2/V3/A1/A1/M4/s1 ),
    .B(\V2/V3/A1/A1/c3 ),
    .Z(\V2/V3/s1 [3]));
 OR2_X1 \V2/V3/A1/A1/M4/_0_  (.A1(\V2/V3/A1/A1/M4/c1 ),
    .A2(\V2/V3/A1/A1/M4/c2 ),
    .ZN(\V2/V3/A1/c1 ));
 AND2_X1 \V2/V3/A1/A2/M1/M1/_0_  (.A1(\V2/V3/v2 [4]),
    .A2(\V2/V3/v3 [4]),
    .ZN(\V2/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M1/M1/_1_  (.A(\V2/V3/v2 [4]),
    .B(\V2/V3/v3 [4]),
    .Z(\V2/V3/A1/A2/M1/s1 ));
 AND2_X1 \V2/V3/A1/A2/M1/M2/_0_  (.A1(\V2/V3/A1/A2/M1/s1 ),
    .A2(\V2/V3/A1/c1 ),
    .ZN(\V2/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M1/M2/_1_  (.A(\V2/V3/A1/A2/M1/s1 ),
    .B(\V2/V3/A1/c1 ),
    .Z(\V2/V3/s1 [4]));
 OR2_X1 \V2/V3/A1/A2/M1/_0_  (.A1(\V2/V3/A1/A2/M1/c1 ),
    .A2(\V2/V3/A1/A2/M1/c2 ),
    .ZN(\V2/V3/A1/A2/c1 ));
 AND2_X1 \V2/V3/A1/A2/M2/M1/_0_  (.A1(\V2/V3/v2 [5]),
    .A2(\V2/V3/v3 [5]),
    .ZN(\V2/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M2/M1/_1_  (.A(\V2/V3/v2 [5]),
    .B(\V2/V3/v3 [5]),
    .Z(\V2/V3/A1/A2/M2/s1 ));
 AND2_X1 \V2/V3/A1/A2/M2/M2/_0_  (.A1(\V2/V3/A1/A2/M2/s1 ),
    .A2(\V2/V3/A1/A2/c1 ),
    .ZN(\V2/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M2/M2/_1_  (.A(\V2/V3/A1/A2/M2/s1 ),
    .B(\V2/V3/A1/A2/c1 ),
    .Z(\V2/V3/s1 [5]));
 OR2_X1 \V2/V3/A1/A2/M2/_0_  (.A1(\V2/V3/A1/A2/M2/c1 ),
    .A2(\V2/V3/A1/A2/M2/c2 ),
    .ZN(\V2/V3/A1/A2/c2 ));
 AND2_X1 \V2/V3/A1/A2/M3/M1/_0_  (.A1(\V2/V3/v2 [6]),
    .A2(\V2/V3/v3 [6]),
    .ZN(\V2/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M3/M1/_1_  (.A(\V2/V3/v2 [6]),
    .B(\V2/V3/v3 [6]),
    .Z(\V2/V3/A1/A2/M3/s1 ));
 AND2_X1 \V2/V3/A1/A2/M3/M2/_0_  (.A1(\V2/V3/A1/A2/M3/s1 ),
    .A2(\V2/V3/A1/A2/c2 ),
    .ZN(\V2/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M3/M2/_1_  (.A(\V2/V3/A1/A2/M3/s1 ),
    .B(\V2/V3/A1/A2/c2 ),
    .Z(\V2/V3/s1 [6]));
 OR2_X1 \V2/V3/A1/A2/M3/_0_  (.A1(\V2/V3/A1/A2/M3/c1 ),
    .A2(\V2/V3/A1/A2/M3/c2 ),
    .ZN(\V2/V3/A1/A2/c3 ));
 AND2_X1 \V2/V3/A1/A2/M4/M1/_0_  (.A1(\V2/V3/v2 [7]),
    .A2(\V2/V3/v3 [7]),
    .ZN(\V2/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M4/M1/_1_  (.A(\V2/V3/v2 [7]),
    .B(\V2/V3/v3 [7]),
    .Z(\V2/V3/A1/A2/M4/s1 ));
 AND2_X1 \V2/V3/A1/A2/M4/M2/_0_  (.A1(\V2/V3/A1/A2/M4/s1 ),
    .A2(\V2/V3/A1/A2/c3 ),
    .ZN(\V2/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M4/M2/_1_  (.A(\V2/V3/A1/A2/M4/s1 ),
    .B(\V2/V3/A1/A2/c3 ),
    .Z(\V2/V3/s1 [7]));
 OR2_X1 \V2/V3/A1/A2/M4/_0_  (.A1(\V2/V3/A1/A2/M4/c1 ),
    .A2(\V2/V3/A1/A2/M4/c2 ),
    .ZN(\V2/V3/c1 ));
 AND2_X1 \V2/V3/A2/A1/M1/M1/_0_  (.A1(\V2/V3/s1 [0]),
    .A2(\V2/V3/v1 [4]),
    .ZN(\V2/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M1/M1/_1_  (.A(\V2/V3/s1 [0]),
    .B(\V2/V3/v1 [4]),
    .Z(\V2/V3/A2/A1/M1/s1 ));
 AND2_X1 \V2/V3/A2/A1/M1/M2/_0_  (.A1(\V2/V3/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M1/M2/_1_  (.A(\V2/V3/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v3 [4]));
 OR2_X1 \V2/V3/A2/A1/M1/_0_  (.A1(\V2/V3/A2/A1/M1/c1 ),
    .A2(\V2/V3/A2/A1/M1/c2 ),
    .ZN(\V2/V3/A2/A1/c1 ));
 AND2_X1 \V2/V3/A2/A1/M2/M1/_0_  (.A1(\V2/V3/s1 [1]),
    .A2(\V2/V3/v1 [5]),
    .ZN(\V2/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M2/M1/_1_  (.A(\V2/V3/s1 [1]),
    .B(\V2/V3/v1 [5]),
    .Z(\V2/V3/A2/A1/M2/s1 ));
 AND2_X1 \V2/V3/A2/A1/M2/M2/_0_  (.A1(\V2/V3/A2/A1/M2/s1 ),
    .A2(\V2/V3/A2/A1/c1 ),
    .ZN(\V2/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M2/M2/_1_  (.A(\V2/V3/A2/A1/M2/s1 ),
    .B(\V2/V3/A2/A1/c1 ),
    .Z(\V2/v3 [5]));
 OR2_X1 \V2/V3/A2/A1/M2/_0_  (.A1(\V2/V3/A2/A1/M2/c1 ),
    .A2(\V2/V3/A2/A1/M2/c2 ),
    .ZN(\V2/V3/A2/A1/c2 ));
 AND2_X1 \V2/V3/A2/A1/M3/M1/_0_  (.A1(\V2/V3/s1 [2]),
    .A2(\V2/V3/v1 [6]),
    .ZN(\V2/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M3/M1/_1_  (.A(\V2/V3/s1 [2]),
    .B(\V2/V3/v1 [6]),
    .Z(\V2/V3/A2/A1/M3/s1 ));
 AND2_X1 \V2/V3/A2/A1/M3/M2/_0_  (.A1(\V2/V3/A2/A1/M3/s1 ),
    .A2(\V2/V3/A2/A1/c2 ),
    .ZN(\V2/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M3/M2/_1_  (.A(\V2/V3/A2/A1/M3/s1 ),
    .B(\V2/V3/A2/A1/c2 ),
    .Z(\V2/v3 [6]));
 OR2_X1 \V2/V3/A2/A1/M3/_0_  (.A1(\V2/V3/A2/A1/M3/c1 ),
    .A2(\V2/V3/A2/A1/M3/c2 ),
    .ZN(\V2/V3/A2/A1/c3 ));
 AND2_X1 \V2/V3/A2/A1/M4/M1/_0_  (.A1(\V2/V3/s1 [3]),
    .A2(\V2/V3/v1 [7]),
    .ZN(\V2/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M4/M1/_1_  (.A(\V2/V3/s1 [3]),
    .B(\V2/V3/v1 [7]),
    .Z(\V2/V3/A2/A1/M4/s1 ));
 AND2_X1 \V2/V3/A2/A1/M4/M2/_0_  (.A1(\V2/V3/A2/A1/M4/s1 ),
    .A2(\V2/V3/A2/A1/c3 ),
    .ZN(\V2/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M4/M2/_1_  (.A(\V2/V3/A2/A1/M4/s1 ),
    .B(\V2/V3/A2/A1/c3 ),
    .Z(\V2/v3 [7]));
 OR2_X1 \V2/V3/A2/A1/M4/_0_  (.A1(\V2/V3/A2/A1/M4/c1 ),
    .A2(\V2/V3/A2/A1/M4/c2 ),
    .ZN(\V2/V3/A2/c1 ));
 AND2_X1 \V2/V3/A2/A2/M1/M1/_0_  (.A1(\V2/V3/s1 [4]),
    .A2(ground),
    .ZN(\V2/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M1/M1/_1_  (.A(\V2/V3/s1 [4]),
    .B(ground),
    .Z(\V2/V3/A2/A2/M1/s1 ));
 AND2_X1 \V2/V3/A2/A2/M1/M2/_0_  (.A1(\V2/V3/A2/A2/M1/s1 ),
    .A2(\V2/V3/A2/c1 ),
    .ZN(\V2/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M1/M2/_1_  (.A(\V2/V3/A2/A2/M1/s1 ),
    .B(\V2/V3/A2/c1 ),
    .Z(\V2/V3/s2 [4]));
 OR2_X1 \V2/V3/A2/A2/M1/_0_  (.A1(\V2/V3/A2/A2/M1/c1 ),
    .A2(\V2/V3/A2/A2/M1/c2 ),
    .ZN(\V2/V3/A2/A2/c1 ));
 AND2_X1 \V2/V3/A2/A2/M2/M1/_0_  (.A1(\V2/V3/s1 [5]),
    .A2(ground),
    .ZN(\V2/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M2/M1/_1_  (.A(\V2/V3/s1 [5]),
    .B(ground),
    .Z(\V2/V3/A2/A2/M2/s1 ));
 AND2_X1 \V2/V3/A2/A2/M2/M2/_0_  (.A1(\V2/V3/A2/A2/M2/s1 ),
    .A2(\V2/V3/A2/A2/c1 ),
    .ZN(\V2/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M2/M2/_1_  (.A(\V2/V3/A2/A2/M2/s1 ),
    .B(\V2/V3/A2/A2/c1 ),
    .Z(\V2/V3/s2 [5]));
 OR2_X1 \V2/V3/A2/A2/M2/_0_  (.A1(\V2/V3/A2/A2/M2/c1 ),
    .A2(\V2/V3/A2/A2/M2/c2 ),
    .ZN(\V2/V3/A2/A2/c2 ));
 AND2_X1 \V2/V3/A2/A2/M3/M1/_0_  (.A1(\V2/V3/s1 [6]),
    .A2(ground),
    .ZN(\V2/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M3/M1/_1_  (.A(\V2/V3/s1 [6]),
    .B(ground),
    .Z(\V2/V3/A2/A2/M3/s1 ));
 AND2_X1 \V2/V3/A2/A2/M3/M2/_0_  (.A1(\V2/V3/A2/A2/M3/s1 ),
    .A2(\V2/V3/A2/A2/c2 ),
    .ZN(\V2/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M3/M2/_1_  (.A(\V2/V3/A2/A2/M3/s1 ),
    .B(\V2/V3/A2/A2/c2 ),
    .Z(\V2/V3/s2 [6]));
 OR2_X1 \V2/V3/A2/A2/M3/_0_  (.A1(\V2/V3/A2/A2/M3/c1 ),
    .A2(\V2/V3/A2/A2/M3/c2 ),
    .ZN(\V2/V3/A2/A2/c3 ));
 AND2_X1 \V2/V3/A2/A2/M4/M1/_0_  (.A1(\V2/V3/s1 [7]),
    .A2(ground),
    .ZN(\V2/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M4/M1/_1_  (.A(\V2/V3/s1 [7]),
    .B(ground),
    .Z(\V2/V3/A2/A2/M4/s1 ));
 AND2_X1 \V2/V3/A2/A2/M4/M2/_0_  (.A1(\V2/V3/A2/A2/M4/s1 ),
    .A2(\V2/V3/A2/A2/c3 ),
    .ZN(\V2/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M4/M2/_1_  (.A(\V2/V3/A2/A2/M4/s1 ),
    .B(\V2/V3/A2/A2/c3 ),
    .Z(\V2/V3/s2 [7]));
 OR2_X1 \V2/V3/A2/A2/M4/_0_  (.A1(\V2/V3/A2/A2/M4/c1 ),
    .A2(\V2/V3/A2/A2/M4/c2 ),
    .ZN(\V2/V3/c2 ));
 AND2_X1 \V2/V3/A3/A1/M1/M1/_0_  (.A1(\V2/V3/v4 [0]),
    .A2(\V2/V3/s2 [4]),
    .ZN(\V2/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M1/M1/_1_  (.A(\V2/V3/v4 [0]),
    .B(\V2/V3/s2 [4]),
    .Z(\V2/V3/A3/A1/M1/s1 ));
 AND2_X1 \V2/V3/A3/A1/M1/M2/_0_  (.A1(\V2/V3/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M1/M2/_1_  (.A(\V2/V3/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v3 [8]));
 OR2_X1 \V2/V3/A3/A1/M1/_0_  (.A1(\V2/V3/A3/A1/M1/c1 ),
    .A2(\V2/V3/A3/A1/M1/c2 ),
    .ZN(\V2/V3/A3/A1/c1 ));
 AND2_X1 \V2/V3/A3/A1/M2/M1/_0_  (.A1(\V2/V3/v4 [1]),
    .A2(\V2/V3/s2 [5]),
    .ZN(\V2/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M2/M1/_1_  (.A(\V2/V3/v4 [1]),
    .B(\V2/V3/s2 [5]),
    .Z(\V2/V3/A3/A1/M2/s1 ));
 AND2_X1 \V2/V3/A3/A1/M2/M2/_0_  (.A1(\V2/V3/A3/A1/M2/s1 ),
    .A2(\V2/V3/A3/A1/c1 ),
    .ZN(\V2/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M2/M2/_1_  (.A(\V2/V3/A3/A1/M2/s1 ),
    .B(\V2/V3/A3/A1/c1 ),
    .Z(\V2/v3 [9]));
 OR2_X1 \V2/V3/A3/A1/M2/_0_  (.A1(\V2/V3/A3/A1/M2/c1 ),
    .A2(\V2/V3/A3/A1/M2/c2 ),
    .ZN(\V2/V3/A3/A1/c2 ));
 AND2_X1 \V2/V3/A3/A1/M3/M1/_0_  (.A1(\V2/V3/v4 [2]),
    .A2(\V2/V3/s2 [6]),
    .ZN(\V2/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M3/M1/_1_  (.A(\V2/V3/v4 [2]),
    .B(\V2/V3/s2 [6]),
    .Z(\V2/V3/A3/A1/M3/s1 ));
 AND2_X1 \V2/V3/A3/A1/M3/M2/_0_  (.A1(\V2/V3/A3/A1/M3/s1 ),
    .A2(\V2/V3/A3/A1/c2 ),
    .ZN(\V2/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M3/M2/_1_  (.A(\V2/V3/A3/A1/M3/s1 ),
    .B(\V2/V3/A3/A1/c2 ),
    .Z(\V2/v3 [10]));
 OR2_X1 \V2/V3/A3/A1/M3/_0_  (.A1(\V2/V3/A3/A1/M3/c1 ),
    .A2(\V2/V3/A3/A1/M3/c2 ),
    .ZN(\V2/V3/A3/A1/c3 ));
 AND2_X1 \V2/V3/A3/A1/M4/M1/_0_  (.A1(\V2/V3/v4 [3]),
    .A2(\V2/V3/s2 [7]),
    .ZN(\V2/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M4/M1/_1_  (.A(\V2/V3/v4 [3]),
    .B(\V2/V3/s2 [7]),
    .Z(\V2/V3/A3/A1/M4/s1 ));
 AND2_X1 \V2/V3/A3/A1/M4/M2/_0_  (.A1(\V2/V3/A3/A1/M4/s1 ),
    .A2(\V2/V3/A3/A1/c3 ),
    .ZN(\V2/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M4/M2/_1_  (.A(\V2/V3/A3/A1/M4/s1 ),
    .B(\V2/V3/A3/A1/c3 ),
    .Z(\V2/v3 [11]));
 OR2_X1 \V2/V3/A3/A1/M4/_0_  (.A1(\V2/V3/A3/A1/M4/c1 ),
    .A2(\V2/V3/A3/A1/M4/c2 ),
    .ZN(\V2/V3/A3/c1 ));
 AND2_X1 \V2/V3/A3/A2/M1/M1/_0_  (.A1(\V2/V3/v4 [4]),
    .A2(\V2/V3/c3 ),
    .ZN(\V2/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M1/M1/_1_  (.A(\V2/V3/v4 [4]),
    .B(\V2/V3/c3 ),
    .Z(\V2/V3/A3/A2/M1/s1 ));
 AND2_X1 \V2/V3/A3/A2/M1/M2/_0_  (.A1(\V2/V3/A3/A2/M1/s1 ),
    .A2(\V2/V3/A3/c1 ),
    .ZN(\V2/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M1/M2/_1_  (.A(\V2/V3/A3/A2/M1/s1 ),
    .B(\V2/V3/A3/c1 ),
    .Z(\V2/v3 [12]));
 OR2_X1 \V2/V3/A3/A2/M1/_0_  (.A1(\V2/V3/A3/A2/M1/c1 ),
    .A2(\V2/V3/A3/A2/M1/c2 ),
    .ZN(\V2/V3/A3/A2/c1 ));
 AND2_X1 \V2/V3/A3/A2/M2/M1/_0_  (.A1(\V2/V3/v4 [5]),
    .A2(ground),
    .ZN(\V2/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M2/M1/_1_  (.A(\V2/V3/v4 [5]),
    .B(ground),
    .Z(\V2/V3/A3/A2/M2/s1 ));
 AND2_X1 \V2/V3/A3/A2/M2/M2/_0_  (.A1(\V2/V3/A3/A2/M2/s1 ),
    .A2(\V2/V3/A3/A2/c1 ),
    .ZN(\V2/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M2/M2/_1_  (.A(\V2/V3/A3/A2/M2/s1 ),
    .B(\V2/V3/A3/A2/c1 ),
    .Z(\V2/v3 [13]));
 OR2_X1 \V2/V3/A3/A2/M2/_0_  (.A1(\V2/V3/A3/A2/M2/c1 ),
    .A2(\V2/V3/A3/A2/M2/c2 ),
    .ZN(\V2/V3/A3/A2/c2 ));
 AND2_X1 \V2/V3/A3/A2/M3/M1/_0_  (.A1(\V2/V3/v4 [6]),
    .A2(ground),
    .ZN(\V2/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M3/M1/_1_  (.A(\V2/V3/v4 [6]),
    .B(ground),
    .Z(\V2/V3/A3/A2/M3/s1 ));
 AND2_X1 \V2/V3/A3/A2/M3/M2/_0_  (.A1(\V2/V3/A3/A2/M3/s1 ),
    .A2(\V2/V3/A3/A2/c2 ),
    .ZN(\V2/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M3/M2/_1_  (.A(\V2/V3/A3/A2/M3/s1 ),
    .B(\V2/V3/A3/A2/c2 ),
    .Z(\V2/v3 [14]));
 OR2_X1 \V2/V3/A3/A2/M3/_0_  (.A1(\V2/V3/A3/A2/M3/c1 ),
    .A2(\V2/V3/A3/A2/M3/c2 ),
    .ZN(\V2/V3/A3/A2/c3 ));
 AND2_X1 \V2/V3/A3/A2/M4/M1/_0_  (.A1(\V2/V3/v4 [7]),
    .A2(ground),
    .ZN(\V2/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M4/M1/_1_  (.A(\V2/V3/v4 [7]),
    .B(ground),
    .Z(\V2/V3/A3/A2/M4/s1 ));
 AND2_X1 \V2/V3/A3/A2/M4/M2/_0_  (.A1(\V2/V3/A3/A2/M4/s1 ),
    .A2(\V2/V3/A3/A2/c3 ),
    .ZN(\V2/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M4/M2/_1_  (.A(\V2/V3/A3/A2/M4/s1 ),
    .B(\V2/V3/A3/A2/c3 ),
    .Z(\V2/v3 [15]));
 OR2_X1 \V2/V3/A3/A2/M4/_0_  (.A1(\V2/V3/A3/A2/M4/c1 ),
    .A2(\V2/V3/A3/A2/M4/c2 ),
    .ZN(\V2/V3/overflow ));
 AND2_X1 \V2/V3/V1/A1/M1/M1/_0_  (.A1(\V2/V3/V1/v2 [0]),
    .A2(\V2/V3/V1/v3 [0]),
    .ZN(\V2/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M1/M1/_1_  (.A(\V2/V3/V1/v2 [0]),
    .B(\V2/V3/V1/v3 [0]),
    .Z(\V2/V3/V1/A1/M1/s1 ));
 AND2_X1 \V2/V3/V1/A1/M1/M2/_0_  (.A1(\V2/V3/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M1/M2/_1_  (.A(\V2/V3/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/V1/s1 [0]));
 OR2_X1 \V2/V3/V1/A1/M1/_0_  (.A1(\V2/V3/V1/A1/M1/c1 ),
    .A2(\V2/V3/V1/A1/M1/c2 ),
    .ZN(\V2/V3/V1/A1/c1 ));
 AND2_X1 \V2/V3/V1/A1/M2/M1/_0_  (.A1(\V2/V3/V1/v2 [1]),
    .A2(\V2/V3/V1/v3 [1]),
    .ZN(\V2/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M2/M1/_1_  (.A(\V2/V3/V1/v2 [1]),
    .B(\V2/V3/V1/v3 [1]),
    .Z(\V2/V3/V1/A1/M2/s1 ));
 AND2_X1 \V2/V3/V1/A1/M2/M2/_0_  (.A1(\V2/V3/V1/A1/M2/s1 ),
    .A2(\V2/V3/V1/A1/c1 ),
    .ZN(\V2/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M2/M2/_1_  (.A(\V2/V3/V1/A1/M2/s1 ),
    .B(\V2/V3/V1/A1/c1 ),
    .Z(\V2/V3/V1/s1 [1]));
 OR2_X1 \V2/V3/V1/A1/M2/_0_  (.A1(\V2/V3/V1/A1/M2/c1 ),
    .A2(\V2/V3/V1/A1/M2/c2 ),
    .ZN(\V2/V3/V1/A1/c2 ));
 AND2_X1 \V2/V3/V1/A1/M3/M1/_0_  (.A1(\V2/V3/V1/v2 [2]),
    .A2(\V2/V3/V1/v3 [2]),
    .ZN(\V2/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M3/M1/_1_  (.A(\V2/V3/V1/v2 [2]),
    .B(\V2/V3/V1/v3 [2]),
    .Z(\V2/V3/V1/A1/M3/s1 ));
 AND2_X1 \V2/V3/V1/A1/M3/M2/_0_  (.A1(\V2/V3/V1/A1/M3/s1 ),
    .A2(\V2/V3/V1/A1/c2 ),
    .ZN(\V2/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M3/M2/_1_  (.A(\V2/V3/V1/A1/M3/s1 ),
    .B(\V2/V3/V1/A1/c2 ),
    .Z(\V2/V3/V1/s1 [2]));
 OR2_X1 \V2/V3/V1/A1/M3/_0_  (.A1(\V2/V3/V1/A1/M3/c1 ),
    .A2(\V2/V3/V1/A1/M3/c2 ),
    .ZN(\V2/V3/V1/A1/c3 ));
 AND2_X1 \V2/V3/V1/A1/M4/M1/_0_  (.A1(\V2/V3/V1/v2 [3]),
    .A2(\V2/V3/V1/v3 [3]),
    .ZN(\V2/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M4/M1/_1_  (.A(\V2/V3/V1/v2 [3]),
    .B(\V2/V3/V1/v3 [3]),
    .Z(\V2/V3/V1/A1/M4/s1 ));
 AND2_X1 \V2/V3/V1/A1/M4/M2/_0_  (.A1(\V2/V3/V1/A1/M4/s1 ),
    .A2(\V2/V3/V1/A1/c3 ),
    .ZN(\V2/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M4/M2/_1_  (.A(\V2/V3/V1/A1/M4/s1 ),
    .B(\V2/V3/V1/A1/c3 ),
    .Z(\V2/V3/V1/s1 [3]));
 OR2_X1 \V2/V3/V1/A1/M4/_0_  (.A1(\V2/V3/V1/A1/M4/c1 ),
    .A2(\V2/V3/V1/A1/M4/c2 ),
    .ZN(\V2/V3/V1/c1 ));
 AND2_X1 \V2/V3/V1/A2/M1/M1/_0_  (.A1(\V2/V3/V1/s1 [0]),
    .A2(\V2/V3/V1/v1 [2]),
    .ZN(\V2/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M1/M1/_1_  (.A(\V2/V3/V1/s1 [0]),
    .B(\V2/V3/V1/v1 [2]),
    .Z(\V2/V3/V1/A2/M1/s1 ));
 AND2_X1 \V2/V3/V1/A2/M1/M2/_0_  (.A1(\V2/V3/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M1/M2/_1_  (.A(\V2/V3/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/v3 [2]));
 OR2_X1 \V2/V3/V1/A2/M1/_0_  (.A1(\V2/V3/V1/A2/M1/c1 ),
    .A2(\V2/V3/V1/A2/M1/c2 ),
    .ZN(\V2/V3/V1/A2/c1 ));
 AND2_X1 \V2/V3/V1/A2/M2/M1/_0_  (.A1(\V2/V3/V1/s1 [1]),
    .A2(\V2/V3/V1/v1 [3]),
    .ZN(\V2/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M2/M1/_1_  (.A(\V2/V3/V1/s1 [1]),
    .B(\V2/V3/V1/v1 [3]),
    .Z(\V2/V3/V1/A2/M2/s1 ));
 AND2_X1 \V2/V3/V1/A2/M2/M2/_0_  (.A1(\V2/V3/V1/A2/M2/s1 ),
    .A2(\V2/V3/V1/A2/c1 ),
    .ZN(\V2/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M2/M2/_1_  (.A(\V2/V3/V1/A2/M2/s1 ),
    .B(\V2/V3/V1/A2/c1 ),
    .Z(\V2/v3 [3]));
 OR2_X1 \V2/V3/V1/A2/M2/_0_  (.A1(\V2/V3/V1/A2/M2/c1 ),
    .A2(\V2/V3/V1/A2/M2/c2 ),
    .ZN(\V2/V3/V1/A2/c2 ));
 AND2_X1 \V2/V3/V1/A2/M3/M1/_0_  (.A1(\V2/V3/V1/s1 [2]),
    .A2(ground),
    .ZN(\V2/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M3/M1/_1_  (.A(\V2/V3/V1/s1 [2]),
    .B(ground),
    .Z(\V2/V3/V1/A2/M3/s1 ));
 AND2_X1 \V2/V3/V1/A2/M3/M2/_0_  (.A1(\V2/V3/V1/A2/M3/s1 ),
    .A2(\V2/V3/V1/A2/c2 ),
    .ZN(\V2/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M3/M2/_1_  (.A(\V2/V3/V1/A2/M3/s1 ),
    .B(\V2/V3/V1/A2/c2 ),
    .Z(\V2/V3/V1/s2 [2]));
 OR2_X1 \V2/V3/V1/A2/M3/_0_  (.A1(\V2/V3/V1/A2/M3/c1 ),
    .A2(\V2/V3/V1/A2/M3/c2 ),
    .ZN(\V2/V3/V1/A2/c3 ));
 AND2_X1 \V2/V3/V1/A2/M4/M1/_0_  (.A1(\V2/V3/V1/s1 [3]),
    .A2(ground),
    .ZN(\V2/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M4/M1/_1_  (.A(\V2/V3/V1/s1 [3]),
    .B(ground),
    .Z(\V2/V3/V1/A2/M4/s1 ));
 AND2_X1 \V2/V3/V1/A2/M4/M2/_0_  (.A1(\V2/V3/V1/A2/M4/s1 ),
    .A2(\V2/V3/V1/A2/c3 ),
    .ZN(\V2/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M4/M2/_1_  (.A(\V2/V3/V1/A2/M4/s1 ),
    .B(\V2/V3/V1/A2/c3 ),
    .Z(\V2/V3/V1/s2 [3]));
 OR2_X1 \V2/V3/V1/A2/M4/_0_  (.A1(\V2/V3/V1/A2/M4/c1 ),
    .A2(\V2/V3/V1/A2/M4/c2 ),
    .ZN(\V2/V3/V1/c2 ));
 AND2_X1 \V2/V3/V1/A3/M1/M1/_0_  (.A1(\V2/V3/V1/v4 [0]),
    .A2(\V2/V3/V1/s2 [2]),
    .ZN(\V2/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M1/M1/_1_  (.A(\V2/V3/V1/v4 [0]),
    .B(\V2/V3/V1/s2 [2]),
    .Z(\V2/V3/V1/A3/M1/s1 ));
 AND2_X1 \V2/V3/V1/A3/M1/M2/_0_  (.A1(\V2/V3/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M1/M2/_1_  (.A(\V2/V3/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v1 [4]));
 OR2_X1 \V2/V3/V1/A3/M1/_0_  (.A1(\V2/V3/V1/A3/M1/c1 ),
    .A2(\V2/V3/V1/A3/M1/c2 ),
    .ZN(\V2/V3/V1/A3/c1 ));
 AND2_X1 \V2/V3/V1/A3/M2/M1/_0_  (.A1(\V2/V3/V1/v4 [1]),
    .A2(\V2/V3/V1/s2 [3]),
    .ZN(\V2/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M2/M1/_1_  (.A(\V2/V3/V1/v4 [1]),
    .B(\V2/V3/V1/s2 [3]),
    .Z(\V2/V3/V1/A3/M2/s1 ));
 AND2_X1 \V2/V3/V1/A3/M2/M2/_0_  (.A1(\V2/V3/V1/A3/M2/s1 ),
    .A2(\V2/V3/V1/A3/c1 ),
    .ZN(\V2/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M2/M2/_1_  (.A(\V2/V3/V1/A3/M2/s1 ),
    .B(\V2/V3/V1/A3/c1 ),
    .Z(\V2/V3/v1 [5]));
 OR2_X1 \V2/V3/V1/A3/M2/_0_  (.A1(\V2/V3/V1/A3/M2/c1 ),
    .A2(\V2/V3/V1/A3/M2/c2 ),
    .ZN(\V2/V3/V1/A3/c2 ));
 AND2_X1 \V2/V3/V1/A3/M3/M1/_0_  (.A1(\V2/V3/V1/v4 [2]),
    .A2(\V2/V3/V1/c3 ),
    .ZN(\V2/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M3/M1/_1_  (.A(\V2/V3/V1/v4 [2]),
    .B(\V2/V3/V1/c3 ),
    .Z(\V2/V3/V1/A3/M3/s1 ));
 AND2_X1 \V2/V3/V1/A3/M3/M2/_0_  (.A1(\V2/V3/V1/A3/M3/s1 ),
    .A2(\V2/V3/V1/A3/c2 ),
    .ZN(\V2/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M3/M2/_1_  (.A(\V2/V3/V1/A3/M3/s1 ),
    .B(\V2/V3/V1/A3/c2 ),
    .Z(\V2/V3/v1 [6]));
 OR2_X1 \V2/V3/V1/A3/M3/_0_  (.A1(\V2/V3/V1/A3/M3/c1 ),
    .A2(\V2/V3/V1/A3/M3/c2 ),
    .ZN(\V2/V3/V1/A3/c3 ));
 AND2_X1 \V2/V3/V1/A3/M4/M1/_0_  (.A1(\V2/V3/V1/v4 [3]),
    .A2(ground),
    .ZN(\V2/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M4/M1/_1_  (.A(\V2/V3/V1/v4 [3]),
    .B(ground),
    .Z(\V2/V3/V1/A3/M4/s1 ));
 AND2_X1 \V2/V3/V1/A3/M4/M2/_0_  (.A1(\V2/V3/V1/A3/M4/s1 ),
    .A2(\V2/V3/V1/A3/c3 ),
    .ZN(\V2/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M4/M2/_1_  (.A(\V2/V3/V1/A3/M4/s1 ),
    .B(\V2/V3/V1/A3/c3 ),
    .Z(\V2/V3/v1 [7]));
 OR2_X1 \V2/V3/V1/A3/M4/_0_  (.A1(\V2/V3/V1/A3/M4/c1 ),
    .A2(\V2/V3/V1/A3/M4/c2 ),
    .ZN(\V2/V3/V1/overflow ));
 AND2_X1 \V2/V3/V1/V1/HA1/_0_  (.A1(\V2/V3/V1/V1/w2 ),
    .A2(\V2/V3/V1/V1/w1 ),
    .ZN(\V2/V3/V1/V1/w4 ));
 XOR2_X2 \V2/V3/V1/V1/HA1/_1_  (.A(\V2/V3/V1/V1/w2 ),
    .B(\V2/V3/V1/V1/w1 ),
    .Z(\V2/v3 [1]));
 AND2_X1 \V2/V3/V1/V1/HA2/_0_  (.A1(\V2/V3/V1/V1/w4 ),
    .A2(\V2/V3/V1/V1/w3 ),
    .ZN(\V2/V3/V1/v1 [3]));
 XOR2_X2 \V2/V3/V1/V1/HA2/_1_  (.A(\V2/V3/V1/V1/w4 ),
    .B(\V2/V3/V1/V1/w3 ),
    .Z(\V2/V3/V1/v1 [2]));
 AND2_X1 \V2/V3/V1/V1/_0_  (.A1(A[16]),
    .A2(B[8]),
    .ZN(\V2/v3 [0]));
 AND2_X1 \V2/V3/V1/V1/_1_  (.A1(A[16]),
    .A2(B[9]),
    .ZN(\V2/V3/V1/V1/w1 ));
 AND2_X1 \V2/V3/V1/V1/_2_  (.A1(B[8]),
    .A2(A[17]),
    .ZN(\V2/V3/V1/V1/w2 ));
 AND2_X1 \V2/V3/V1/V1/_3_  (.A1(B[9]),
    .A2(A[17]),
    .ZN(\V2/V3/V1/V1/w3 ));
 AND2_X1 \V2/V3/V1/V2/HA1/_0_  (.A1(\V2/V3/V1/V2/w2 ),
    .A2(\V2/V3/V1/V2/w1 ),
    .ZN(\V2/V3/V1/V2/w4 ));
 XOR2_X2 \V2/V3/V1/V2/HA1/_1_  (.A(\V2/V3/V1/V2/w2 ),
    .B(\V2/V3/V1/V2/w1 ),
    .Z(\V2/V3/V1/v2 [1]));
 AND2_X1 \V2/V3/V1/V2/HA2/_0_  (.A1(\V2/V3/V1/V2/w4 ),
    .A2(\V2/V3/V1/V2/w3 ),
    .ZN(\V2/V3/V1/v2 [3]));
 XOR2_X2 \V2/V3/V1/V2/HA2/_1_  (.A(\V2/V3/V1/V2/w4 ),
    .B(\V2/V3/V1/V2/w3 ),
    .Z(\V2/V3/V1/v2 [2]));
 AND2_X1 \V2/V3/V1/V2/_0_  (.A1(A[18]),
    .A2(B[8]),
    .ZN(\V2/V3/V1/v2 [0]));
 AND2_X1 \V2/V3/V1/V2/_1_  (.A1(A[18]),
    .A2(B[9]),
    .ZN(\V2/V3/V1/V2/w1 ));
 AND2_X1 \V2/V3/V1/V2/_2_  (.A1(B[8]),
    .A2(A[19]),
    .ZN(\V2/V3/V1/V2/w2 ));
 AND2_X1 \V2/V3/V1/V2/_3_  (.A1(B[9]),
    .A2(A[19]),
    .ZN(\V2/V3/V1/V2/w3 ));
 AND2_X1 \V2/V3/V1/V3/HA1/_0_  (.A1(\V2/V3/V1/V3/w2 ),
    .A2(\V2/V3/V1/V3/w1 ),
    .ZN(\V2/V3/V1/V3/w4 ));
 XOR2_X2 \V2/V3/V1/V3/HA1/_1_  (.A(\V2/V3/V1/V3/w2 ),
    .B(\V2/V3/V1/V3/w1 ),
    .Z(\V2/V3/V1/v3 [1]));
 AND2_X1 \V2/V3/V1/V3/HA2/_0_  (.A1(\V2/V3/V1/V3/w4 ),
    .A2(\V2/V3/V1/V3/w3 ),
    .ZN(\V2/V3/V1/v3 [3]));
 XOR2_X2 \V2/V3/V1/V3/HA2/_1_  (.A(\V2/V3/V1/V3/w4 ),
    .B(\V2/V3/V1/V3/w3 ),
    .Z(\V2/V3/V1/v3 [2]));
 AND2_X1 \V2/V3/V1/V3/_0_  (.A1(A[16]),
    .A2(B[10]),
    .ZN(\V2/V3/V1/v3 [0]));
 AND2_X1 \V2/V3/V1/V3/_1_  (.A1(A[16]),
    .A2(B[11]),
    .ZN(\V2/V3/V1/V3/w1 ));
 AND2_X1 \V2/V3/V1/V3/_2_  (.A1(B[10]),
    .A2(A[17]),
    .ZN(\V2/V3/V1/V3/w2 ));
 AND2_X1 \V2/V3/V1/V3/_3_  (.A1(B[11]),
    .A2(A[17]),
    .ZN(\V2/V3/V1/V3/w3 ));
 AND2_X1 \V2/V3/V1/V4/HA1/_0_  (.A1(\V2/V3/V1/V4/w2 ),
    .A2(\V2/V3/V1/V4/w1 ),
    .ZN(\V2/V3/V1/V4/w4 ));
 XOR2_X2 \V2/V3/V1/V4/HA1/_1_  (.A(\V2/V3/V1/V4/w2 ),
    .B(\V2/V3/V1/V4/w1 ),
    .Z(\V2/V3/V1/v4 [1]));
 AND2_X1 \V2/V3/V1/V4/HA2/_0_  (.A1(\V2/V3/V1/V4/w4 ),
    .A2(\V2/V3/V1/V4/w3 ),
    .ZN(\V2/V3/V1/v4 [3]));
 XOR2_X2 \V2/V3/V1/V4/HA2/_1_  (.A(\V2/V3/V1/V4/w4 ),
    .B(\V2/V3/V1/V4/w3 ),
    .Z(\V2/V3/V1/v4 [2]));
 AND2_X1 \V2/V3/V1/V4/_0_  (.A1(A[18]),
    .A2(B[10]),
    .ZN(\V2/V3/V1/v4 [0]));
 AND2_X1 \V2/V3/V1/V4/_1_  (.A1(A[18]),
    .A2(B[11]),
    .ZN(\V2/V3/V1/V4/w1 ));
 AND2_X1 \V2/V3/V1/V4/_2_  (.A1(B[10]),
    .A2(A[19]),
    .ZN(\V2/V3/V1/V4/w2 ));
 AND2_X1 \V2/V3/V1/V4/_3_  (.A1(B[11]),
    .A2(A[19]),
    .ZN(\V2/V3/V1/V4/w3 ));
 OR2_X1 \V2/V3/V1/_0_  (.A1(\V2/V3/V1/c1 ),
    .A2(\V2/V3/V1/c2 ),
    .ZN(\V2/V3/V1/c3 ));
 AND2_X1 \V2/V3/V2/A1/M1/M1/_0_  (.A1(\V2/V3/V2/v2 [0]),
    .A2(\V2/V3/V2/v3 [0]),
    .ZN(\V2/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M1/M1/_1_  (.A(\V2/V3/V2/v2 [0]),
    .B(\V2/V3/V2/v3 [0]),
    .Z(\V2/V3/V2/A1/M1/s1 ));
 AND2_X1 \V2/V3/V2/A1/M1/M2/_0_  (.A1(\V2/V3/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M1/M2/_1_  (.A(\V2/V3/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/V2/s1 [0]));
 OR2_X1 \V2/V3/V2/A1/M1/_0_  (.A1(\V2/V3/V2/A1/M1/c1 ),
    .A2(\V2/V3/V2/A1/M1/c2 ),
    .ZN(\V2/V3/V2/A1/c1 ));
 AND2_X1 \V2/V3/V2/A1/M2/M1/_0_  (.A1(\V2/V3/V2/v2 [1]),
    .A2(\V2/V3/V2/v3 [1]),
    .ZN(\V2/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M2/M1/_1_  (.A(\V2/V3/V2/v2 [1]),
    .B(\V2/V3/V2/v3 [1]),
    .Z(\V2/V3/V2/A1/M2/s1 ));
 AND2_X1 \V2/V3/V2/A1/M2/M2/_0_  (.A1(\V2/V3/V2/A1/M2/s1 ),
    .A2(\V2/V3/V2/A1/c1 ),
    .ZN(\V2/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M2/M2/_1_  (.A(\V2/V3/V2/A1/M2/s1 ),
    .B(\V2/V3/V2/A1/c1 ),
    .Z(\V2/V3/V2/s1 [1]));
 OR2_X1 \V2/V3/V2/A1/M2/_0_  (.A1(\V2/V3/V2/A1/M2/c1 ),
    .A2(\V2/V3/V2/A1/M2/c2 ),
    .ZN(\V2/V3/V2/A1/c2 ));
 AND2_X1 \V2/V3/V2/A1/M3/M1/_0_  (.A1(\V2/V3/V2/v2 [2]),
    .A2(\V2/V3/V2/v3 [2]),
    .ZN(\V2/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M3/M1/_1_  (.A(\V2/V3/V2/v2 [2]),
    .B(\V2/V3/V2/v3 [2]),
    .Z(\V2/V3/V2/A1/M3/s1 ));
 AND2_X1 \V2/V3/V2/A1/M3/M2/_0_  (.A1(\V2/V3/V2/A1/M3/s1 ),
    .A2(\V2/V3/V2/A1/c2 ),
    .ZN(\V2/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M3/M2/_1_  (.A(\V2/V3/V2/A1/M3/s1 ),
    .B(\V2/V3/V2/A1/c2 ),
    .Z(\V2/V3/V2/s1 [2]));
 OR2_X1 \V2/V3/V2/A1/M3/_0_  (.A1(\V2/V3/V2/A1/M3/c1 ),
    .A2(\V2/V3/V2/A1/M3/c2 ),
    .ZN(\V2/V3/V2/A1/c3 ));
 AND2_X1 \V2/V3/V2/A1/M4/M1/_0_  (.A1(\V2/V3/V2/v2 [3]),
    .A2(\V2/V3/V2/v3 [3]),
    .ZN(\V2/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M4/M1/_1_  (.A(\V2/V3/V2/v2 [3]),
    .B(\V2/V3/V2/v3 [3]),
    .Z(\V2/V3/V2/A1/M4/s1 ));
 AND2_X1 \V2/V3/V2/A1/M4/M2/_0_  (.A1(\V2/V3/V2/A1/M4/s1 ),
    .A2(\V2/V3/V2/A1/c3 ),
    .ZN(\V2/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M4/M2/_1_  (.A(\V2/V3/V2/A1/M4/s1 ),
    .B(\V2/V3/V2/A1/c3 ),
    .Z(\V2/V3/V2/s1 [3]));
 OR2_X1 \V2/V3/V2/A1/M4/_0_  (.A1(\V2/V3/V2/A1/M4/c1 ),
    .A2(\V2/V3/V2/A1/M4/c2 ),
    .ZN(\V2/V3/V2/c1 ));
 AND2_X1 \V2/V3/V2/A2/M1/M1/_0_  (.A1(\V2/V3/V2/s1 [0]),
    .A2(\V2/V3/V2/v1 [2]),
    .ZN(\V2/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M1/M1/_1_  (.A(\V2/V3/V2/s1 [0]),
    .B(\V2/V3/V2/v1 [2]),
    .Z(\V2/V3/V2/A2/M1/s1 ));
 AND2_X1 \V2/V3/V2/A2/M1/M2/_0_  (.A1(\V2/V3/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M1/M2/_1_  (.A(\V2/V3/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v2 [2]));
 OR2_X1 \V2/V3/V2/A2/M1/_0_  (.A1(\V2/V3/V2/A2/M1/c1 ),
    .A2(\V2/V3/V2/A2/M1/c2 ),
    .ZN(\V2/V3/V2/A2/c1 ));
 AND2_X1 \V2/V3/V2/A2/M2/M1/_0_  (.A1(\V2/V3/V2/s1 [1]),
    .A2(\V2/V3/V2/v1 [3]),
    .ZN(\V2/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M2/M1/_1_  (.A(\V2/V3/V2/s1 [1]),
    .B(\V2/V3/V2/v1 [3]),
    .Z(\V2/V3/V2/A2/M2/s1 ));
 AND2_X1 \V2/V3/V2/A2/M2/M2/_0_  (.A1(\V2/V3/V2/A2/M2/s1 ),
    .A2(\V2/V3/V2/A2/c1 ),
    .ZN(\V2/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M2/M2/_1_  (.A(\V2/V3/V2/A2/M2/s1 ),
    .B(\V2/V3/V2/A2/c1 ),
    .Z(\V2/V3/v2 [3]));
 OR2_X1 \V2/V3/V2/A2/M2/_0_  (.A1(\V2/V3/V2/A2/M2/c1 ),
    .A2(\V2/V3/V2/A2/M2/c2 ),
    .ZN(\V2/V3/V2/A2/c2 ));
 AND2_X1 \V2/V3/V2/A2/M3/M1/_0_  (.A1(\V2/V3/V2/s1 [2]),
    .A2(ground),
    .ZN(\V2/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M3/M1/_1_  (.A(\V2/V3/V2/s1 [2]),
    .B(ground),
    .Z(\V2/V3/V2/A2/M3/s1 ));
 AND2_X1 \V2/V3/V2/A2/M3/M2/_0_  (.A1(\V2/V3/V2/A2/M3/s1 ),
    .A2(\V2/V3/V2/A2/c2 ),
    .ZN(\V2/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M3/M2/_1_  (.A(\V2/V3/V2/A2/M3/s1 ),
    .B(\V2/V3/V2/A2/c2 ),
    .Z(\V2/V3/V2/s2 [2]));
 OR2_X1 \V2/V3/V2/A2/M3/_0_  (.A1(\V2/V3/V2/A2/M3/c1 ),
    .A2(\V2/V3/V2/A2/M3/c2 ),
    .ZN(\V2/V3/V2/A2/c3 ));
 AND2_X1 \V2/V3/V2/A2/M4/M1/_0_  (.A1(\V2/V3/V2/s1 [3]),
    .A2(ground),
    .ZN(\V2/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M4/M1/_1_  (.A(\V2/V3/V2/s1 [3]),
    .B(ground),
    .Z(\V2/V3/V2/A2/M4/s1 ));
 AND2_X1 \V2/V3/V2/A2/M4/M2/_0_  (.A1(\V2/V3/V2/A2/M4/s1 ),
    .A2(\V2/V3/V2/A2/c3 ),
    .ZN(\V2/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M4/M2/_1_  (.A(\V2/V3/V2/A2/M4/s1 ),
    .B(\V2/V3/V2/A2/c3 ),
    .Z(\V2/V3/V2/s2 [3]));
 OR2_X1 \V2/V3/V2/A2/M4/_0_  (.A1(\V2/V3/V2/A2/M4/c1 ),
    .A2(\V2/V3/V2/A2/M4/c2 ),
    .ZN(\V2/V3/V2/c2 ));
 AND2_X1 \V2/V3/V2/A3/M1/M1/_0_  (.A1(\V2/V3/V2/v4 [0]),
    .A2(\V2/V3/V2/s2 [2]),
    .ZN(\V2/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M1/M1/_1_  (.A(\V2/V3/V2/v4 [0]),
    .B(\V2/V3/V2/s2 [2]),
    .Z(\V2/V3/V2/A3/M1/s1 ));
 AND2_X1 \V2/V3/V2/A3/M1/M2/_0_  (.A1(\V2/V3/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M1/M2/_1_  (.A(\V2/V3/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v2 [4]));
 OR2_X1 \V2/V3/V2/A3/M1/_0_  (.A1(\V2/V3/V2/A3/M1/c1 ),
    .A2(\V2/V3/V2/A3/M1/c2 ),
    .ZN(\V2/V3/V2/A3/c1 ));
 AND2_X1 \V2/V3/V2/A3/M2/M1/_0_  (.A1(\V2/V3/V2/v4 [1]),
    .A2(\V2/V3/V2/s2 [3]),
    .ZN(\V2/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M2/M1/_1_  (.A(\V2/V3/V2/v4 [1]),
    .B(\V2/V3/V2/s2 [3]),
    .Z(\V2/V3/V2/A3/M2/s1 ));
 AND2_X1 \V2/V3/V2/A3/M2/M2/_0_  (.A1(\V2/V3/V2/A3/M2/s1 ),
    .A2(\V2/V3/V2/A3/c1 ),
    .ZN(\V2/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M2/M2/_1_  (.A(\V2/V3/V2/A3/M2/s1 ),
    .B(\V2/V3/V2/A3/c1 ),
    .Z(\V2/V3/v2 [5]));
 OR2_X1 \V2/V3/V2/A3/M2/_0_  (.A1(\V2/V3/V2/A3/M2/c1 ),
    .A2(\V2/V3/V2/A3/M2/c2 ),
    .ZN(\V2/V3/V2/A3/c2 ));
 AND2_X1 \V2/V3/V2/A3/M3/M1/_0_  (.A1(\V2/V3/V2/v4 [2]),
    .A2(\V2/V3/V2/c3 ),
    .ZN(\V2/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M3/M1/_1_  (.A(\V2/V3/V2/v4 [2]),
    .B(\V2/V3/V2/c3 ),
    .Z(\V2/V3/V2/A3/M3/s1 ));
 AND2_X1 \V2/V3/V2/A3/M3/M2/_0_  (.A1(\V2/V3/V2/A3/M3/s1 ),
    .A2(\V2/V3/V2/A3/c2 ),
    .ZN(\V2/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M3/M2/_1_  (.A(\V2/V3/V2/A3/M3/s1 ),
    .B(\V2/V3/V2/A3/c2 ),
    .Z(\V2/V3/v2 [6]));
 OR2_X1 \V2/V3/V2/A3/M3/_0_  (.A1(\V2/V3/V2/A3/M3/c1 ),
    .A2(\V2/V3/V2/A3/M3/c2 ),
    .ZN(\V2/V3/V2/A3/c3 ));
 AND2_X1 \V2/V3/V2/A3/M4/M1/_0_  (.A1(\V2/V3/V2/v4 [3]),
    .A2(ground),
    .ZN(\V2/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M4/M1/_1_  (.A(\V2/V3/V2/v4 [3]),
    .B(ground),
    .Z(\V2/V3/V2/A3/M4/s1 ));
 AND2_X1 \V2/V3/V2/A3/M4/M2/_0_  (.A1(\V2/V3/V2/A3/M4/s1 ),
    .A2(\V2/V3/V2/A3/c3 ),
    .ZN(\V2/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M4/M2/_1_  (.A(\V2/V3/V2/A3/M4/s1 ),
    .B(\V2/V3/V2/A3/c3 ),
    .Z(\V2/V3/v2 [7]));
 OR2_X1 \V2/V3/V2/A3/M4/_0_  (.A1(\V2/V3/V2/A3/M4/c1 ),
    .A2(\V2/V3/V2/A3/M4/c2 ),
    .ZN(\V2/V3/V2/overflow ));
 AND2_X1 \V2/V3/V2/V1/HA1/_0_  (.A1(\V2/V3/V2/V1/w2 ),
    .A2(\V2/V3/V2/V1/w1 ),
    .ZN(\V2/V3/V2/V1/w4 ));
 XOR2_X2 \V2/V3/V2/V1/HA1/_1_  (.A(\V2/V3/V2/V1/w2 ),
    .B(\V2/V3/V2/V1/w1 ),
    .Z(\V2/V3/v2 [1]));
 AND2_X1 \V2/V3/V2/V1/HA2/_0_  (.A1(\V2/V3/V2/V1/w4 ),
    .A2(\V2/V3/V2/V1/w3 ),
    .ZN(\V2/V3/V2/v1 [3]));
 XOR2_X2 \V2/V3/V2/V1/HA2/_1_  (.A(\V2/V3/V2/V1/w4 ),
    .B(\V2/V3/V2/V1/w3 ),
    .Z(\V2/V3/V2/v1 [2]));
 AND2_X1 \V2/V3/V2/V1/_0_  (.A1(A[20]),
    .A2(B[8]),
    .ZN(\V2/V3/v2 [0]));
 AND2_X1 \V2/V3/V2/V1/_1_  (.A1(A[20]),
    .A2(B[9]),
    .ZN(\V2/V3/V2/V1/w1 ));
 AND2_X1 \V2/V3/V2/V1/_2_  (.A1(B[8]),
    .A2(A[21]),
    .ZN(\V2/V3/V2/V1/w2 ));
 AND2_X1 \V2/V3/V2/V1/_3_  (.A1(B[9]),
    .A2(A[21]),
    .ZN(\V2/V3/V2/V1/w3 ));
 AND2_X1 \V2/V3/V2/V2/HA1/_0_  (.A1(\V2/V3/V2/V2/w2 ),
    .A2(\V2/V3/V2/V2/w1 ),
    .ZN(\V2/V3/V2/V2/w4 ));
 XOR2_X2 \V2/V3/V2/V2/HA1/_1_  (.A(\V2/V3/V2/V2/w2 ),
    .B(\V2/V3/V2/V2/w1 ),
    .Z(\V2/V3/V2/v2 [1]));
 AND2_X1 \V2/V3/V2/V2/HA2/_0_  (.A1(\V2/V3/V2/V2/w4 ),
    .A2(\V2/V3/V2/V2/w3 ),
    .ZN(\V2/V3/V2/v2 [3]));
 XOR2_X2 \V2/V3/V2/V2/HA2/_1_  (.A(\V2/V3/V2/V2/w4 ),
    .B(\V2/V3/V2/V2/w3 ),
    .Z(\V2/V3/V2/v2 [2]));
 AND2_X1 \V2/V3/V2/V2/_0_  (.A1(A[22]),
    .A2(B[8]),
    .ZN(\V2/V3/V2/v2 [0]));
 AND2_X1 \V2/V3/V2/V2/_1_  (.A1(A[22]),
    .A2(B[9]),
    .ZN(\V2/V3/V2/V2/w1 ));
 AND2_X1 \V2/V3/V2/V2/_2_  (.A1(B[8]),
    .A2(A[23]),
    .ZN(\V2/V3/V2/V2/w2 ));
 AND2_X1 \V2/V3/V2/V2/_3_  (.A1(B[9]),
    .A2(A[23]),
    .ZN(\V2/V3/V2/V2/w3 ));
 AND2_X1 \V2/V3/V2/V3/HA1/_0_  (.A1(\V2/V3/V2/V3/w2 ),
    .A2(\V2/V3/V2/V3/w1 ),
    .ZN(\V2/V3/V2/V3/w4 ));
 XOR2_X2 \V2/V3/V2/V3/HA1/_1_  (.A(\V2/V3/V2/V3/w2 ),
    .B(\V2/V3/V2/V3/w1 ),
    .Z(\V2/V3/V2/v3 [1]));
 AND2_X1 \V2/V3/V2/V3/HA2/_0_  (.A1(\V2/V3/V2/V3/w4 ),
    .A2(\V2/V3/V2/V3/w3 ),
    .ZN(\V2/V3/V2/v3 [3]));
 XOR2_X2 \V2/V3/V2/V3/HA2/_1_  (.A(\V2/V3/V2/V3/w4 ),
    .B(\V2/V3/V2/V3/w3 ),
    .Z(\V2/V3/V2/v3 [2]));
 AND2_X1 \V2/V3/V2/V3/_0_  (.A1(A[20]),
    .A2(B[10]),
    .ZN(\V2/V3/V2/v3 [0]));
 AND2_X1 \V2/V3/V2/V3/_1_  (.A1(A[20]),
    .A2(B[11]),
    .ZN(\V2/V3/V2/V3/w1 ));
 AND2_X1 \V2/V3/V2/V3/_2_  (.A1(B[10]),
    .A2(A[21]),
    .ZN(\V2/V3/V2/V3/w2 ));
 AND2_X1 \V2/V3/V2/V3/_3_  (.A1(B[11]),
    .A2(A[21]),
    .ZN(\V2/V3/V2/V3/w3 ));
 AND2_X1 \V2/V3/V2/V4/HA1/_0_  (.A1(\V2/V3/V2/V4/w2 ),
    .A2(\V2/V3/V2/V4/w1 ),
    .ZN(\V2/V3/V2/V4/w4 ));
 XOR2_X2 \V2/V3/V2/V4/HA1/_1_  (.A(\V2/V3/V2/V4/w2 ),
    .B(\V2/V3/V2/V4/w1 ),
    .Z(\V2/V3/V2/v4 [1]));
 AND2_X1 \V2/V3/V2/V4/HA2/_0_  (.A1(\V2/V3/V2/V4/w4 ),
    .A2(\V2/V3/V2/V4/w3 ),
    .ZN(\V2/V3/V2/v4 [3]));
 XOR2_X2 \V2/V3/V2/V4/HA2/_1_  (.A(\V2/V3/V2/V4/w4 ),
    .B(\V2/V3/V2/V4/w3 ),
    .Z(\V2/V3/V2/v4 [2]));
 AND2_X1 \V2/V3/V2/V4/_0_  (.A1(A[22]),
    .A2(B[10]),
    .ZN(\V2/V3/V2/v4 [0]));
 AND2_X1 \V2/V3/V2/V4/_1_  (.A1(A[22]),
    .A2(B[11]),
    .ZN(\V2/V3/V2/V4/w1 ));
 AND2_X1 \V2/V3/V2/V4/_2_  (.A1(B[10]),
    .A2(A[23]),
    .ZN(\V2/V3/V2/V4/w2 ));
 AND2_X1 \V2/V3/V2/V4/_3_  (.A1(B[11]),
    .A2(A[23]),
    .ZN(\V2/V3/V2/V4/w3 ));
 OR2_X1 \V2/V3/V2/_0_  (.A1(\V2/V3/V2/c1 ),
    .A2(\V2/V3/V2/c2 ),
    .ZN(\V2/V3/V2/c3 ));
 AND2_X1 \V2/V3/V3/A1/M1/M1/_0_  (.A1(\V2/V3/V3/v2 [0]),
    .A2(\V2/V3/V3/v3 [0]),
    .ZN(\V2/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M1/M1/_1_  (.A(\V2/V3/V3/v2 [0]),
    .B(\V2/V3/V3/v3 [0]),
    .Z(\V2/V3/V3/A1/M1/s1 ));
 AND2_X1 \V2/V3/V3/A1/M1/M2/_0_  (.A1(\V2/V3/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M1/M2/_1_  (.A(\V2/V3/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/V3/s1 [0]));
 OR2_X1 \V2/V3/V3/A1/M1/_0_  (.A1(\V2/V3/V3/A1/M1/c1 ),
    .A2(\V2/V3/V3/A1/M1/c2 ),
    .ZN(\V2/V3/V3/A1/c1 ));
 AND2_X1 \V2/V3/V3/A1/M2/M1/_0_  (.A1(\V2/V3/V3/v2 [1]),
    .A2(\V2/V3/V3/v3 [1]),
    .ZN(\V2/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M2/M1/_1_  (.A(\V2/V3/V3/v2 [1]),
    .B(\V2/V3/V3/v3 [1]),
    .Z(\V2/V3/V3/A1/M2/s1 ));
 AND2_X1 \V2/V3/V3/A1/M2/M2/_0_  (.A1(\V2/V3/V3/A1/M2/s1 ),
    .A2(\V2/V3/V3/A1/c1 ),
    .ZN(\V2/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M2/M2/_1_  (.A(\V2/V3/V3/A1/M2/s1 ),
    .B(\V2/V3/V3/A1/c1 ),
    .Z(\V2/V3/V3/s1 [1]));
 OR2_X1 \V2/V3/V3/A1/M2/_0_  (.A1(\V2/V3/V3/A1/M2/c1 ),
    .A2(\V2/V3/V3/A1/M2/c2 ),
    .ZN(\V2/V3/V3/A1/c2 ));
 AND2_X1 \V2/V3/V3/A1/M3/M1/_0_  (.A1(\V2/V3/V3/v2 [2]),
    .A2(\V2/V3/V3/v3 [2]),
    .ZN(\V2/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M3/M1/_1_  (.A(\V2/V3/V3/v2 [2]),
    .B(\V2/V3/V3/v3 [2]),
    .Z(\V2/V3/V3/A1/M3/s1 ));
 AND2_X1 \V2/V3/V3/A1/M3/M2/_0_  (.A1(\V2/V3/V3/A1/M3/s1 ),
    .A2(\V2/V3/V3/A1/c2 ),
    .ZN(\V2/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M3/M2/_1_  (.A(\V2/V3/V3/A1/M3/s1 ),
    .B(\V2/V3/V3/A1/c2 ),
    .Z(\V2/V3/V3/s1 [2]));
 OR2_X1 \V2/V3/V3/A1/M3/_0_  (.A1(\V2/V3/V3/A1/M3/c1 ),
    .A2(\V2/V3/V3/A1/M3/c2 ),
    .ZN(\V2/V3/V3/A1/c3 ));
 AND2_X1 \V2/V3/V3/A1/M4/M1/_0_  (.A1(\V2/V3/V3/v2 [3]),
    .A2(\V2/V3/V3/v3 [3]),
    .ZN(\V2/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M4/M1/_1_  (.A(\V2/V3/V3/v2 [3]),
    .B(\V2/V3/V3/v3 [3]),
    .Z(\V2/V3/V3/A1/M4/s1 ));
 AND2_X1 \V2/V3/V3/A1/M4/M2/_0_  (.A1(\V2/V3/V3/A1/M4/s1 ),
    .A2(\V2/V3/V3/A1/c3 ),
    .ZN(\V2/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M4/M2/_1_  (.A(\V2/V3/V3/A1/M4/s1 ),
    .B(\V2/V3/V3/A1/c3 ),
    .Z(\V2/V3/V3/s1 [3]));
 OR2_X1 \V2/V3/V3/A1/M4/_0_  (.A1(\V2/V3/V3/A1/M4/c1 ),
    .A2(\V2/V3/V3/A1/M4/c2 ),
    .ZN(\V2/V3/V3/c1 ));
 AND2_X1 \V2/V3/V3/A2/M1/M1/_0_  (.A1(\V2/V3/V3/s1 [0]),
    .A2(\V2/V3/V3/v1 [2]),
    .ZN(\V2/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M1/M1/_1_  (.A(\V2/V3/V3/s1 [0]),
    .B(\V2/V3/V3/v1 [2]),
    .Z(\V2/V3/V3/A2/M1/s1 ));
 AND2_X1 \V2/V3/V3/A2/M1/M2/_0_  (.A1(\V2/V3/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M1/M2/_1_  (.A(\V2/V3/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v3 [2]));
 OR2_X1 \V2/V3/V3/A2/M1/_0_  (.A1(\V2/V3/V3/A2/M1/c1 ),
    .A2(\V2/V3/V3/A2/M1/c2 ),
    .ZN(\V2/V3/V3/A2/c1 ));
 AND2_X1 \V2/V3/V3/A2/M2/M1/_0_  (.A1(\V2/V3/V3/s1 [1]),
    .A2(\V2/V3/V3/v1 [3]),
    .ZN(\V2/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M2/M1/_1_  (.A(\V2/V3/V3/s1 [1]),
    .B(\V2/V3/V3/v1 [3]),
    .Z(\V2/V3/V3/A2/M2/s1 ));
 AND2_X1 \V2/V3/V3/A2/M2/M2/_0_  (.A1(\V2/V3/V3/A2/M2/s1 ),
    .A2(\V2/V3/V3/A2/c1 ),
    .ZN(\V2/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M2/M2/_1_  (.A(\V2/V3/V3/A2/M2/s1 ),
    .B(\V2/V3/V3/A2/c1 ),
    .Z(\V2/V3/v3 [3]));
 OR2_X1 \V2/V3/V3/A2/M2/_0_  (.A1(\V2/V3/V3/A2/M2/c1 ),
    .A2(\V2/V3/V3/A2/M2/c2 ),
    .ZN(\V2/V3/V3/A2/c2 ));
 AND2_X1 \V2/V3/V3/A2/M3/M1/_0_  (.A1(\V2/V3/V3/s1 [2]),
    .A2(ground),
    .ZN(\V2/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M3/M1/_1_  (.A(\V2/V3/V3/s1 [2]),
    .B(ground),
    .Z(\V2/V3/V3/A2/M3/s1 ));
 AND2_X1 \V2/V3/V3/A2/M3/M2/_0_  (.A1(\V2/V3/V3/A2/M3/s1 ),
    .A2(\V2/V3/V3/A2/c2 ),
    .ZN(\V2/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M3/M2/_1_  (.A(\V2/V3/V3/A2/M3/s1 ),
    .B(\V2/V3/V3/A2/c2 ),
    .Z(\V2/V3/V3/s2 [2]));
 OR2_X1 \V2/V3/V3/A2/M3/_0_  (.A1(\V2/V3/V3/A2/M3/c1 ),
    .A2(\V2/V3/V3/A2/M3/c2 ),
    .ZN(\V2/V3/V3/A2/c3 ));
 AND2_X1 \V2/V3/V3/A2/M4/M1/_0_  (.A1(\V2/V3/V3/s1 [3]),
    .A2(ground),
    .ZN(\V2/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M4/M1/_1_  (.A(\V2/V3/V3/s1 [3]),
    .B(ground),
    .Z(\V2/V3/V3/A2/M4/s1 ));
 AND2_X1 \V2/V3/V3/A2/M4/M2/_0_  (.A1(\V2/V3/V3/A2/M4/s1 ),
    .A2(\V2/V3/V3/A2/c3 ),
    .ZN(\V2/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M4/M2/_1_  (.A(\V2/V3/V3/A2/M4/s1 ),
    .B(\V2/V3/V3/A2/c3 ),
    .Z(\V2/V3/V3/s2 [3]));
 OR2_X1 \V2/V3/V3/A2/M4/_0_  (.A1(\V2/V3/V3/A2/M4/c1 ),
    .A2(\V2/V3/V3/A2/M4/c2 ),
    .ZN(\V2/V3/V3/c2 ));
 AND2_X1 \V2/V3/V3/A3/M1/M1/_0_  (.A1(\V2/V3/V3/v4 [0]),
    .A2(\V2/V3/V3/s2 [2]),
    .ZN(\V2/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M1/M1/_1_  (.A(\V2/V3/V3/v4 [0]),
    .B(\V2/V3/V3/s2 [2]),
    .Z(\V2/V3/V3/A3/M1/s1 ));
 AND2_X1 \V2/V3/V3/A3/M1/M2/_0_  (.A1(\V2/V3/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M1/M2/_1_  (.A(\V2/V3/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v3 [4]));
 OR2_X1 \V2/V3/V3/A3/M1/_0_  (.A1(\V2/V3/V3/A3/M1/c1 ),
    .A2(\V2/V3/V3/A3/M1/c2 ),
    .ZN(\V2/V3/V3/A3/c1 ));
 AND2_X1 \V2/V3/V3/A3/M2/M1/_0_  (.A1(\V2/V3/V3/v4 [1]),
    .A2(\V2/V3/V3/s2 [3]),
    .ZN(\V2/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M2/M1/_1_  (.A(\V2/V3/V3/v4 [1]),
    .B(\V2/V3/V3/s2 [3]),
    .Z(\V2/V3/V3/A3/M2/s1 ));
 AND2_X1 \V2/V3/V3/A3/M2/M2/_0_  (.A1(\V2/V3/V3/A3/M2/s1 ),
    .A2(\V2/V3/V3/A3/c1 ),
    .ZN(\V2/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M2/M2/_1_  (.A(\V2/V3/V3/A3/M2/s1 ),
    .B(\V2/V3/V3/A3/c1 ),
    .Z(\V2/V3/v3 [5]));
 OR2_X1 \V2/V3/V3/A3/M2/_0_  (.A1(\V2/V3/V3/A3/M2/c1 ),
    .A2(\V2/V3/V3/A3/M2/c2 ),
    .ZN(\V2/V3/V3/A3/c2 ));
 AND2_X1 \V2/V3/V3/A3/M3/M1/_0_  (.A1(\V2/V3/V3/v4 [2]),
    .A2(\V2/V3/V3/c3 ),
    .ZN(\V2/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M3/M1/_1_  (.A(\V2/V3/V3/v4 [2]),
    .B(\V2/V3/V3/c3 ),
    .Z(\V2/V3/V3/A3/M3/s1 ));
 AND2_X1 \V2/V3/V3/A3/M3/M2/_0_  (.A1(\V2/V3/V3/A3/M3/s1 ),
    .A2(\V2/V3/V3/A3/c2 ),
    .ZN(\V2/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M3/M2/_1_  (.A(\V2/V3/V3/A3/M3/s1 ),
    .B(\V2/V3/V3/A3/c2 ),
    .Z(\V2/V3/v3 [6]));
 OR2_X1 \V2/V3/V3/A3/M3/_0_  (.A1(\V2/V3/V3/A3/M3/c1 ),
    .A2(\V2/V3/V3/A3/M3/c2 ),
    .ZN(\V2/V3/V3/A3/c3 ));
 AND2_X1 \V2/V3/V3/A3/M4/M1/_0_  (.A1(\V2/V3/V3/v4 [3]),
    .A2(ground),
    .ZN(\V2/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M4/M1/_1_  (.A(\V2/V3/V3/v4 [3]),
    .B(ground),
    .Z(\V2/V3/V3/A3/M4/s1 ));
 AND2_X1 \V2/V3/V3/A3/M4/M2/_0_  (.A1(\V2/V3/V3/A3/M4/s1 ),
    .A2(\V2/V3/V3/A3/c3 ),
    .ZN(\V2/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M4/M2/_1_  (.A(\V2/V3/V3/A3/M4/s1 ),
    .B(\V2/V3/V3/A3/c3 ),
    .Z(\V2/V3/v3 [7]));
 OR2_X1 \V2/V3/V3/A3/M4/_0_  (.A1(\V2/V3/V3/A3/M4/c1 ),
    .A2(\V2/V3/V3/A3/M4/c2 ),
    .ZN(\V2/V3/V3/overflow ));
 AND2_X1 \V2/V3/V3/V1/HA1/_0_  (.A1(\V2/V3/V3/V1/w2 ),
    .A2(\V2/V3/V3/V1/w1 ),
    .ZN(\V2/V3/V3/V1/w4 ));
 XOR2_X2 \V2/V3/V3/V1/HA1/_1_  (.A(\V2/V3/V3/V1/w2 ),
    .B(\V2/V3/V3/V1/w1 ),
    .Z(\V2/V3/v3 [1]));
 AND2_X1 \V2/V3/V3/V1/HA2/_0_  (.A1(\V2/V3/V3/V1/w4 ),
    .A2(\V2/V3/V3/V1/w3 ),
    .ZN(\V2/V3/V3/v1 [3]));
 XOR2_X2 \V2/V3/V3/V1/HA2/_1_  (.A(\V2/V3/V3/V1/w4 ),
    .B(\V2/V3/V3/V1/w3 ),
    .Z(\V2/V3/V3/v1 [2]));
 AND2_X1 \V2/V3/V3/V1/_0_  (.A1(A[16]),
    .A2(B[12]),
    .ZN(\V2/V3/v3 [0]));
 AND2_X1 \V2/V3/V3/V1/_1_  (.A1(A[16]),
    .A2(B[13]),
    .ZN(\V2/V3/V3/V1/w1 ));
 AND2_X1 \V2/V3/V3/V1/_2_  (.A1(B[12]),
    .A2(A[17]),
    .ZN(\V2/V3/V3/V1/w2 ));
 AND2_X1 \V2/V3/V3/V1/_3_  (.A1(B[13]),
    .A2(A[17]),
    .ZN(\V2/V3/V3/V1/w3 ));
 AND2_X1 \V2/V3/V3/V2/HA1/_0_  (.A1(\V2/V3/V3/V2/w2 ),
    .A2(\V2/V3/V3/V2/w1 ),
    .ZN(\V2/V3/V3/V2/w4 ));
 XOR2_X2 \V2/V3/V3/V2/HA1/_1_  (.A(\V2/V3/V3/V2/w2 ),
    .B(\V2/V3/V3/V2/w1 ),
    .Z(\V2/V3/V3/v2 [1]));
 AND2_X1 \V2/V3/V3/V2/HA2/_0_  (.A1(\V2/V3/V3/V2/w4 ),
    .A2(\V2/V3/V3/V2/w3 ),
    .ZN(\V2/V3/V3/v2 [3]));
 XOR2_X2 \V2/V3/V3/V2/HA2/_1_  (.A(\V2/V3/V3/V2/w4 ),
    .B(\V2/V3/V3/V2/w3 ),
    .Z(\V2/V3/V3/v2 [2]));
 AND2_X1 \V2/V3/V3/V2/_0_  (.A1(A[18]),
    .A2(B[12]),
    .ZN(\V2/V3/V3/v2 [0]));
 AND2_X1 \V2/V3/V3/V2/_1_  (.A1(A[18]),
    .A2(B[13]),
    .ZN(\V2/V3/V3/V2/w1 ));
 AND2_X1 \V2/V3/V3/V2/_2_  (.A1(B[12]),
    .A2(A[19]),
    .ZN(\V2/V3/V3/V2/w2 ));
 AND2_X1 \V2/V3/V3/V2/_3_  (.A1(B[13]),
    .A2(A[19]),
    .ZN(\V2/V3/V3/V2/w3 ));
 AND2_X1 \V2/V3/V3/V3/HA1/_0_  (.A1(\V2/V3/V3/V3/w2 ),
    .A2(\V2/V3/V3/V3/w1 ),
    .ZN(\V2/V3/V3/V3/w4 ));
 XOR2_X2 \V2/V3/V3/V3/HA1/_1_  (.A(\V2/V3/V3/V3/w2 ),
    .B(\V2/V3/V3/V3/w1 ),
    .Z(\V2/V3/V3/v3 [1]));
 AND2_X1 \V2/V3/V3/V3/HA2/_0_  (.A1(\V2/V3/V3/V3/w4 ),
    .A2(\V2/V3/V3/V3/w3 ),
    .ZN(\V2/V3/V3/v3 [3]));
 XOR2_X2 \V2/V3/V3/V3/HA2/_1_  (.A(\V2/V3/V3/V3/w4 ),
    .B(\V2/V3/V3/V3/w3 ),
    .Z(\V2/V3/V3/v3 [2]));
 AND2_X1 \V2/V3/V3/V3/_0_  (.A1(A[16]),
    .A2(B[14]),
    .ZN(\V2/V3/V3/v3 [0]));
 AND2_X1 \V2/V3/V3/V3/_1_  (.A1(A[16]),
    .A2(B[15]),
    .ZN(\V2/V3/V3/V3/w1 ));
 AND2_X1 \V2/V3/V3/V3/_2_  (.A1(B[14]),
    .A2(A[17]),
    .ZN(\V2/V3/V3/V3/w2 ));
 AND2_X1 \V2/V3/V3/V3/_3_  (.A1(B[15]),
    .A2(A[17]),
    .ZN(\V2/V3/V3/V3/w3 ));
 AND2_X1 \V2/V3/V3/V4/HA1/_0_  (.A1(\V2/V3/V3/V4/w2 ),
    .A2(\V2/V3/V3/V4/w1 ),
    .ZN(\V2/V3/V3/V4/w4 ));
 XOR2_X2 \V2/V3/V3/V4/HA1/_1_  (.A(\V2/V3/V3/V4/w2 ),
    .B(\V2/V3/V3/V4/w1 ),
    .Z(\V2/V3/V3/v4 [1]));
 AND2_X1 \V2/V3/V3/V4/HA2/_0_  (.A1(\V2/V3/V3/V4/w4 ),
    .A2(\V2/V3/V3/V4/w3 ),
    .ZN(\V2/V3/V3/v4 [3]));
 XOR2_X2 \V2/V3/V3/V4/HA2/_1_  (.A(\V2/V3/V3/V4/w4 ),
    .B(\V2/V3/V3/V4/w3 ),
    .Z(\V2/V3/V3/v4 [2]));
 AND2_X1 \V2/V3/V3/V4/_0_  (.A1(A[18]),
    .A2(B[14]),
    .ZN(\V2/V3/V3/v4 [0]));
 AND2_X1 \V2/V3/V3/V4/_1_  (.A1(A[18]),
    .A2(B[15]),
    .ZN(\V2/V3/V3/V4/w1 ));
 AND2_X1 \V2/V3/V3/V4/_2_  (.A1(B[14]),
    .A2(A[19]),
    .ZN(\V2/V3/V3/V4/w2 ));
 AND2_X1 \V2/V3/V3/V4/_3_  (.A1(B[15]),
    .A2(A[19]),
    .ZN(\V2/V3/V3/V4/w3 ));
 OR2_X1 \V2/V3/V3/_0_  (.A1(\V2/V3/V3/c1 ),
    .A2(\V2/V3/V3/c2 ),
    .ZN(\V2/V3/V3/c3 ));
 AND2_X1 \V2/V3/V4/A1/M1/M1/_0_  (.A1(\V2/V3/V4/v2 [0]),
    .A2(\V2/V3/V4/v3 [0]),
    .ZN(\V2/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M1/M1/_1_  (.A(\V2/V3/V4/v2 [0]),
    .B(\V2/V3/V4/v3 [0]),
    .Z(\V2/V3/V4/A1/M1/s1 ));
 AND2_X1 \V2/V3/V4/A1/M1/M2/_0_  (.A1(\V2/V3/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M1/M2/_1_  (.A(\V2/V3/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/V4/s1 [0]));
 OR2_X1 \V2/V3/V4/A1/M1/_0_  (.A1(\V2/V3/V4/A1/M1/c1 ),
    .A2(\V2/V3/V4/A1/M1/c2 ),
    .ZN(\V2/V3/V4/A1/c1 ));
 AND2_X1 \V2/V3/V4/A1/M2/M1/_0_  (.A1(\V2/V3/V4/v2 [1]),
    .A2(\V2/V3/V4/v3 [1]),
    .ZN(\V2/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M2/M1/_1_  (.A(\V2/V3/V4/v2 [1]),
    .B(\V2/V3/V4/v3 [1]),
    .Z(\V2/V3/V4/A1/M2/s1 ));
 AND2_X1 \V2/V3/V4/A1/M2/M2/_0_  (.A1(\V2/V3/V4/A1/M2/s1 ),
    .A2(\V2/V3/V4/A1/c1 ),
    .ZN(\V2/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M2/M2/_1_  (.A(\V2/V3/V4/A1/M2/s1 ),
    .B(\V2/V3/V4/A1/c1 ),
    .Z(\V2/V3/V4/s1 [1]));
 OR2_X1 \V2/V3/V4/A1/M2/_0_  (.A1(\V2/V3/V4/A1/M2/c1 ),
    .A2(\V2/V3/V4/A1/M2/c2 ),
    .ZN(\V2/V3/V4/A1/c2 ));
 AND2_X1 \V2/V3/V4/A1/M3/M1/_0_  (.A1(\V2/V3/V4/v2 [2]),
    .A2(\V2/V3/V4/v3 [2]),
    .ZN(\V2/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M3/M1/_1_  (.A(\V2/V3/V4/v2 [2]),
    .B(\V2/V3/V4/v3 [2]),
    .Z(\V2/V3/V4/A1/M3/s1 ));
 AND2_X1 \V2/V3/V4/A1/M3/M2/_0_  (.A1(\V2/V3/V4/A1/M3/s1 ),
    .A2(\V2/V3/V4/A1/c2 ),
    .ZN(\V2/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M3/M2/_1_  (.A(\V2/V3/V4/A1/M3/s1 ),
    .B(\V2/V3/V4/A1/c2 ),
    .Z(\V2/V3/V4/s1 [2]));
 OR2_X1 \V2/V3/V4/A1/M3/_0_  (.A1(\V2/V3/V4/A1/M3/c1 ),
    .A2(\V2/V3/V4/A1/M3/c2 ),
    .ZN(\V2/V3/V4/A1/c3 ));
 AND2_X1 \V2/V3/V4/A1/M4/M1/_0_  (.A1(\V2/V3/V4/v2 [3]),
    .A2(\V2/V3/V4/v3 [3]),
    .ZN(\V2/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M4/M1/_1_  (.A(\V2/V3/V4/v2 [3]),
    .B(\V2/V3/V4/v3 [3]),
    .Z(\V2/V3/V4/A1/M4/s1 ));
 AND2_X1 \V2/V3/V4/A1/M4/M2/_0_  (.A1(\V2/V3/V4/A1/M4/s1 ),
    .A2(\V2/V3/V4/A1/c3 ),
    .ZN(\V2/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M4/M2/_1_  (.A(\V2/V3/V4/A1/M4/s1 ),
    .B(\V2/V3/V4/A1/c3 ),
    .Z(\V2/V3/V4/s1 [3]));
 OR2_X1 \V2/V3/V4/A1/M4/_0_  (.A1(\V2/V3/V4/A1/M4/c1 ),
    .A2(\V2/V3/V4/A1/M4/c2 ),
    .ZN(\V2/V3/V4/c1 ));
 AND2_X1 \V2/V3/V4/A2/M1/M1/_0_  (.A1(\V2/V3/V4/s1 [0]),
    .A2(\V2/V3/V4/v1 [2]),
    .ZN(\V2/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M1/M1/_1_  (.A(\V2/V3/V4/s1 [0]),
    .B(\V2/V3/V4/v1 [2]),
    .Z(\V2/V3/V4/A2/M1/s1 ));
 AND2_X1 \V2/V3/V4/A2/M1/M2/_0_  (.A1(\V2/V3/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M1/M2/_1_  (.A(\V2/V3/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v4 [2]));
 OR2_X1 \V2/V3/V4/A2/M1/_0_  (.A1(\V2/V3/V4/A2/M1/c1 ),
    .A2(\V2/V3/V4/A2/M1/c2 ),
    .ZN(\V2/V3/V4/A2/c1 ));
 AND2_X1 \V2/V3/V4/A2/M2/M1/_0_  (.A1(\V2/V3/V4/s1 [1]),
    .A2(\V2/V3/V4/v1 [3]),
    .ZN(\V2/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M2/M1/_1_  (.A(\V2/V3/V4/s1 [1]),
    .B(\V2/V3/V4/v1 [3]),
    .Z(\V2/V3/V4/A2/M2/s1 ));
 AND2_X1 \V2/V3/V4/A2/M2/M2/_0_  (.A1(\V2/V3/V4/A2/M2/s1 ),
    .A2(\V2/V3/V4/A2/c1 ),
    .ZN(\V2/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M2/M2/_1_  (.A(\V2/V3/V4/A2/M2/s1 ),
    .B(\V2/V3/V4/A2/c1 ),
    .Z(\V2/V3/v4 [3]));
 OR2_X1 \V2/V3/V4/A2/M2/_0_  (.A1(\V2/V3/V4/A2/M2/c1 ),
    .A2(\V2/V3/V4/A2/M2/c2 ),
    .ZN(\V2/V3/V4/A2/c2 ));
 AND2_X1 \V2/V3/V4/A2/M3/M1/_0_  (.A1(\V2/V3/V4/s1 [2]),
    .A2(ground),
    .ZN(\V2/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M3/M1/_1_  (.A(\V2/V3/V4/s1 [2]),
    .B(ground),
    .Z(\V2/V3/V4/A2/M3/s1 ));
 AND2_X1 \V2/V3/V4/A2/M3/M2/_0_  (.A1(\V2/V3/V4/A2/M3/s1 ),
    .A2(\V2/V3/V4/A2/c2 ),
    .ZN(\V2/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M3/M2/_1_  (.A(\V2/V3/V4/A2/M3/s1 ),
    .B(\V2/V3/V4/A2/c2 ),
    .Z(\V2/V3/V4/s2 [2]));
 OR2_X1 \V2/V3/V4/A2/M3/_0_  (.A1(\V2/V3/V4/A2/M3/c1 ),
    .A2(\V2/V3/V4/A2/M3/c2 ),
    .ZN(\V2/V3/V4/A2/c3 ));
 AND2_X1 \V2/V3/V4/A2/M4/M1/_0_  (.A1(\V2/V3/V4/s1 [3]),
    .A2(ground),
    .ZN(\V2/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M4/M1/_1_  (.A(\V2/V3/V4/s1 [3]),
    .B(ground),
    .Z(\V2/V3/V4/A2/M4/s1 ));
 AND2_X1 \V2/V3/V4/A2/M4/M2/_0_  (.A1(\V2/V3/V4/A2/M4/s1 ),
    .A2(\V2/V3/V4/A2/c3 ),
    .ZN(\V2/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M4/M2/_1_  (.A(\V2/V3/V4/A2/M4/s1 ),
    .B(\V2/V3/V4/A2/c3 ),
    .Z(\V2/V3/V4/s2 [3]));
 OR2_X1 \V2/V3/V4/A2/M4/_0_  (.A1(\V2/V3/V4/A2/M4/c1 ),
    .A2(\V2/V3/V4/A2/M4/c2 ),
    .ZN(\V2/V3/V4/c2 ));
 AND2_X1 \V2/V3/V4/A3/M1/M1/_0_  (.A1(\V2/V3/V4/v4 [0]),
    .A2(\V2/V3/V4/s2 [2]),
    .ZN(\V2/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M1/M1/_1_  (.A(\V2/V3/V4/v4 [0]),
    .B(\V2/V3/V4/s2 [2]),
    .Z(\V2/V3/V4/A3/M1/s1 ));
 AND2_X1 \V2/V3/V4/A3/M1/M2/_0_  (.A1(\V2/V3/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M1/M2/_1_  (.A(\V2/V3/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V3/v4 [4]));
 OR2_X1 \V2/V3/V4/A3/M1/_0_  (.A1(\V2/V3/V4/A3/M1/c1 ),
    .A2(\V2/V3/V4/A3/M1/c2 ),
    .ZN(\V2/V3/V4/A3/c1 ));
 AND2_X1 \V2/V3/V4/A3/M2/M1/_0_  (.A1(\V2/V3/V4/v4 [1]),
    .A2(\V2/V3/V4/s2 [3]),
    .ZN(\V2/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M2/M1/_1_  (.A(\V2/V3/V4/v4 [1]),
    .B(\V2/V3/V4/s2 [3]),
    .Z(\V2/V3/V4/A3/M2/s1 ));
 AND2_X1 \V2/V3/V4/A3/M2/M2/_0_  (.A1(\V2/V3/V4/A3/M2/s1 ),
    .A2(\V2/V3/V4/A3/c1 ),
    .ZN(\V2/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M2/M2/_1_  (.A(\V2/V3/V4/A3/M2/s1 ),
    .B(\V2/V3/V4/A3/c1 ),
    .Z(\V2/V3/v4 [5]));
 OR2_X1 \V2/V3/V4/A3/M2/_0_  (.A1(\V2/V3/V4/A3/M2/c1 ),
    .A2(\V2/V3/V4/A3/M2/c2 ),
    .ZN(\V2/V3/V4/A3/c2 ));
 AND2_X1 \V2/V3/V4/A3/M3/M1/_0_  (.A1(\V2/V3/V4/v4 [2]),
    .A2(\V2/V3/V4/c3 ),
    .ZN(\V2/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M3/M1/_1_  (.A(\V2/V3/V4/v4 [2]),
    .B(\V2/V3/V4/c3 ),
    .Z(\V2/V3/V4/A3/M3/s1 ));
 AND2_X1 \V2/V3/V4/A3/M3/M2/_0_  (.A1(\V2/V3/V4/A3/M3/s1 ),
    .A2(\V2/V3/V4/A3/c2 ),
    .ZN(\V2/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M3/M2/_1_  (.A(\V2/V3/V4/A3/M3/s1 ),
    .B(\V2/V3/V4/A3/c2 ),
    .Z(\V2/V3/v4 [6]));
 OR2_X1 \V2/V3/V4/A3/M3/_0_  (.A1(\V2/V3/V4/A3/M3/c1 ),
    .A2(\V2/V3/V4/A3/M3/c2 ),
    .ZN(\V2/V3/V4/A3/c3 ));
 AND2_X1 \V2/V3/V4/A3/M4/M1/_0_  (.A1(\V2/V3/V4/v4 [3]),
    .A2(ground),
    .ZN(\V2/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M4/M1/_1_  (.A(\V2/V3/V4/v4 [3]),
    .B(ground),
    .Z(\V2/V3/V4/A3/M4/s1 ));
 AND2_X1 \V2/V3/V4/A3/M4/M2/_0_  (.A1(\V2/V3/V4/A3/M4/s1 ),
    .A2(\V2/V3/V4/A3/c3 ),
    .ZN(\V2/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M4/M2/_1_  (.A(\V2/V3/V4/A3/M4/s1 ),
    .B(\V2/V3/V4/A3/c3 ),
    .Z(\V2/V3/v4 [7]));
 OR2_X1 \V2/V3/V4/A3/M4/_0_  (.A1(\V2/V3/V4/A3/M4/c1 ),
    .A2(\V2/V3/V4/A3/M4/c2 ),
    .ZN(\V2/V3/V4/overflow ));
 AND2_X1 \V2/V3/V4/V1/HA1/_0_  (.A1(\V2/V3/V4/V1/w2 ),
    .A2(\V2/V3/V4/V1/w1 ),
    .ZN(\V2/V3/V4/V1/w4 ));
 XOR2_X2 \V2/V3/V4/V1/HA1/_1_  (.A(\V2/V3/V4/V1/w2 ),
    .B(\V2/V3/V4/V1/w1 ),
    .Z(\V2/V3/v4 [1]));
 AND2_X1 \V2/V3/V4/V1/HA2/_0_  (.A1(\V2/V3/V4/V1/w4 ),
    .A2(\V2/V3/V4/V1/w3 ),
    .ZN(\V2/V3/V4/v1 [3]));
 XOR2_X2 \V2/V3/V4/V1/HA2/_1_  (.A(\V2/V3/V4/V1/w4 ),
    .B(\V2/V3/V4/V1/w3 ),
    .Z(\V2/V3/V4/v1 [2]));
 AND2_X1 \V2/V3/V4/V1/_0_  (.A1(A[20]),
    .A2(B[12]),
    .ZN(\V2/V3/v4 [0]));
 AND2_X1 \V2/V3/V4/V1/_1_  (.A1(A[20]),
    .A2(B[13]),
    .ZN(\V2/V3/V4/V1/w1 ));
 AND2_X1 \V2/V3/V4/V1/_2_  (.A1(B[12]),
    .A2(A[21]),
    .ZN(\V2/V3/V4/V1/w2 ));
 AND2_X1 \V2/V3/V4/V1/_3_  (.A1(B[13]),
    .A2(A[21]),
    .ZN(\V2/V3/V4/V1/w3 ));
 AND2_X1 \V2/V3/V4/V2/HA1/_0_  (.A1(\V2/V3/V4/V2/w2 ),
    .A2(\V2/V3/V4/V2/w1 ),
    .ZN(\V2/V3/V4/V2/w4 ));
 XOR2_X2 \V2/V3/V4/V2/HA1/_1_  (.A(\V2/V3/V4/V2/w2 ),
    .B(\V2/V3/V4/V2/w1 ),
    .Z(\V2/V3/V4/v2 [1]));
 AND2_X1 \V2/V3/V4/V2/HA2/_0_  (.A1(\V2/V3/V4/V2/w4 ),
    .A2(\V2/V3/V4/V2/w3 ),
    .ZN(\V2/V3/V4/v2 [3]));
 XOR2_X2 \V2/V3/V4/V2/HA2/_1_  (.A(\V2/V3/V4/V2/w4 ),
    .B(\V2/V3/V4/V2/w3 ),
    .Z(\V2/V3/V4/v2 [2]));
 AND2_X1 \V2/V3/V4/V2/_0_  (.A1(A[22]),
    .A2(B[12]),
    .ZN(\V2/V3/V4/v2 [0]));
 AND2_X1 \V2/V3/V4/V2/_1_  (.A1(A[22]),
    .A2(B[13]),
    .ZN(\V2/V3/V4/V2/w1 ));
 AND2_X1 \V2/V3/V4/V2/_2_  (.A1(B[12]),
    .A2(A[23]),
    .ZN(\V2/V3/V4/V2/w2 ));
 AND2_X1 \V2/V3/V4/V2/_3_  (.A1(B[13]),
    .A2(A[23]),
    .ZN(\V2/V3/V4/V2/w3 ));
 AND2_X1 \V2/V3/V4/V3/HA1/_0_  (.A1(\V2/V3/V4/V3/w2 ),
    .A2(\V2/V3/V4/V3/w1 ),
    .ZN(\V2/V3/V4/V3/w4 ));
 XOR2_X2 \V2/V3/V4/V3/HA1/_1_  (.A(\V2/V3/V4/V3/w2 ),
    .B(\V2/V3/V4/V3/w1 ),
    .Z(\V2/V3/V4/v3 [1]));
 AND2_X1 \V2/V3/V4/V3/HA2/_0_  (.A1(\V2/V3/V4/V3/w4 ),
    .A2(\V2/V3/V4/V3/w3 ),
    .ZN(\V2/V3/V4/v3 [3]));
 XOR2_X2 \V2/V3/V4/V3/HA2/_1_  (.A(\V2/V3/V4/V3/w4 ),
    .B(\V2/V3/V4/V3/w3 ),
    .Z(\V2/V3/V4/v3 [2]));
 AND2_X1 \V2/V3/V4/V3/_0_  (.A1(A[20]),
    .A2(B[14]),
    .ZN(\V2/V3/V4/v3 [0]));
 AND2_X1 \V2/V3/V4/V3/_1_  (.A1(A[20]),
    .A2(B[15]),
    .ZN(\V2/V3/V4/V3/w1 ));
 AND2_X1 \V2/V3/V4/V3/_2_  (.A1(B[14]),
    .A2(A[21]),
    .ZN(\V2/V3/V4/V3/w2 ));
 AND2_X1 \V2/V3/V4/V3/_3_  (.A1(B[15]),
    .A2(A[21]),
    .ZN(\V2/V3/V4/V3/w3 ));
 AND2_X1 \V2/V3/V4/V4/HA1/_0_  (.A1(\V2/V3/V4/V4/w2 ),
    .A2(\V2/V3/V4/V4/w1 ),
    .ZN(\V2/V3/V4/V4/w4 ));
 XOR2_X2 \V2/V3/V4/V4/HA1/_1_  (.A(\V2/V3/V4/V4/w2 ),
    .B(\V2/V3/V4/V4/w1 ),
    .Z(\V2/V3/V4/v4 [1]));
 AND2_X1 \V2/V3/V4/V4/HA2/_0_  (.A1(\V2/V3/V4/V4/w4 ),
    .A2(\V2/V3/V4/V4/w3 ),
    .ZN(\V2/V3/V4/v4 [3]));
 XOR2_X2 \V2/V3/V4/V4/HA2/_1_  (.A(\V2/V3/V4/V4/w4 ),
    .B(\V2/V3/V4/V4/w3 ),
    .Z(\V2/V3/V4/v4 [2]));
 AND2_X1 \V2/V3/V4/V4/_0_  (.A1(A[22]),
    .A2(B[14]),
    .ZN(\V2/V3/V4/v4 [0]));
 AND2_X1 \V2/V3/V4/V4/_1_  (.A1(A[22]),
    .A2(B[15]),
    .ZN(\V2/V3/V4/V4/w1 ));
 AND2_X1 \V2/V3/V4/V4/_2_  (.A1(B[14]),
    .A2(A[23]),
    .ZN(\V2/V3/V4/V4/w2 ));
 AND2_X1 \V2/V3/V4/V4/_3_  (.A1(B[15]),
    .A2(A[23]),
    .ZN(\V2/V3/V4/V4/w3 ));
 OR2_X1 \V2/V3/V4/_0_  (.A1(\V2/V3/V4/c1 ),
    .A2(\V2/V3/V4/c2 ),
    .ZN(\V2/V3/V4/c3 ));
 OR2_X1 \V2/V3/_0_  (.A1(\V2/V3/c1 ),
    .A2(\V2/V3/c2 ),
    .ZN(\V2/V3/c3 ));
 AND2_X1 \V2/V4/A1/A1/M1/M1/_0_  (.A1(\V2/V4/v2 [0]),
    .A2(\V2/V4/v3 [0]),
    .ZN(\V2/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M1/M1/_1_  (.A(\V2/V4/v2 [0]),
    .B(\V2/V4/v3 [0]),
    .Z(\V2/V4/A1/A1/M1/s1 ));
 AND2_X1 \V2/V4/A1/A1/M1/M2/_0_  (.A1(\V2/V4/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M1/M2/_1_  (.A(\V2/V4/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/s1 [0]));
 OR2_X1 \V2/V4/A1/A1/M1/_0_  (.A1(\V2/V4/A1/A1/M1/c1 ),
    .A2(\V2/V4/A1/A1/M1/c2 ),
    .ZN(\V2/V4/A1/A1/c1 ));
 AND2_X1 \V2/V4/A1/A1/M2/M1/_0_  (.A1(\V2/V4/v2 [1]),
    .A2(\V2/V4/v3 [1]),
    .ZN(\V2/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M2/M1/_1_  (.A(\V2/V4/v2 [1]),
    .B(\V2/V4/v3 [1]),
    .Z(\V2/V4/A1/A1/M2/s1 ));
 AND2_X1 \V2/V4/A1/A1/M2/M2/_0_  (.A1(\V2/V4/A1/A1/M2/s1 ),
    .A2(\V2/V4/A1/A1/c1 ),
    .ZN(\V2/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M2/M2/_1_  (.A(\V2/V4/A1/A1/M2/s1 ),
    .B(\V2/V4/A1/A1/c1 ),
    .Z(\V2/V4/s1 [1]));
 OR2_X1 \V2/V4/A1/A1/M2/_0_  (.A1(\V2/V4/A1/A1/M2/c1 ),
    .A2(\V2/V4/A1/A1/M2/c2 ),
    .ZN(\V2/V4/A1/A1/c2 ));
 AND2_X1 \V2/V4/A1/A1/M3/M1/_0_  (.A1(\V2/V4/v2 [2]),
    .A2(\V2/V4/v3 [2]),
    .ZN(\V2/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M3/M1/_1_  (.A(\V2/V4/v2 [2]),
    .B(\V2/V4/v3 [2]),
    .Z(\V2/V4/A1/A1/M3/s1 ));
 AND2_X1 \V2/V4/A1/A1/M3/M2/_0_  (.A1(\V2/V4/A1/A1/M3/s1 ),
    .A2(\V2/V4/A1/A1/c2 ),
    .ZN(\V2/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M3/M2/_1_  (.A(\V2/V4/A1/A1/M3/s1 ),
    .B(\V2/V4/A1/A1/c2 ),
    .Z(\V2/V4/s1 [2]));
 OR2_X1 \V2/V4/A1/A1/M3/_0_  (.A1(\V2/V4/A1/A1/M3/c1 ),
    .A2(\V2/V4/A1/A1/M3/c2 ),
    .ZN(\V2/V4/A1/A1/c3 ));
 AND2_X1 \V2/V4/A1/A1/M4/M1/_0_  (.A1(\V2/V4/v2 [3]),
    .A2(\V2/V4/v3 [3]),
    .ZN(\V2/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M4/M1/_1_  (.A(\V2/V4/v2 [3]),
    .B(\V2/V4/v3 [3]),
    .Z(\V2/V4/A1/A1/M4/s1 ));
 AND2_X1 \V2/V4/A1/A1/M4/M2/_0_  (.A1(\V2/V4/A1/A1/M4/s1 ),
    .A2(\V2/V4/A1/A1/c3 ),
    .ZN(\V2/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M4/M2/_1_  (.A(\V2/V4/A1/A1/M4/s1 ),
    .B(\V2/V4/A1/A1/c3 ),
    .Z(\V2/V4/s1 [3]));
 OR2_X1 \V2/V4/A1/A1/M4/_0_  (.A1(\V2/V4/A1/A1/M4/c1 ),
    .A2(\V2/V4/A1/A1/M4/c2 ),
    .ZN(\V2/V4/A1/c1 ));
 AND2_X1 \V2/V4/A1/A2/M1/M1/_0_  (.A1(\V2/V4/v2 [4]),
    .A2(\V2/V4/v3 [4]),
    .ZN(\V2/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M1/M1/_1_  (.A(\V2/V4/v2 [4]),
    .B(\V2/V4/v3 [4]),
    .Z(\V2/V4/A1/A2/M1/s1 ));
 AND2_X1 \V2/V4/A1/A2/M1/M2/_0_  (.A1(\V2/V4/A1/A2/M1/s1 ),
    .A2(\V2/V4/A1/c1 ),
    .ZN(\V2/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M1/M2/_1_  (.A(\V2/V4/A1/A2/M1/s1 ),
    .B(\V2/V4/A1/c1 ),
    .Z(\V2/V4/s1 [4]));
 OR2_X1 \V2/V4/A1/A2/M1/_0_  (.A1(\V2/V4/A1/A2/M1/c1 ),
    .A2(\V2/V4/A1/A2/M1/c2 ),
    .ZN(\V2/V4/A1/A2/c1 ));
 AND2_X1 \V2/V4/A1/A2/M2/M1/_0_  (.A1(\V2/V4/v2 [5]),
    .A2(\V2/V4/v3 [5]),
    .ZN(\V2/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M2/M1/_1_  (.A(\V2/V4/v2 [5]),
    .B(\V2/V4/v3 [5]),
    .Z(\V2/V4/A1/A2/M2/s1 ));
 AND2_X1 \V2/V4/A1/A2/M2/M2/_0_  (.A1(\V2/V4/A1/A2/M2/s1 ),
    .A2(\V2/V4/A1/A2/c1 ),
    .ZN(\V2/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M2/M2/_1_  (.A(\V2/V4/A1/A2/M2/s1 ),
    .B(\V2/V4/A1/A2/c1 ),
    .Z(\V2/V4/s1 [5]));
 OR2_X1 \V2/V4/A1/A2/M2/_0_  (.A1(\V2/V4/A1/A2/M2/c1 ),
    .A2(\V2/V4/A1/A2/M2/c2 ),
    .ZN(\V2/V4/A1/A2/c2 ));
 AND2_X1 \V2/V4/A1/A2/M3/M1/_0_  (.A1(\V2/V4/v2 [6]),
    .A2(\V2/V4/v3 [6]),
    .ZN(\V2/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M3/M1/_1_  (.A(\V2/V4/v2 [6]),
    .B(\V2/V4/v3 [6]),
    .Z(\V2/V4/A1/A2/M3/s1 ));
 AND2_X1 \V2/V4/A1/A2/M3/M2/_0_  (.A1(\V2/V4/A1/A2/M3/s1 ),
    .A2(\V2/V4/A1/A2/c2 ),
    .ZN(\V2/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M3/M2/_1_  (.A(\V2/V4/A1/A2/M3/s1 ),
    .B(\V2/V4/A1/A2/c2 ),
    .Z(\V2/V4/s1 [6]));
 OR2_X1 \V2/V4/A1/A2/M3/_0_  (.A1(\V2/V4/A1/A2/M3/c1 ),
    .A2(\V2/V4/A1/A2/M3/c2 ),
    .ZN(\V2/V4/A1/A2/c3 ));
 AND2_X1 \V2/V4/A1/A2/M4/M1/_0_  (.A1(\V2/V4/v2 [7]),
    .A2(\V2/V4/v3 [7]),
    .ZN(\V2/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M4/M1/_1_  (.A(\V2/V4/v2 [7]),
    .B(\V2/V4/v3 [7]),
    .Z(\V2/V4/A1/A2/M4/s1 ));
 AND2_X1 \V2/V4/A1/A2/M4/M2/_0_  (.A1(\V2/V4/A1/A2/M4/s1 ),
    .A2(\V2/V4/A1/A2/c3 ),
    .ZN(\V2/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M4/M2/_1_  (.A(\V2/V4/A1/A2/M4/s1 ),
    .B(\V2/V4/A1/A2/c3 ),
    .Z(\V2/V4/s1 [7]));
 OR2_X1 \V2/V4/A1/A2/M4/_0_  (.A1(\V2/V4/A1/A2/M4/c1 ),
    .A2(\V2/V4/A1/A2/M4/c2 ),
    .ZN(\V2/V4/c1 ));
 AND2_X1 \V2/V4/A2/A1/M1/M1/_0_  (.A1(\V2/V4/s1 [0]),
    .A2(\V2/V4/v1 [4]),
    .ZN(\V2/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M1/M1/_1_  (.A(\V2/V4/s1 [0]),
    .B(\V2/V4/v1 [4]),
    .Z(\V2/V4/A2/A1/M1/s1 ));
 AND2_X1 \V2/V4/A2/A1/M1/M2/_0_  (.A1(\V2/V4/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M1/M2/_1_  (.A(\V2/V4/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v4 [4]));
 OR2_X1 \V2/V4/A2/A1/M1/_0_  (.A1(\V2/V4/A2/A1/M1/c1 ),
    .A2(\V2/V4/A2/A1/M1/c2 ),
    .ZN(\V2/V4/A2/A1/c1 ));
 AND2_X1 \V2/V4/A2/A1/M2/M1/_0_  (.A1(\V2/V4/s1 [1]),
    .A2(\V2/V4/v1 [5]),
    .ZN(\V2/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M2/M1/_1_  (.A(\V2/V4/s1 [1]),
    .B(\V2/V4/v1 [5]),
    .Z(\V2/V4/A2/A1/M2/s1 ));
 AND2_X1 \V2/V4/A2/A1/M2/M2/_0_  (.A1(\V2/V4/A2/A1/M2/s1 ),
    .A2(\V2/V4/A2/A1/c1 ),
    .ZN(\V2/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M2/M2/_1_  (.A(\V2/V4/A2/A1/M2/s1 ),
    .B(\V2/V4/A2/A1/c1 ),
    .Z(\V2/v4 [5]));
 OR2_X1 \V2/V4/A2/A1/M2/_0_  (.A1(\V2/V4/A2/A1/M2/c1 ),
    .A2(\V2/V4/A2/A1/M2/c2 ),
    .ZN(\V2/V4/A2/A1/c2 ));
 AND2_X1 \V2/V4/A2/A1/M3/M1/_0_  (.A1(\V2/V4/s1 [2]),
    .A2(\V2/V4/v1 [6]),
    .ZN(\V2/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M3/M1/_1_  (.A(\V2/V4/s1 [2]),
    .B(\V2/V4/v1 [6]),
    .Z(\V2/V4/A2/A1/M3/s1 ));
 AND2_X1 \V2/V4/A2/A1/M3/M2/_0_  (.A1(\V2/V4/A2/A1/M3/s1 ),
    .A2(\V2/V4/A2/A1/c2 ),
    .ZN(\V2/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M3/M2/_1_  (.A(\V2/V4/A2/A1/M3/s1 ),
    .B(\V2/V4/A2/A1/c2 ),
    .Z(\V2/v4 [6]));
 OR2_X1 \V2/V4/A2/A1/M3/_0_  (.A1(\V2/V4/A2/A1/M3/c1 ),
    .A2(\V2/V4/A2/A1/M3/c2 ),
    .ZN(\V2/V4/A2/A1/c3 ));
 AND2_X1 \V2/V4/A2/A1/M4/M1/_0_  (.A1(\V2/V4/s1 [3]),
    .A2(\V2/V4/v1 [7]),
    .ZN(\V2/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M4/M1/_1_  (.A(\V2/V4/s1 [3]),
    .B(\V2/V4/v1 [7]),
    .Z(\V2/V4/A2/A1/M4/s1 ));
 AND2_X1 \V2/V4/A2/A1/M4/M2/_0_  (.A1(\V2/V4/A2/A1/M4/s1 ),
    .A2(\V2/V4/A2/A1/c3 ),
    .ZN(\V2/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M4/M2/_1_  (.A(\V2/V4/A2/A1/M4/s1 ),
    .B(\V2/V4/A2/A1/c3 ),
    .Z(\V2/v4 [7]));
 OR2_X1 \V2/V4/A2/A1/M4/_0_  (.A1(\V2/V4/A2/A1/M4/c1 ),
    .A2(\V2/V4/A2/A1/M4/c2 ),
    .ZN(\V2/V4/A2/c1 ));
 AND2_X1 \V2/V4/A2/A2/M1/M1/_0_  (.A1(\V2/V4/s1 [4]),
    .A2(ground),
    .ZN(\V2/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M1/M1/_1_  (.A(\V2/V4/s1 [4]),
    .B(ground),
    .Z(\V2/V4/A2/A2/M1/s1 ));
 AND2_X1 \V2/V4/A2/A2/M1/M2/_0_  (.A1(\V2/V4/A2/A2/M1/s1 ),
    .A2(\V2/V4/A2/c1 ),
    .ZN(\V2/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M1/M2/_1_  (.A(\V2/V4/A2/A2/M1/s1 ),
    .B(\V2/V4/A2/c1 ),
    .Z(\V2/V4/s2 [4]));
 OR2_X1 \V2/V4/A2/A2/M1/_0_  (.A1(\V2/V4/A2/A2/M1/c1 ),
    .A2(\V2/V4/A2/A2/M1/c2 ),
    .ZN(\V2/V4/A2/A2/c1 ));
 AND2_X1 \V2/V4/A2/A2/M2/M1/_0_  (.A1(\V2/V4/s1 [5]),
    .A2(ground),
    .ZN(\V2/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M2/M1/_1_  (.A(\V2/V4/s1 [5]),
    .B(ground),
    .Z(\V2/V4/A2/A2/M2/s1 ));
 AND2_X1 \V2/V4/A2/A2/M2/M2/_0_  (.A1(\V2/V4/A2/A2/M2/s1 ),
    .A2(\V2/V4/A2/A2/c1 ),
    .ZN(\V2/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M2/M2/_1_  (.A(\V2/V4/A2/A2/M2/s1 ),
    .B(\V2/V4/A2/A2/c1 ),
    .Z(\V2/V4/s2 [5]));
 OR2_X1 \V2/V4/A2/A2/M2/_0_  (.A1(\V2/V4/A2/A2/M2/c1 ),
    .A2(\V2/V4/A2/A2/M2/c2 ),
    .ZN(\V2/V4/A2/A2/c2 ));
 AND2_X1 \V2/V4/A2/A2/M3/M1/_0_  (.A1(\V2/V4/s1 [6]),
    .A2(ground),
    .ZN(\V2/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M3/M1/_1_  (.A(\V2/V4/s1 [6]),
    .B(ground),
    .Z(\V2/V4/A2/A2/M3/s1 ));
 AND2_X1 \V2/V4/A2/A2/M3/M2/_0_  (.A1(\V2/V4/A2/A2/M3/s1 ),
    .A2(\V2/V4/A2/A2/c2 ),
    .ZN(\V2/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M3/M2/_1_  (.A(\V2/V4/A2/A2/M3/s1 ),
    .B(\V2/V4/A2/A2/c2 ),
    .Z(\V2/V4/s2 [6]));
 OR2_X1 \V2/V4/A2/A2/M3/_0_  (.A1(\V2/V4/A2/A2/M3/c1 ),
    .A2(\V2/V4/A2/A2/M3/c2 ),
    .ZN(\V2/V4/A2/A2/c3 ));
 AND2_X1 \V2/V4/A2/A2/M4/M1/_0_  (.A1(\V2/V4/s1 [7]),
    .A2(ground),
    .ZN(\V2/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M4/M1/_1_  (.A(\V2/V4/s1 [7]),
    .B(ground),
    .Z(\V2/V4/A2/A2/M4/s1 ));
 AND2_X1 \V2/V4/A2/A2/M4/M2/_0_  (.A1(\V2/V4/A2/A2/M4/s1 ),
    .A2(\V2/V4/A2/A2/c3 ),
    .ZN(\V2/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M4/M2/_1_  (.A(\V2/V4/A2/A2/M4/s1 ),
    .B(\V2/V4/A2/A2/c3 ),
    .Z(\V2/V4/s2 [7]));
 OR2_X1 \V2/V4/A2/A2/M4/_0_  (.A1(\V2/V4/A2/A2/M4/c1 ),
    .A2(\V2/V4/A2/A2/M4/c2 ),
    .ZN(\V2/V4/c2 ));
 AND2_X1 \V2/V4/A3/A1/M1/M1/_0_  (.A1(\V2/V4/v4 [0]),
    .A2(\V2/V4/s2 [4]),
    .ZN(\V2/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M1/M1/_1_  (.A(\V2/V4/v4 [0]),
    .B(\V2/V4/s2 [4]),
    .Z(\V2/V4/A3/A1/M1/s1 ));
 AND2_X1 \V2/V4/A3/A1/M1/M2/_0_  (.A1(\V2/V4/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M1/M2/_1_  (.A(\V2/V4/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/v4 [8]));
 OR2_X1 \V2/V4/A3/A1/M1/_0_  (.A1(\V2/V4/A3/A1/M1/c1 ),
    .A2(\V2/V4/A3/A1/M1/c2 ),
    .ZN(\V2/V4/A3/A1/c1 ));
 AND2_X1 \V2/V4/A3/A1/M2/M1/_0_  (.A1(\V2/V4/v4 [1]),
    .A2(\V2/V4/s2 [5]),
    .ZN(\V2/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M2/M1/_1_  (.A(\V2/V4/v4 [1]),
    .B(\V2/V4/s2 [5]),
    .Z(\V2/V4/A3/A1/M2/s1 ));
 AND2_X1 \V2/V4/A3/A1/M2/M2/_0_  (.A1(\V2/V4/A3/A1/M2/s1 ),
    .A2(\V2/V4/A3/A1/c1 ),
    .ZN(\V2/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M2/M2/_1_  (.A(\V2/V4/A3/A1/M2/s1 ),
    .B(\V2/V4/A3/A1/c1 ),
    .Z(\V2/v4 [9]));
 OR2_X1 \V2/V4/A3/A1/M2/_0_  (.A1(\V2/V4/A3/A1/M2/c1 ),
    .A2(\V2/V4/A3/A1/M2/c2 ),
    .ZN(\V2/V4/A3/A1/c2 ));
 AND2_X1 \V2/V4/A3/A1/M3/M1/_0_  (.A1(\V2/V4/v4 [2]),
    .A2(\V2/V4/s2 [6]),
    .ZN(\V2/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M3/M1/_1_  (.A(\V2/V4/v4 [2]),
    .B(\V2/V4/s2 [6]),
    .Z(\V2/V4/A3/A1/M3/s1 ));
 AND2_X1 \V2/V4/A3/A1/M3/M2/_0_  (.A1(\V2/V4/A3/A1/M3/s1 ),
    .A2(\V2/V4/A3/A1/c2 ),
    .ZN(\V2/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M3/M2/_1_  (.A(\V2/V4/A3/A1/M3/s1 ),
    .B(\V2/V4/A3/A1/c2 ),
    .Z(\V2/v4 [10]));
 OR2_X1 \V2/V4/A3/A1/M3/_0_  (.A1(\V2/V4/A3/A1/M3/c1 ),
    .A2(\V2/V4/A3/A1/M3/c2 ),
    .ZN(\V2/V4/A3/A1/c3 ));
 AND2_X1 \V2/V4/A3/A1/M4/M1/_0_  (.A1(\V2/V4/v4 [3]),
    .A2(\V2/V4/s2 [7]),
    .ZN(\V2/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M4/M1/_1_  (.A(\V2/V4/v4 [3]),
    .B(\V2/V4/s2 [7]),
    .Z(\V2/V4/A3/A1/M4/s1 ));
 AND2_X1 \V2/V4/A3/A1/M4/M2/_0_  (.A1(\V2/V4/A3/A1/M4/s1 ),
    .A2(\V2/V4/A3/A1/c3 ),
    .ZN(\V2/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M4/M2/_1_  (.A(\V2/V4/A3/A1/M4/s1 ),
    .B(\V2/V4/A3/A1/c3 ),
    .Z(\V2/v4 [11]));
 OR2_X1 \V2/V4/A3/A1/M4/_0_  (.A1(\V2/V4/A3/A1/M4/c1 ),
    .A2(\V2/V4/A3/A1/M4/c2 ),
    .ZN(\V2/V4/A3/c1 ));
 AND2_X1 \V2/V4/A3/A2/M1/M1/_0_  (.A1(\V2/V4/v4 [4]),
    .A2(\V2/V4/c3 ),
    .ZN(\V2/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M1/M1/_1_  (.A(\V2/V4/v4 [4]),
    .B(\V2/V4/c3 ),
    .Z(\V2/V4/A3/A2/M1/s1 ));
 AND2_X1 \V2/V4/A3/A2/M1/M2/_0_  (.A1(\V2/V4/A3/A2/M1/s1 ),
    .A2(\V2/V4/A3/c1 ),
    .ZN(\V2/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M1/M2/_1_  (.A(\V2/V4/A3/A2/M1/s1 ),
    .B(\V2/V4/A3/c1 ),
    .Z(\V2/v4 [12]));
 OR2_X1 \V2/V4/A3/A2/M1/_0_  (.A1(\V2/V4/A3/A2/M1/c1 ),
    .A2(\V2/V4/A3/A2/M1/c2 ),
    .ZN(\V2/V4/A3/A2/c1 ));
 AND2_X1 \V2/V4/A3/A2/M2/M1/_0_  (.A1(\V2/V4/v4 [5]),
    .A2(ground),
    .ZN(\V2/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M2/M1/_1_  (.A(\V2/V4/v4 [5]),
    .B(ground),
    .Z(\V2/V4/A3/A2/M2/s1 ));
 AND2_X1 \V2/V4/A3/A2/M2/M2/_0_  (.A1(\V2/V4/A3/A2/M2/s1 ),
    .A2(\V2/V4/A3/A2/c1 ),
    .ZN(\V2/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M2/M2/_1_  (.A(\V2/V4/A3/A2/M2/s1 ),
    .B(\V2/V4/A3/A2/c1 ),
    .Z(\V2/v4 [13]));
 OR2_X1 \V2/V4/A3/A2/M2/_0_  (.A1(\V2/V4/A3/A2/M2/c1 ),
    .A2(\V2/V4/A3/A2/M2/c2 ),
    .ZN(\V2/V4/A3/A2/c2 ));
 AND2_X1 \V2/V4/A3/A2/M3/M1/_0_  (.A1(\V2/V4/v4 [6]),
    .A2(ground),
    .ZN(\V2/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M3/M1/_1_  (.A(\V2/V4/v4 [6]),
    .B(ground),
    .Z(\V2/V4/A3/A2/M3/s1 ));
 AND2_X1 \V2/V4/A3/A2/M3/M2/_0_  (.A1(\V2/V4/A3/A2/M3/s1 ),
    .A2(\V2/V4/A3/A2/c2 ),
    .ZN(\V2/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M3/M2/_1_  (.A(\V2/V4/A3/A2/M3/s1 ),
    .B(\V2/V4/A3/A2/c2 ),
    .Z(\V2/v4 [14]));
 OR2_X1 \V2/V4/A3/A2/M3/_0_  (.A1(\V2/V4/A3/A2/M3/c1 ),
    .A2(\V2/V4/A3/A2/M3/c2 ),
    .ZN(\V2/V4/A3/A2/c3 ));
 AND2_X1 \V2/V4/A3/A2/M4/M1/_0_  (.A1(\V2/V4/v4 [7]),
    .A2(ground),
    .ZN(\V2/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M4/M1/_1_  (.A(\V2/V4/v4 [7]),
    .B(ground),
    .Z(\V2/V4/A3/A2/M4/s1 ));
 AND2_X1 \V2/V4/A3/A2/M4/M2/_0_  (.A1(\V2/V4/A3/A2/M4/s1 ),
    .A2(\V2/V4/A3/A2/c3 ),
    .ZN(\V2/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M4/M2/_1_  (.A(\V2/V4/A3/A2/M4/s1 ),
    .B(\V2/V4/A3/A2/c3 ),
    .Z(\V2/v4 [15]));
 OR2_X1 \V2/V4/A3/A2/M4/_0_  (.A1(\V2/V4/A3/A2/M4/c1 ),
    .A2(\V2/V4/A3/A2/M4/c2 ),
    .ZN(\V2/V4/overflow ));
 AND2_X1 \V2/V4/V1/A1/M1/M1/_0_  (.A1(\V2/V4/V1/v2 [0]),
    .A2(\V2/V4/V1/v3 [0]),
    .ZN(\V2/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M1/M1/_1_  (.A(\V2/V4/V1/v2 [0]),
    .B(\V2/V4/V1/v3 [0]),
    .Z(\V2/V4/V1/A1/M1/s1 ));
 AND2_X1 \V2/V4/V1/A1/M1/M2/_0_  (.A1(\V2/V4/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M1/M2/_1_  (.A(\V2/V4/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/V1/s1 [0]));
 OR2_X1 \V2/V4/V1/A1/M1/_0_  (.A1(\V2/V4/V1/A1/M1/c1 ),
    .A2(\V2/V4/V1/A1/M1/c2 ),
    .ZN(\V2/V4/V1/A1/c1 ));
 AND2_X1 \V2/V4/V1/A1/M2/M1/_0_  (.A1(\V2/V4/V1/v2 [1]),
    .A2(\V2/V4/V1/v3 [1]),
    .ZN(\V2/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M2/M1/_1_  (.A(\V2/V4/V1/v2 [1]),
    .B(\V2/V4/V1/v3 [1]),
    .Z(\V2/V4/V1/A1/M2/s1 ));
 AND2_X1 \V2/V4/V1/A1/M2/M2/_0_  (.A1(\V2/V4/V1/A1/M2/s1 ),
    .A2(\V2/V4/V1/A1/c1 ),
    .ZN(\V2/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M2/M2/_1_  (.A(\V2/V4/V1/A1/M2/s1 ),
    .B(\V2/V4/V1/A1/c1 ),
    .Z(\V2/V4/V1/s1 [1]));
 OR2_X1 \V2/V4/V1/A1/M2/_0_  (.A1(\V2/V4/V1/A1/M2/c1 ),
    .A2(\V2/V4/V1/A1/M2/c2 ),
    .ZN(\V2/V4/V1/A1/c2 ));
 AND2_X1 \V2/V4/V1/A1/M3/M1/_0_  (.A1(\V2/V4/V1/v2 [2]),
    .A2(\V2/V4/V1/v3 [2]),
    .ZN(\V2/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M3/M1/_1_  (.A(\V2/V4/V1/v2 [2]),
    .B(\V2/V4/V1/v3 [2]),
    .Z(\V2/V4/V1/A1/M3/s1 ));
 AND2_X1 \V2/V4/V1/A1/M3/M2/_0_  (.A1(\V2/V4/V1/A1/M3/s1 ),
    .A2(\V2/V4/V1/A1/c2 ),
    .ZN(\V2/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M3/M2/_1_  (.A(\V2/V4/V1/A1/M3/s1 ),
    .B(\V2/V4/V1/A1/c2 ),
    .Z(\V2/V4/V1/s1 [2]));
 OR2_X1 \V2/V4/V1/A1/M3/_0_  (.A1(\V2/V4/V1/A1/M3/c1 ),
    .A2(\V2/V4/V1/A1/M3/c2 ),
    .ZN(\V2/V4/V1/A1/c3 ));
 AND2_X1 \V2/V4/V1/A1/M4/M1/_0_  (.A1(\V2/V4/V1/v2 [3]),
    .A2(\V2/V4/V1/v3 [3]),
    .ZN(\V2/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M4/M1/_1_  (.A(\V2/V4/V1/v2 [3]),
    .B(\V2/V4/V1/v3 [3]),
    .Z(\V2/V4/V1/A1/M4/s1 ));
 AND2_X1 \V2/V4/V1/A1/M4/M2/_0_  (.A1(\V2/V4/V1/A1/M4/s1 ),
    .A2(\V2/V4/V1/A1/c3 ),
    .ZN(\V2/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M4/M2/_1_  (.A(\V2/V4/V1/A1/M4/s1 ),
    .B(\V2/V4/V1/A1/c3 ),
    .Z(\V2/V4/V1/s1 [3]));
 OR2_X1 \V2/V4/V1/A1/M4/_0_  (.A1(\V2/V4/V1/A1/M4/c1 ),
    .A2(\V2/V4/V1/A1/M4/c2 ),
    .ZN(\V2/V4/V1/c1 ));
 AND2_X1 \V2/V4/V1/A2/M1/M1/_0_  (.A1(\V2/V4/V1/s1 [0]),
    .A2(\V2/V4/V1/v1 [2]),
    .ZN(\V2/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M1/M1/_1_  (.A(\V2/V4/V1/s1 [0]),
    .B(\V2/V4/V1/v1 [2]),
    .Z(\V2/V4/V1/A2/M1/s1 ));
 AND2_X1 \V2/V4/V1/A2/M1/M2/_0_  (.A1(\V2/V4/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M1/M2/_1_  (.A(\V2/V4/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/v4 [2]));
 OR2_X1 \V2/V4/V1/A2/M1/_0_  (.A1(\V2/V4/V1/A2/M1/c1 ),
    .A2(\V2/V4/V1/A2/M1/c2 ),
    .ZN(\V2/V4/V1/A2/c1 ));
 AND2_X1 \V2/V4/V1/A2/M2/M1/_0_  (.A1(\V2/V4/V1/s1 [1]),
    .A2(\V2/V4/V1/v1 [3]),
    .ZN(\V2/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M2/M1/_1_  (.A(\V2/V4/V1/s1 [1]),
    .B(\V2/V4/V1/v1 [3]),
    .Z(\V2/V4/V1/A2/M2/s1 ));
 AND2_X1 \V2/V4/V1/A2/M2/M2/_0_  (.A1(\V2/V4/V1/A2/M2/s1 ),
    .A2(\V2/V4/V1/A2/c1 ),
    .ZN(\V2/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M2/M2/_1_  (.A(\V2/V4/V1/A2/M2/s1 ),
    .B(\V2/V4/V1/A2/c1 ),
    .Z(\V2/v4 [3]));
 OR2_X1 \V2/V4/V1/A2/M2/_0_  (.A1(\V2/V4/V1/A2/M2/c1 ),
    .A2(\V2/V4/V1/A2/M2/c2 ),
    .ZN(\V2/V4/V1/A2/c2 ));
 AND2_X1 \V2/V4/V1/A2/M3/M1/_0_  (.A1(\V2/V4/V1/s1 [2]),
    .A2(ground),
    .ZN(\V2/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M3/M1/_1_  (.A(\V2/V4/V1/s1 [2]),
    .B(ground),
    .Z(\V2/V4/V1/A2/M3/s1 ));
 AND2_X1 \V2/V4/V1/A2/M3/M2/_0_  (.A1(\V2/V4/V1/A2/M3/s1 ),
    .A2(\V2/V4/V1/A2/c2 ),
    .ZN(\V2/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M3/M2/_1_  (.A(\V2/V4/V1/A2/M3/s1 ),
    .B(\V2/V4/V1/A2/c2 ),
    .Z(\V2/V4/V1/s2 [2]));
 OR2_X1 \V2/V4/V1/A2/M3/_0_  (.A1(\V2/V4/V1/A2/M3/c1 ),
    .A2(\V2/V4/V1/A2/M3/c2 ),
    .ZN(\V2/V4/V1/A2/c3 ));
 AND2_X1 \V2/V4/V1/A2/M4/M1/_0_  (.A1(\V2/V4/V1/s1 [3]),
    .A2(ground),
    .ZN(\V2/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M4/M1/_1_  (.A(\V2/V4/V1/s1 [3]),
    .B(ground),
    .Z(\V2/V4/V1/A2/M4/s1 ));
 AND2_X1 \V2/V4/V1/A2/M4/M2/_0_  (.A1(\V2/V4/V1/A2/M4/s1 ),
    .A2(\V2/V4/V1/A2/c3 ),
    .ZN(\V2/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M4/M2/_1_  (.A(\V2/V4/V1/A2/M4/s1 ),
    .B(\V2/V4/V1/A2/c3 ),
    .Z(\V2/V4/V1/s2 [3]));
 OR2_X1 \V2/V4/V1/A2/M4/_0_  (.A1(\V2/V4/V1/A2/M4/c1 ),
    .A2(\V2/V4/V1/A2/M4/c2 ),
    .ZN(\V2/V4/V1/c2 ));
 AND2_X1 \V2/V4/V1/A3/M1/M1/_0_  (.A1(\V2/V4/V1/v4 [0]),
    .A2(\V2/V4/V1/s2 [2]),
    .ZN(\V2/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M1/M1/_1_  (.A(\V2/V4/V1/v4 [0]),
    .B(\V2/V4/V1/s2 [2]),
    .Z(\V2/V4/V1/A3/M1/s1 ));
 AND2_X1 \V2/V4/V1/A3/M1/M2/_0_  (.A1(\V2/V4/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M1/M2/_1_  (.A(\V2/V4/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v1 [4]));
 OR2_X1 \V2/V4/V1/A3/M1/_0_  (.A1(\V2/V4/V1/A3/M1/c1 ),
    .A2(\V2/V4/V1/A3/M1/c2 ),
    .ZN(\V2/V4/V1/A3/c1 ));
 AND2_X1 \V2/V4/V1/A3/M2/M1/_0_  (.A1(\V2/V4/V1/v4 [1]),
    .A2(\V2/V4/V1/s2 [3]),
    .ZN(\V2/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M2/M1/_1_  (.A(\V2/V4/V1/v4 [1]),
    .B(\V2/V4/V1/s2 [3]),
    .Z(\V2/V4/V1/A3/M2/s1 ));
 AND2_X1 \V2/V4/V1/A3/M2/M2/_0_  (.A1(\V2/V4/V1/A3/M2/s1 ),
    .A2(\V2/V4/V1/A3/c1 ),
    .ZN(\V2/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M2/M2/_1_  (.A(\V2/V4/V1/A3/M2/s1 ),
    .B(\V2/V4/V1/A3/c1 ),
    .Z(\V2/V4/v1 [5]));
 OR2_X1 \V2/V4/V1/A3/M2/_0_  (.A1(\V2/V4/V1/A3/M2/c1 ),
    .A2(\V2/V4/V1/A3/M2/c2 ),
    .ZN(\V2/V4/V1/A3/c2 ));
 AND2_X1 \V2/V4/V1/A3/M3/M1/_0_  (.A1(\V2/V4/V1/v4 [2]),
    .A2(\V2/V4/V1/c3 ),
    .ZN(\V2/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M3/M1/_1_  (.A(\V2/V4/V1/v4 [2]),
    .B(\V2/V4/V1/c3 ),
    .Z(\V2/V4/V1/A3/M3/s1 ));
 AND2_X1 \V2/V4/V1/A3/M3/M2/_0_  (.A1(\V2/V4/V1/A3/M3/s1 ),
    .A2(\V2/V4/V1/A3/c2 ),
    .ZN(\V2/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M3/M2/_1_  (.A(\V2/V4/V1/A3/M3/s1 ),
    .B(\V2/V4/V1/A3/c2 ),
    .Z(\V2/V4/v1 [6]));
 OR2_X1 \V2/V4/V1/A3/M3/_0_  (.A1(\V2/V4/V1/A3/M3/c1 ),
    .A2(\V2/V4/V1/A3/M3/c2 ),
    .ZN(\V2/V4/V1/A3/c3 ));
 AND2_X1 \V2/V4/V1/A3/M4/M1/_0_  (.A1(\V2/V4/V1/v4 [3]),
    .A2(ground),
    .ZN(\V2/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M4/M1/_1_  (.A(\V2/V4/V1/v4 [3]),
    .B(ground),
    .Z(\V2/V4/V1/A3/M4/s1 ));
 AND2_X1 \V2/V4/V1/A3/M4/M2/_0_  (.A1(\V2/V4/V1/A3/M4/s1 ),
    .A2(\V2/V4/V1/A3/c3 ),
    .ZN(\V2/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M4/M2/_1_  (.A(\V2/V4/V1/A3/M4/s1 ),
    .B(\V2/V4/V1/A3/c3 ),
    .Z(\V2/V4/v1 [7]));
 OR2_X1 \V2/V4/V1/A3/M4/_0_  (.A1(\V2/V4/V1/A3/M4/c1 ),
    .A2(\V2/V4/V1/A3/M4/c2 ),
    .ZN(\V2/V4/V1/overflow ));
 AND2_X1 \V2/V4/V1/V1/HA1/_0_  (.A1(\V2/V4/V1/V1/w2 ),
    .A2(\V2/V4/V1/V1/w1 ),
    .ZN(\V2/V4/V1/V1/w4 ));
 XOR2_X2 \V2/V4/V1/V1/HA1/_1_  (.A(\V2/V4/V1/V1/w2 ),
    .B(\V2/V4/V1/V1/w1 ),
    .Z(\V2/v4 [1]));
 AND2_X1 \V2/V4/V1/V1/HA2/_0_  (.A1(\V2/V4/V1/V1/w4 ),
    .A2(\V2/V4/V1/V1/w3 ),
    .ZN(\V2/V4/V1/v1 [3]));
 XOR2_X2 \V2/V4/V1/V1/HA2/_1_  (.A(\V2/V4/V1/V1/w4 ),
    .B(\V2/V4/V1/V1/w3 ),
    .Z(\V2/V4/V1/v1 [2]));
 AND2_X1 \V2/V4/V1/V1/_0_  (.A1(A[24]),
    .A2(B[8]),
    .ZN(\V2/v4 [0]));
 AND2_X1 \V2/V4/V1/V1/_1_  (.A1(A[24]),
    .A2(B[9]),
    .ZN(\V2/V4/V1/V1/w1 ));
 AND2_X1 \V2/V4/V1/V1/_2_  (.A1(B[8]),
    .A2(A[25]),
    .ZN(\V2/V4/V1/V1/w2 ));
 AND2_X1 \V2/V4/V1/V1/_3_  (.A1(B[9]),
    .A2(A[25]),
    .ZN(\V2/V4/V1/V1/w3 ));
 AND2_X1 \V2/V4/V1/V2/HA1/_0_  (.A1(\V2/V4/V1/V2/w2 ),
    .A2(\V2/V4/V1/V2/w1 ),
    .ZN(\V2/V4/V1/V2/w4 ));
 XOR2_X2 \V2/V4/V1/V2/HA1/_1_  (.A(\V2/V4/V1/V2/w2 ),
    .B(\V2/V4/V1/V2/w1 ),
    .Z(\V2/V4/V1/v2 [1]));
 AND2_X1 \V2/V4/V1/V2/HA2/_0_  (.A1(\V2/V4/V1/V2/w4 ),
    .A2(\V2/V4/V1/V2/w3 ),
    .ZN(\V2/V4/V1/v2 [3]));
 XOR2_X2 \V2/V4/V1/V2/HA2/_1_  (.A(\V2/V4/V1/V2/w4 ),
    .B(\V2/V4/V1/V2/w3 ),
    .Z(\V2/V4/V1/v2 [2]));
 AND2_X1 \V2/V4/V1/V2/_0_  (.A1(A[26]),
    .A2(B[8]),
    .ZN(\V2/V4/V1/v2 [0]));
 AND2_X1 \V2/V4/V1/V2/_1_  (.A1(A[26]),
    .A2(B[9]),
    .ZN(\V2/V4/V1/V2/w1 ));
 AND2_X1 \V2/V4/V1/V2/_2_  (.A1(B[8]),
    .A2(A[27]),
    .ZN(\V2/V4/V1/V2/w2 ));
 AND2_X1 \V2/V4/V1/V2/_3_  (.A1(B[9]),
    .A2(A[27]),
    .ZN(\V2/V4/V1/V2/w3 ));
 AND2_X1 \V2/V4/V1/V3/HA1/_0_  (.A1(\V2/V4/V1/V3/w2 ),
    .A2(\V2/V4/V1/V3/w1 ),
    .ZN(\V2/V4/V1/V3/w4 ));
 XOR2_X2 \V2/V4/V1/V3/HA1/_1_  (.A(\V2/V4/V1/V3/w2 ),
    .B(\V2/V4/V1/V3/w1 ),
    .Z(\V2/V4/V1/v3 [1]));
 AND2_X1 \V2/V4/V1/V3/HA2/_0_  (.A1(\V2/V4/V1/V3/w4 ),
    .A2(\V2/V4/V1/V3/w3 ),
    .ZN(\V2/V4/V1/v3 [3]));
 XOR2_X2 \V2/V4/V1/V3/HA2/_1_  (.A(\V2/V4/V1/V3/w4 ),
    .B(\V2/V4/V1/V3/w3 ),
    .Z(\V2/V4/V1/v3 [2]));
 AND2_X1 \V2/V4/V1/V3/_0_  (.A1(A[24]),
    .A2(B[10]),
    .ZN(\V2/V4/V1/v3 [0]));
 AND2_X1 \V2/V4/V1/V3/_1_  (.A1(A[24]),
    .A2(B[11]),
    .ZN(\V2/V4/V1/V3/w1 ));
 AND2_X1 \V2/V4/V1/V3/_2_  (.A1(B[10]),
    .A2(A[25]),
    .ZN(\V2/V4/V1/V3/w2 ));
 AND2_X1 \V2/V4/V1/V3/_3_  (.A1(B[11]),
    .A2(A[25]),
    .ZN(\V2/V4/V1/V3/w3 ));
 AND2_X1 \V2/V4/V1/V4/HA1/_0_  (.A1(\V2/V4/V1/V4/w2 ),
    .A2(\V2/V4/V1/V4/w1 ),
    .ZN(\V2/V4/V1/V4/w4 ));
 XOR2_X2 \V2/V4/V1/V4/HA1/_1_  (.A(\V2/V4/V1/V4/w2 ),
    .B(\V2/V4/V1/V4/w1 ),
    .Z(\V2/V4/V1/v4 [1]));
 AND2_X1 \V2/V4/V1/V4/HA2/_0_  (.A1(\V2/V4/V1/V4/w4 ),
    .A2(\V2/V4/V1/V4/w3 ),
    .ZN(\V2/V4/V1/v4 [3]));
 XOR2_X2 \V2/V4/V1/V4/HA2/_1_  (.A(\V2/V4/V1/V4/w4 ),
    .B(\V2/V4/V1/V4/w3 ),
    .Z(\V2/V4/V1/v4 [2]));
 AND2_X1 \V2/V4/V1/V4/_0_  (.A1(A[26]),
    .A2(B[10]),
    .ZN(\V2/V4/V1/v4 [0]));
 AND2_X1 \V2/V4/V1/V4/_1_  (.A1(A[26]),
    .A2(B[11]),
    .ZN(\V2/V4/V1/V4/w1 ));
 AND2_X1 \V2/V4/V1/V4/_2_  (.A1(B[10]),
    .A2(A[27]),
    .ZN(\V2/V4/V1/V4/w2 ));
 AND2_X1 \V2/V4/V1/V4/_3_  (.A1(B[11]),
    .A2(A[27]),
    .ZN(\V2/V4/V1/V4/w3 ));
 OR2_X1 \V2/V4/V1/_0_  (.A1(\V2/V4/V1/c1 ),
    .A2(\V2/V4/V1/c2 ),
    .ZN(\V2/V4/V1/c3 ));
 AND2_X1 \V2/V4/V2/A1/M1/M1/_0_  (.A1(\V2/V4/V2/v2 [0]),
    .A2(\V2/V4/V2/v3 [0]),
    .ZN(\V2/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M1/M1/_1_  (.A(\V2/V4/V2/v2 [0]),
    .B(\V2/V4/V2/v3 [0]),
    .Z(\V2/V4/V2/A1/M1/s1 ));
 AND2_X1 \V2/V4/V2/A1/M1/M2/_0_  (.A1(\V2/V4/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M1/M2/_1_  (.A(\V2/V4/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/V2/s1 [0]));
 OR2_X1 \V2/V4/V2/A1/M1/_0_  (.A1(\V2/V4/V2/A1/M1/c1 ),
    .A2(\V2/V4/V2/A1/M1/c2 ),
    .ZN(\V2/V4/V2/A1/c1 ));
 AND2_X1 \V2/V4/V2/A1/M2/M1/_0_  (.A1(\V2/V4/V2/v2 [1]),
    .A2(\V2/V4/V2/v3 [1]),
    .ZN(\V2/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M2/M1/_1_  (.A(\V2/V4/V2/v2 [1]),
    .B(\V2/V4/V2/v3 [1]),
    .Z(\V2/V4/V2/A1/M2/s1 ));
 AND2_X1 \V2/V4/V2/A1/M2/M2/_0_  (.A1(\V2/V4/V2/A1/M2/s1 ),
    .A2(\V2/V4/V2/A1/c1 ),
    .ZN(\V2/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M2/M2/_1_  (.A(\V2/V4/V2/A1/M2/s1 ),
    .B(\V2/V4/V2/A1/c1 ),
    .Z(\V2/V4/V2/s1 [1]));
 OR2_X1 \V2/V4/V2/A1/M2/_0_  (.A1(\V2/V4/V2/A1/M2/c1 ),
    .A2(\V2/V4/V2/A1/M2/c2 ),
    .ZN(\V2/V4/V2/A1/c2 ));
 AND2_X1 \V2/V4/V2/A1/M3/M1/_0_  (.A1(\V2/V4/V2/v2 [2]),
    .A2(\V2/V4/V2/v3 [2]),
    .ZN(\V2/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M3/M1/_1_  (.A(\V2/V4/V2/v2 [2]),
    .B(\V2/V4/V2/v3 [2]),
    .Z(\V2/V4/V2/A1/M3/s1 ));
 AND2_X1 \V2/V4/V2/A1/M3/M2/_0_  (.A1(\V2/V4/V2/A1/M3/s1 ),
    .A2(\V2/V4/V2/A1/c2 ),
    .ZN(\V2/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M3/M2/_1_  (.A(\V2/V4/V2/A1/M3/s1 ),
    .B(\V2/V4/V2/A1/c2 ),
    .Z(\V2/V4/V2/s1 [2]));
 OR2_X1 \V2/V4/V2/A1/M3/_0_  (.A1(\V2/V4/V2/A1/M3/c1 ),
    .A2(\V2/V4/V2/A1/M3/c2 ),
    .ZN(\V2/V4/V2/A1/c3 ));
 AND2_X1 \V2/V4/V2/A1/M4/M1/_0_  (.A1(\V2/V4/V2/v2 [3]),
    .A2(\V2/V4/V2/v3 [3]),
    .ZN(\V2/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M4/M1/_1_  (.A(\V2/V4/V2/v2 [3]),
    .B(\V2/V4/V2/v3 [3]),
    .Z(\V2/V4/V2/A1/M4/s1 ));
 AND2_X1 \V2/V4/V2/A1/M4/M2/_0_  (.A1(\V2/V4/V2/A1/M4/s1 ),
    .A2(\V2/V4/V2/A1/c3 ),
    .ZN(\V2/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M4/M2/_1_  (.A(\V2/V4/V2/A1/M4/s1 ),
    .B(\V2/V4/V2/A1/c3 ),
    .Z(\V2/V4/V2/s1 [3]));
 OR2_X1 \V2/V4/V2/A1/M4/_0_  (.A1(\V2/V4/V2/A1/M4/c1 ),
    .A2(\V2/V4/V2/A1/M4/c2 ),
    .ZN(\V2/V4/V2/c1 ));
 AND2_X1 \V2/V4/V2/A2/M1/M1/_0_  (.A1(\V2/V4/V2/s1 [0]),
    .A2(\V2/V4/V2/v1 [2]),
    .ZN(\V2/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M1/M1/_1_  (.A(\V2/V4/V2/s1 [0]),
    .B(\V2/V4/V2/v1 [2]),
    .Z(\V2/V4/V2/A2/M1/s1 ));
 AND2_X1 \V2/V4/V2/A2/M1/M2/_0_  (.A1(\V2/V4/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M1/M2/_1_  (.A(\V2/V4/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v2 [2]));
 OR2_X1 \V2/V4/V2/A2/M1/_0_  (.A1(\V2/V4/V2/A2/M1/c1 ),
    .A2(\V2/V4/V2/A2/M1/c2 ),
    .ZN(\V2/V4/V2/A2/c1 ));
 AND2_X1 \V2/V4/V2/A2/M2/M1/_0_  (.A1(\V2/V4/V2/s1 [1]),
    .A2(\V2/V4/V2/v1 [3]),
    .ZN(\V2/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M2/M1/_1_  (.A(\V2/V4/V2/s1 [1]),
    .B(\V2/V4/V2/v1 [3]),
    .Z(\V2/V4/V2/A2/M2/s1 ));
 AND2_X1 \V2/V4/V2/A2/M2/M2/_0_  (.A1(\V2/V4/V2/A2/M2/s1 ),
    .A2(\V2/V4/V2/A2/c1 ),
    .ZN(\V2/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M2/M2/_1_  (.A(\V2/V4/V2/A2/M2/s1 ),
    .B(\V2/V4/V2/A2/c1 ),
    .Z(\V2/V4/v2 [3]));
 OR2_X1 \V2/V4/V2/A2/M2/_0_  (.A1(\V2/V4/V2/A2/M2/c1 ),
    .A2(\V2/V4/V2/A2/M2/c2 ),
    .ZN(\V2/V4/V2/A2/c2 ));
 AND2_X1 \V2/V4/V2/A2/M3/M1/_0_  (.A1(\V2/V4/V2/s1 [2]),
    .A2(ground),
    .ZN(\V2/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M3/M1/_1_  (.A(\V2/V4/V2/s1 [2]),
    .B(ground),
    .Z(\V2/V4/V2/A2/M3/s1 ));
 AND2_X1 \V2/V4/V2/A2/M3/M2/_0_  (.A1(\V2/V4/V2/A2/M3/s1 ),
    .A2(\V2/V4/V2/A2/c2 ),
    .ZN(\V2/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M3/M2/_1_  (.A(\V2/V4/V2/A2/M3/s1 ),
    .B(\V2/V4/V2/A2/c2 ),
    .Z(\V2/V4/V2/s2 [2]));
 OR2_X1 \V2/V4/V2/A2/M3/_0_  (.A1(\V2/V4/V2/A2/M3/c1 ),
    .A2(\V2/V4/V2/A2/M3/c2 ),
    .ZN(\V2/V4/V2/A2/c3 ));
 AND2_X1 \V2/V4/V2/A2/M4/M1/_0_  (.A1(\V2/V4/V2/s1 [3]),
    .A2(ground),
    .ZN(\V2/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M4/M1/_1_  (.A(\V2/V4/V2/s1 [3]),
    .B(ground),
    .Z(\V2/V4/V2/A2/M4/s1 ));
 AND2_X1 \V2/V4/V2/A2/M4/M2/_0_  (.A1(\V2/V4/V2/A2/M4/s1 ),
    .A2(\V2/V4/V2/A2/c3 ),
    .ZN(\V2/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M4/M2/_1_  (.A(\V2/V4/V2/A2/M4/s1 ),
    .B(\V2/V4/V2/A2/c3 ),
    .Z(\V2/V4/V2/s2 [3]));
 OR2_X1 \V2/V4/V2/A2/M4/_0_  (.A1(\V2/V4/V2/A2/M4/c1 ),
    .A2(\V2/V4/V2/A2/M4/c2 ),
    .ZN(\V2/V4/V2/c2 ));
 AND2_X1 \V2/V4/V2/A3/M1/M1/_0_  (.A1(\V2/V4/V2/v4 [0]),
    .A2(\V2/V4/V2/s2 [2]),
    .ZN(\V2/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M1/M1/_1_  (.A(\V2/V4/V2/v4 [0]),
    .B(\V2/V4/V2/s2 [2]),
    .Z(\V2/V4/V2/A3/M1/s1 ));
 AND2_X1 \V2/V4/V2/A3/M1/M2/_0_  (.A1(\V2/V4/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M1/M2/_1_  (.A(\V2/V4/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v2 [4]));
 OR2_X1 \V2/V4/V2/A3/M1/_0_  (.A1(\V2/V4/V2/A3/M1/c1 ),
    .A2(\V2/V4/V2/A3/M1/c2 ),
    .ZN(\V2/V4/V2/A3/c1 ));
 AND2_X1 \V2/V4/V2/A3/M2/M1/_0_  (.A1(\V2/V4/V2/v4 [1]),
    .A2(\V2/V4/V2/s2 [3]),
    .ZN(\V2/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M2/M1/_1_  (.A(\V2/V4/V2/v4 [1]),
    .B(\V2/V4/V2/s2 [3]),
    .Z(\V2/V4/V2/A3/M2/s1 ));
 AND2_X1 \V2/V4/V2/A3/M2/M2/_0_  (.A1(\V2/V4/V2/A3/M2/s1 ),
    .A2(\V2/V4/V2/A3/c1 ),
    .ZN(\V2/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M2/M2/_1_  (.A(\V2/V4/V2/A3/M2/s1 ),
    .B(\V2/V4/V2/A3/c1 ),
    .Z(\V2/V4/v2 [5]));
 OR2_X1 \V2/V4/V2/A3/M2/_0_  (.A1(\V2/V4/V2/A3/M2/c1 ),
    .A2(\V2/V4/V2/A3/M2/c2 ),
    .ZN(\V2/V4/V2/A3/c2 ));
 AND2_X1 \V2/V4/V2/A3/M3/M1/_0_  (.A1(\V2/V4/V2/v4 [2]),
    .A2(\V2/V4/V2/c3 ),
    .ZN(\V2/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M3/M1/_1_  (.A(\V2/V4/V2/v4 [2]),
    .B(\V2/V4/V2/c3 ),
    .Z(\V2/V4/V2/A3/M3/s1 ));
 AND2_X1 \V2/V4/V2/A3/M3/M2/_0_  (.A1(\V2/V4/V2/A3/M3/s1 ),
    .A2(\V2/V4/V2/A3/c2 ),
    .ZN(\V2/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M3/M2/_1_  (.A(\V2/V4/V2/A3/M3/s1 ),
    .B(\V2/V4/V2/A3/c2 ),
    .Z(\V2/V4/v2 [6]));
 OR2_X1 \V2/V4/V2/A3/M3/_0_  (.A1(\V2/V4/V2/A3/M3/c1 ),
    .A2(\V2/V4/V2/A3/M3/c2 ),
    .ZN(\V2/V4/V2/A3/c3 ));
 AND2_X1 \V2/V4/V2/A3/M4/M1/_0_  (.A1(\V2/V4/V2/v4 [3]),
    .A2(ground),
    .ZN(\V2/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M4/M1/_1_  (.A(\V2/V4/V2/v4 [3]),
    .B(ground),
    .Z(\V2/V4/V2/A3/M4/s1 ));
 AND2_X1 \V2/V4/V2/A3/M4/M2/_0_  (.A1(\V2/V4/V2/A3/M4/s1 ),
    .A2(\V2/V4/V2/A3/c3 ),
    .ZN(\V2/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M4/M2/_1_  (.A(\V2/V4/V2/A3/M4/s1 ),
    .B(\V2/V4/V2/A3/c3 ),
    .Z(\V2/V4/v2 [7]));
 OR2_X1 \V2/V4/V2/A3/M4/_0_  (.A1(\V2/V4/V2/A3/M4/c1 ),
    .A2(\V2/V4/V2/A3/M4/c2 ),
    .ZN(\V2/V4/V2/overflow ));
 AND2_X1 \V2/V4/V2/V1/HA1/_0_  (.A1(\V2/V4/V2/V1/w2 ),
    .A2(\V2/V4/V2/V1/w1 ),
    .ZN(\V2/V4/V2/V1/w4 ));
 XOR2_X2 \V2/V4/V2/V1/HA1/_1_  (.A(\V2/V4/V2/V1/w2 ),
    .B(\V2/V4/V2/V1/w1 ),
    .Z(\V2/V4/v2 [1]));
 AND2_X1 \V2/V4/V2/V1/HA2/_0_  (.A1(\V2/V4/V2/V1/w4 ),
    .A2(\V2/V4/V2/V1/w3 ),
    .ZN(\V2/V4/V2/v1 [3]));
 XOR2_X2 \V2/V4/V2/V1/HA2/_1_  (.A(\V2/V4/V2/V1/w4 ),
    .B(\V2/V4/V2/V1/w3 ),
    .Z(\V2/V4/V2/v1 [2]));
 AND2_X1 \V2/V4/V2/V1/_0_  (.A1(A[28]),
    .A2(B[8]),
    .ZN(\V2/V4/v2 [0]));
 AND2_X1 \V2/V4/V2/V1/_1_  (.A1(A[28]),
    .A2(B[9]),
    .ZN(\V2/V4/V2/V1/w1 ));
 AND2_X1 \V2/V4/V2/V1/_2_  (.A1(B[8]),
    .A2(A[29]),
    .ZN(\V2/V4/V2/V1/w2 ));
 AND2_X1 \V2/V4/V2/V1/_3_  (.A1(B[9]),
    .A2(A[29]),
    .ZN(\V2/V4/V2/V1/w3 ));
 AND2_X1 \V2/V4/V2/V2/HA1/_0_  (.A1(\V2/V4/V2/V2/w2 ),
    .A2(\V2/V4/V2/V2/w1 ),
    .ZN(\V2/V4/V2/V2/w4 ));
 XOR2_X2 \V2/V4/V2/V2/HA1/_1_  (.A(\V2/V4/V2/V2/w2 ),
    .B(\V2/V4/V2/V2/w1 ),
    .Z(\V2/V4/V2/v2 [1]));
 AND2_X1 \V2/V4/V2/V2/HA2/_0_  (.A1(\V2/V4/V2/V2/w4 ),
    .A2(\V2/V4/V2/V2/w3 ),
    .ZN(\V2/V4/V2/v2 [3]));
 XOR2_X2 \V2/V4/V2/V2/HA2/_1_  (.A(\V2/V4/V2/V2/w4 ),
    .B(\V2/V4/V2/V2/w3 ),
    .Z(\V2/V4/V2/v2 [2]));
 AND2_X1 \V2/V4/V2/V2/_0_  (.A1(A[30]),
    .A2(B[8]),
    .ZN(\V2/V4/V2/v2 [0]));
 AND2_X1 \V2/V4/V2/V2/_1_  (.A1(A[30]),
    .A2(B[9]),
    .ZN(\V2/V4/V2/V2/w1 ));
 AND2_X1 \V2/V4/V2/V2/_2_  (.A1(B[8]),
    .A2(A[31]),
    .ZN(\V2/V4/V2/V2/w2 ));
 AND2_X1 \V2/V4/V2/V2/_3_  (.A1(B[9]),
    .A2(A[31]),
    .ZN(\V2/V4/V2/V2/w3 ));
 AND2_X1 \V2/V4/V2/V3/HA1/_0_  (.A1(\V2/V4/V2/V3/w2 ),
    .A2(\V2/V4/V2/V3/w1 ),
    .ZN(\V2/V4/V2/V3/w4 ));
 XOR2_X2 \V2/V4/V2/V3/HA1/_1_  (.A(\V2/V4/V2/V3/w2 ),
    .B(\V2/V4/V2/V3/w1 ),
    .Z(\V2/V4/V2/v3 [1]));
 AND2_X1 \V2/V4/V2/V3/HA2/_0_  (.A1(\V2/V4/V2/V3/w4 ),
    .A2(\V2/V4/V2/V3/w3 ),
    .ZN(\V2/V4/V2/v3 [3]));
 XOR2_X2 \V2/V4/V2/V3/HA2/_1_  (.A(\V2/V4/V2/V3/w4 ),
    .B(\V2/V4/V2/V3/w3 ),
    .Z(\V2/V4/V2/v3 [2]));
 AND2_X1 \V2/V4/V2/V3/_0_  (.A1(A[28]),
    .A2(B[10]),
    .ZN(\V2/V4/V2/v3 [0]));
 AND2_X1 \V2/V4/V2/V3/_1_  (.A1(A[28]),
    .A2(B[11]),
    .ZN(\V2/V4/V2/V3/w1 ));
 AND2_X1 \V2/V4/V2/V3/_2_  (.A1(B[10]),
    .A2(A[29]),
    .ZN(\V2/V4/V2/V3/w2 ));
 AND2_X1 \V2/V4/V2/V3/_3_  (.A1(B[11]),
    .A2(A[29]),
    .ZN(\V2/V4/V2/V3/w3 ));
 AND2_X1 \V2/V4/V2/V4/HA1/_0_  (.A1(\V2/V4/V2/V4/w2 ),
    .A2(\V2/V4/V2/V4/w1 ),
    .ZN(\V2/V4/V2/V4/w4 ));
 XOR2_X2 \V2/V4/V2/V4/HA1/_1_  (.A(\V2/V4/V2/V4/w2 ),
    .B(\V2/V4/V2/V4/w1 ),
    .Z(\V2/V4/V2/v4 [1]));
 AND2_X1 \V2/V4/V2/V4/HA2/_0_  (.A1(\V2/V4/V2/V4/w4 ),
    .A2(\V2/V4/V2/V4/w3 ),
    .ZN(\V2/V4/V2/v4 [3]));
 XOR2_X2 \V2/V4/V2/V4/HA2/_1_  (.A(\V2/V4/V2/V4/w4 ),
    .B(\V2/V4/V2/V4/w3 ),
    .Z(\V2/V4/V2/v4 [2]));
 AND2_X1 \V2/V4/V2/V4/_0_  (.A1(A[30]),
    .A2(B[10]),
    .ZN(\V2/V4/V2/v4 [0]));
 AND2_X1 \V2/V4/V2/V4/_1_  (.A1(A[30]),
    .A2(B[11]),
    .ZN(\V2/V4/V2/V4/w1 ));
 AND2_X1 \V2/V4/V2/V4/_2_  (.A1(B[10]),
    .A2(A[31]),
    .ZN(\V2/V4/V2/V4/w2 ));
 AND2_X1 \V2/V4/V2/V4/_3_  (.A1(B[11]),
    .A2(A[31]),
    .ZN(\V2/V4/V2/V4/w3 ));
 OR2_X1 \V2/V4/V2/_0_  (.A1(\V2/V4/V2/c1 ),
    .A2(\V2/V4/V2/c2 ),
    .ZN(\V2/V4/V2/c3 ));
 AND2_X1 \V2/V4/V3/A1/M1/M1/_0_  (.A1(\V2/V4/V3/v2 [0]),
    .A2(\V2/V4/V3/v3 [0]),
    .ZN(\V2/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M1/M1/_1_  (.A(\V2/V4/V3/v2 [0]),
    .B(\V2/V4/V3/v3 [0]),
    .Z(\V2/V4/V3/A1/M1/s1 ));
 AND2_X1 \V2/V4/V3/A1/M1/M2/_0_  (.A1(\V2/V4/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M1/M2/_1_  (.A(\V2/V4/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/V3/s1 [0]));
 OR2_X1 \V2/V4/V3/A1/M1/_0_  (.A1(\V2/V4/V3/A1/M1/c1 ),
    .A2(\V2/V4/V3/A1/M1/c2 ),
    .ZN(\V2/V4/V3/A1/c1 ));
 AND2_X1 \V2/V4/V3/A1/M2/M1/_0_  (.A1(\V2/V4/V3/v2 [1]),
    .A2(\V2/V4/V3/v3 [1]),
    .ZN(\V2/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M2/M1/_1_  (.A(\V2/V4/V3/v2 [1]),
    .B(\V2/V4/V3/v3 [1]),
    .Z(\V2/V4/V3/A1/M2/s1 ));
 AND2_X1 \V2/V4/V3/A1/M2/M2/_0_  (.A1(\V2/V4/V3/A1/M2/s1 ),
    .A2(\V2/V4/V3/A1/c1 ),
    .ZN(\V2/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M2/M2/_1_  (.A(\V2/V4/V3/A1/M2/s1 ),
    .B(\V2/V4/V3/A1/c1 ),
    .Z(\V2/V4/V3/s1 [1]));
 OR2_X1 \V2/V4/V3/A1/M2/_0_  (.A1(\V2/V4/V3/A1/M2/c1 ),
    .A2(\V2/V4/V3/A1/M2/c2 ),
    .ZN(\V2/V4/V3/A1/c2 ));
 AND2_X1 \V2/V4/V3/A1/M3/M1/_0_  (.A1(\V2/V4/V3/v2 [2]),
    .A2(\V2/V4/V3/v3 [2]),
    .ZN(\V2/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M3/M1/_1_  (.A(\V2/V4/V3/v2 [2]),
    .B(\V2/V4/V3/v3 [2]),
    .Z(\V2/V4/V3/A1/M3/s1 ));
 AND2_X1 \V2/V4/V3/A1/M3/M2/_0_  (.A1(\V2/V4/V3/A1/M3/s1 ),
    .A2(\V2/V4/V3/A1/c2 ),
    .ZN(\V2/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M3/M2/_1_  (.A(\V2/V4/V3/A1/M3/s1 ),
    .B(\V2/V4/V3/A1/c2 ),
    .Z(\V2/V4/V3/s1 [2]));
 OR2_X1 \V2/V4/V3/A1/M3/_0_  (.A1(\V2/V4/V3/A1/M3/c1 ),
    .A2(\V2/V4/V3/A1/M3/c2 ),
    .ZN(\V2/V4/V3/A1/c3 ));
 AND2_X1 \V2/V4/V3/A1/M4/M1/_0_  (.A1(\V2/V4/V3/v2 [3]),
    .A2(\V2/V4/V3/v3 [3]),
    .ZN(\V2/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M4/M1/_1_  (.A(\V2/V4/V3/v2 [3]),
    .B(\V2/V4/V3/v3 [3]),
    .Z(\V2/V4/V3/A1/M4/s1 ));
 AND2_X1 \V2/V4/V3/A1/M4/M2/_0_  (.A1(\V2/V4/V3/A1/M4/s1 ),
    .A2(\V2/V4/V3/A1/c3 ),
    .ZN(\V2/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M4/M2/_1_  (.A(\V2/V4/V3/A1/M4/s1 ),
    .B(\V2/V4/V3/A1/c3 ),
    .Z(\V2/V4/V3/s1 [3]));
 OR2_X1 \V2/V4/V3/A1/M4/_0_  (.A1(\V2/V4/V3/A1/M4/c1 ),
    .A2(\V2/V4/V3/A1/M4/c2 ),
    .ZN(\V2/V4/V3/c1 ));
 AND2_X1 \V2/V4/V3/A2/M1/M1/_0_  (.A1(\V2/V4/V3/s1 [0]),
    .A2(\V2/V4/V3/v1 [2]),
    .ZN(\V2/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M1/M1/_1_  (.A(\V2/V4/V3/s1 [0]),
    .B(\V2/V4/V3/v1 [2]),
    .Z(\V2/V4/V3/A2/M1/s1 ));
 AND2_X1 \V2/V4/V3/A2/M1/M2/_0_  (.A1(\V2/V4/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M1/M2/_1_  (.A(\V2/V4/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v3 [2]));
 OR2_X1 \V2/V4/V3/A2/M1/_0_  (.A1(\V2/V4/V3/A2/M1/c1 ),
    .A2(\V2/V4/V3/A2/M1/c2 ),
    .ZN(\V2/V4/V3/A2/c1 ));
 AND2_X1 \V2/V4/V3/A2/M2/M1/_0_  (.A1(\V2/V4/V3/s1 [1]),
    .A2(\V2/V4/V3/v1 [3]),
    .ZN(\V2/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M2/M1/_1_  (.A(\V2/V4/V3/s1 [1]),
    .B(\V2/V4/V3/v1 [3]),
    .Z(\V2/V4/V3/A2/M2/s1 ));
 AND2_X1 \V2/V4/V3/A2/M2/M2/_0_  (.A1(\V2/V4/V3/A2/M2/s1 ),
    .A2(\V2/V4/V3/A2/c1 ),
    .ZN(\V2/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M2/M2/_1_  (.A(\V2/V4/V3/A2/M2/s1 ),
    .B(\V2/V4/V3/A2/c1 ),
    .Z(\V2/V4/v3 [3]));
 OR2_X1 \V2/V4/V3/A2/M2/_0_  (.A1(\V2/V4/V3/A2/M2/c1 ),
    .A2(\V2/V4/V3/A2/M2/c2 ),
    .ZN(\V2/V4/V3/A2/c2 ));
 AND2_X1 \V2/V4/V3/A2/M3/M1/_0_  (.A1(\V2/V4/V3/s1 [2]),
    .A2(ground),
    .ZN(\V2/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M3/M1/_1_  (.A(\V2/V4/V3/s1 [2]),
    .B(ground),
    .Z(\V2/V4/V3/A2/M3/s1 ));
 AND2_X1 \V2/V4/V3/A2/M3/M2/_0_  (.A1(\V2/V4/V3/A2/M3/s1 ),
    .A2(\V2/V4/V3/A2/c2 ),
    .ZN(\V2/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M3/M2/_1_  (.A(\V2/V4/V3/A2/M3/s1 ),
    .B(\V2/V4/V3/A2/c2 ),
    .Z(\V2/V4/V3/s2 [2]));
 OR2_X1 \V2/V4/V3/A2/M3/_0_  (.A1(\V2/V4/V3/A2/M3/c1 ),
    .A2(\V2/V4/V3/A2/M3/c2 ),
    .ZN(\V2/V4/V3/A2/c3 ));
 AND2_X1 \V2/V4/V3/A2/M4/M1/_0_  (.A1(\V2/V4/V3/s1 [3]),
    .A2(ground),
    .ZN(\V2/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M4/M1/_1_  (.A(\V2/V4/V3/s1 [3]),
    .B(ground),
    .Z(\V2/V4/V3/A2/M4/s1 ));
 AND2_X1 \V2/V4/V3/A2/M4/M2/_0_  (.A1(\V2/V4/V3/A2/M4/s1 ),
    .A2(\V2/V4/V3/A2/c3 ),
    .ZN(\V2/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M4/M2/_1_  (.A(\V2/V4/V3/A2/M4/s1 ),
    .B(\V2/V4/V3/A2/c3 ),
    .Z(\V2/V4/V3/s2 [3]));
 OR2_X1 \V2/V4/V3/A2/M4/_0_  (.A1(\V2/V4/V3/A2/M4/c1 ),
    .A2(\V2/V4/V3/A2/M4/c2 ),
    .ZN(\V2/V4/V3/c2 ));
 AND2_X1 \V2/V4/V3/A3/M1/M1/_0_  (.A1(\V2/V4/V3/v4 [0]),
    .A2(\V2/V4/V3/s2 [2]),
    .ZN(\V2/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M1/M1/_1_  (.A(\V2/V4/V3/v4 [0]),
    .B(\V2/V4/V3/s2 [2]),
    .Z(\V2/V4/V3/A3/M1/s1 ));
 AND2_X1 \V2/V4/V3/A3/M1/M2/_0_  (.A1(\V2/V4/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M1/M2/_1_  (.A(\V2/V4/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v3 [4]));
 OR2_X1 \V2/V4/V3/A3/M1/_0_  (.A1(\V2/V4/V3/A3/M1/c1 ),
    .A2(\V2/V4/V3/A3/M1/c2 ),
    .ZN(\V2/V4/V3/A3/c1 ));
 AND2_X1 \V2/V4/V3/A3/M2/M1/_0_  (.A1(\V2/V4/V3/v4 [1]),
    .A2(\V2/V4/V3/s2 [3]),
    .ZN(\V2/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M2/M1/_1_  (.A(\V2/V4/V3/v4 [1]),
    .B(\V2/V4/V3/s2 [3]),
    .Z(\V2/V4/V3/A3/M2/s1 ));
 AND2_X1 \V2/V4/V3/A3/M2/M2/_0_  (.A1(\V2/V4/V3/A3/M2/s1 ),
    .A2(\V2/V4/V3/A3/c1 ),
    .ZN(\V2/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M2/M2/_1_  (.A(\V2/V4/V3/A3/M2/s1 ),
    .B(\V2/V4/V3/A3/c1 ),
    .Z(\V2/V4/v3 [5]));
 OR2_X1 \V2/V4/V3/A3/M2/_0_  (.A1(\V2/V4/V3/A3/M2/c1 ),
    .A2(\V2/V4/V3/A3/M2/c2 ),
    .ZN(\V2/V4/V3/A3/c2 ));
 AND2_X1 \V2/V4/V3/A3/M3/M1/_0_  (.A1(\V2/V4/V3/v4 [2]),
    .A2(\V2/V4/V3/c3 ),
    .ZN(\V2/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M3/M1/_1_  (.A(\V2/V4/V3/v4 [2]),
    .B(\V2/V4/V3/c3 ),
    .Z(\V2/V4/V3/A3/M3/s1 ));
 AND2_X1 \V2/V4/V3/A3/M3/M2/_0_  (.A1(\V2/V4/V3/A3/M3/s1 ),
    .A2(\V2/V4/V3/A3/c2 ),
    .ZN(\V2/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M3/M2/_1_  (.A(\V2/V4/V3/A3/M3/s1 ),
    .B(\V2/V4/V3/A3/c2 ),
    .Z(\V2/V4/v3 [6]));
 OR2_X1 \V2/V4/V3/A3/M3/_0_  (.A1(\V2/V4/V3/A3/M3/c1 ),
    .A2(\V2/V4/V3/A3/M3/c2 ),
    .ZN(\V2/V4/V3/A3/c3 ));
 AND2_X1 \V2/V4/V3/A3/M4/M1/_0_  (.A1(\V2/V4/V3/v4 [3]),
    .A2(ground),
    .ZN(\V2/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M4/M1/_1_  (.A(\V2/V4/V3/v4 [3]),
    .B(ground),
    .Z(\V2/V4/V3/A3/M4/s1 ));
 AND2_X1 \V2/V4/V3/A3/M4/M2/_0_  (.A1(\V2/V4/V3/A3/M4/s1 ),
    .A2(\V2/V4/V3/A3/c3 ),
    .ZN(\V2/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M4/M2/_1_  (.A(\V2/V4/V3/A3/M4/s1 ),
    .B(\V2/V4/V3/A3/c3 ),
    .Z(\V2/V4/v3 [7]));
 OR2_X1 \V2/V4/V3/A3/M4/_0_  (.A1(\V2/V4/V3/A3/M4/c1 ),
    .A2(\V2/V4/V3/A3/M4/c2 ),
    .ZN(\V2/V4/V3/overflow ));
 AND2_X1 \V2/V4/V3/V1/HA1/_0_  (.A1(\V2/V4/V3/V1/w2 ),
    .A2(\V2/V4/V3/V1/w1 ),
    .ZN(\V2/V4/V3/V1/w4 ));
 XOR2_X2 \V2/V4/V3/V1/HA1/_1_  (.A(\V2/V4/V3/V1/w2 ),
    .B(\V2/V4/V3/V1/w1 ),
    .Z(\V2/V4/v3 [1]));
 AND2_X1 \V2/V4/V3/V1/HA2/_0_  (.A1(\V2/V4/V3/V1/w4 ),
    .A2(\V2/V4/V3/V1/w3 ),
    .ZN(\V2/V4/V3/v1 [3]));
 XOR2_X2 \V2/V4/V3/V1/HA2/_1_  (.A(\V2/V4/V3/V1/w4 ),
    .B(\V2/V4/V3/V1/w3 ),
    .Z(\V2/V4/V3/v1 [2]));
 AND2_X1 \V2/V4/V3/V1/_0_  (.A1(A[24]),
    .A2(B[12]),
    .ZN(\V2/V4/v3 [0]));
 AND2_X1 \V2/V4/V3/V1/_1_  (.A1(A[24]),
    .A2(B[13]),
    .ZN(\V2/V4/V3/V1/w1 ));
 AND2_X1 \V2/V4/V3/V1/_2_  (.A1(B[12]),
    .A2(A[25]),
    .ZN(\V2/V4/V3/V1/w2 ));
 AND2_X1 \V2/V4/V3/V1/_3_  (.A1(B[13]),
    .A2(A[25]),
    .ZN(\V2/V4/V3/V1/w3 ));
 AND2_X1 \V2/V4/V3/V2/HA1/_0_  (.A1(\V2/V4/V3/V2/w2 ),
    .A2(\V2/V4/V3/V2/w1 ),
    .ZN(\V2/V4/V3/V2/w4 ));
 XOR2_X2 \V2/V4/V3/V2/HA1/_1_  (.A(\V2/V4/V3/V2/w2 ),
    .B(\V2/V4/V3/V2/w1 ),
    .Z(\V2/V4/V3/v2 [1]));
 AND2_X1 \V2/V4/V3/V2/HA2/_0_  (.A1(\V2/V4/V3/V2/w4 ),
    .A2(\V2/V4/V3/V2/w3 ),
    .ZN(\V2/V4/V3/v2 [3]));
 XOR2_X2 \V2/V4/V3/V2/HA2/_1_  (.A(\V2/V4/V3/V2/w4 ),
    .B(\V2/V4/V3/V2/w3 ),
    .Z(\V2/V4/V3/v2 [2]));
 AND2_X1 \V2/V4/V3/V2/_0_  (.A1(A[26]),
    .A2(B[12]),
    .ZN(\V2/V4/V3/v2 [0]));
 AND2_X1 \V2/V4/V3/V2/_1_  (.A1(A[26]),
    .A2(B[13]),
    .ZN(\V2/V4/V3/V2/w1 ));
 AND2_X1 \V2/V4/V3/V2/_2_  (.A1(B[12]),
    .A2(A[27]),
    .ZN(\V2/V4/V3/V2/w2 ));
 AND2_X1 \V2/V4/V3/V2/_3_  (.A1(B[13]),
    .A2(A[27]),
    .ZN(\V2/V4/V3/V2/w3 ));
 AND2_X1 \V2/V4/V3/V3/HA1/_0_  (.A1(\V2/V4/V3/V3/w2 ),
    .A2(\V2/V4/V3/V3/w1 ),
    .ZN(\V2/V4/V3/V3/w4 ));
 XOR2_X2 \V2/V4/V3/V3/HA1/_1_  (.A(\V2/V4/V3/V3/w2 ),
    .B(\V2/V4/V3/V3/w1 ),
    .Z(\V2/V4/V3/v3 [1]));
 AND2_X1 \V2/V4/V3/V3/HA2/_0_  (.A1(\V2/V4/V3/V3/w4 ),
    .A2(\V2/V4/V3/V3/w3 ),
    .ZN(\V2/V4/V3/v3 [3]));
 XOR2_X2 \V2/V4/V3/V3/HA2/_1_  (.A(\V2/V4/V3/V3/w4 ),
    .B(\V2/V4/V3/V3/w3 ),
    .Z(\V2/V4/V3/v3 [2]));
 AND2_X1 \V2/V4/V3/V3/_0_  (.A1(A[24]),
    .A2(B[14]),
    .ZN(\V2/V4/V3/v3 [0]));
 AND2_X1 \V2/V4/V3/V3/_1_  (.A1(A[24]),
    .A2(B[15]),
    .ZN(\V2/V4/V3/V3/w1 ));
 AND2_X1 \V2/V4/V3/V3/_2_  (.A1(B[14]),
    .A2(A[25]),
    .ZN(\V2/V4/V3/V3/w2 ));
 AND2_X1 \V2/V4/V3/V3/_3_  (.A1(B[15]),
    .A2(A[25]),
    .ZN(\V2/V4/V3/V3/w3 ));
 AND2_X1 \V2/V4/V3/V4/HA1/_0_  (.A1(\V2/V4/V3/V4/w2 ),
    .A2(\V2/V4/V3/V4/w1 ),
    .ZN(\V2/V4/V3/V4/w4 ));
 XOR2_X2 \V2/V4/V3/V4/HA1/_1_  (.A(\V2/V4/V3/V4/w2 ),
    .B(\V2/V4/V3/V4/w1 ),
    .Z(\V2/V4/V3/v4 [1]));
 AND2_X1 \V2/V4/V3/V4/HA2/_0_  (.A1(\V2/V4/V3/V4/w4 ),
    .A2(\V2/V4/V3/V4/w3 ),
    .ZN(\V2/V4/V3/v4 [3]));
 XOR2_X2 \V2/V4/V3/V4/HA2/_1_  (.A(\V2/V4/V3/V4/w4 ),
    .B(\V2/V4/V3/V4/w3 ),
    .Z(\V2/V4/V3/v4 [2]));
 AND2_X1 \V2/V4/V3/V4/_0_  (.A1(A[26]),
    .A2(B[14]),
    .ZN(\V2/V4/V3/v4 [0]));
 AND2_X1 \V2/V4/V3/V4/_1_  (.A1(A[26]),
    .A2(B[15]),
    .ZN(\V2/V4/V3/V4/w1 ));
 AND2_X1 \V2/V4/V3/V4/_2_  (.A1(B[14]),
    .A2(A[27]),
    .ZN(\V2/V4/V3/V4/w2 ));
 AND2_X1 \V2/V4/V3/V4/_3_  (.A1(B[15]),
    .A2(A[27]),
    .ZN(\V2/V4/V3/V4/w3 ));
 OR2_X1 \V2/V4/V3/_0_  (.A1(\V2/V4/V3/c1 ),
    .A2(\V2/V4/V3/c2 ),
    .ZN(\V2/V4/V3/c3 ));
 AND2_X1 \V2/V4/V4/A1/M1/M1/_0_  (.A1(\V2/V4/V4/v2 [0]),
    .A2(\V2/V4/V4/v3 [0]),
    .ZN(\V2/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M1/M1/_1_  (.A(\V2/V4/V4/v2 [0]),
    .B(\V2/V4/V4/v3 [0]),
    .Z(\V2/V4/V4/A1/M1/s1 ));
 AND2_X1 \V2/V4/V4/A1/M1/M2/_0_  (.A1(\V2/V4/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M1/M2/_1_  (.A(\V2/V4/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/V4/s1 [0]));
 OR2_X1 \V2/V4/V4/A1/M1/_0_  (.A1(\V2/V4/V4/A1/M1/c1 ),
    .A2(\V2/V4/V4/A1/M1/c2 ),
    .ZN(\V2/V4/V4/A1/c1 ));
 AND2_X1 \V2/V4/V4/A1/M2/M1/_0_  (.A1(\V2/V4/V4/v2 [1]),
    .A2(\V2/V4/V4/v3 [1]),
    .ZN(\V2/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M2/M1/_1_  (.A(\V2/V4/V4/v2 [1]),
    .B(\V2/V4/V4/v3 [1]),
    .Z(\V2/V4/V4/A1/M2/s1 ));
 AND2_X1 \V2/V4/V4/A1/M2/M2/_0_  (.A1(\V2/V4/V4/A1/M2/s1 ),
    .A2(\V2/V4/V4/A1/c1 ),
    .ZN(\V2/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M2/M2/_1_  (.A(\V2/V4/V4/A1/M2/s1 ),
    .B(\V2/V4/V4/A1/c1 ),
    .Z(\V2/V4/V4/s1 [1]));
 OR2_X1 \V2/V4/V4/A1/M2/_0_  (.A1(\V2/V4/V4/A1/M2/c1 ),
    .A2(\V2/V4/V4/A1/M2/c2 ),
    .ZN(\V2/V4/V4/A1/c2 ));
 AND2_X1 \V2/V4/V4/A1/M3/M1/_0_  (.A1(\V2/V4/V4/v2 [2]),
    .A2(\V2/V4/V4/v3 [2]),
    .ZN(\V2/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M3/M1/_1_  (.A(\V2/V4/V4/v2 [2]),
    .B(\V2/V4/V4/v3 [2]),
    .Z(\V2/V4/V4/A1/M3/s1 ));
 AND2_X1 \V2/V4/V4/A1/M3/M2/_0_  (.A1(\V2/V4/V4/A1/M3/s1 ),
    .A2(\V2/V4/V4/A1/c2 ),
    .ZN(\V2/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M3/M2/_1_  (.A(\V2/V4/V4/A1/M3/s1 ),
    .B(\V2/V4/V4/A1/c2 ),
    .Z(\V2/V4/V4/s1 [2]));
 OR2_X1 \V2/V4/V4/A1/M3/_0_  (.A1(\V2/V4/V4/A1/M3/c1 ),
    .A2(\V2/V4/V4/A1/M3/c2 ),
    .ZN(\V2/V4/V4/A1/c3 ));
 AND2_X1 \V2/V4/V4/A1/M4/M1/_0_  (.A1(\V2/V4/V4/v2 [3]),
    .A2(\V2/V4/V4/v3 [3]),
    .ZN(\V2/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M4/M1/_1_  (.A(\V2/V4/V4/v2 [3]),
    .B(\V2/V4/V4/v3 [3]),
    .Z(\V2/V4/V4/A1/M4/s1 ));
 AND2_X1 \V2/V4/V4/A1/M4/M2/_0_  (.A1(\V2/V4/V4/A1/M4/s1 ),
    .A2(\V2/V4/V4/A1/c3 ),
    .ZN(\V2/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M4/M2/_1_  (.A(\V2/V4/V4/A1/M4/s1 ),
    .B(\V2/V4/V4/A1/c3 ),
    .Z(\V2/V4/V4/s1 [3]));
 OR2_X1 \V2/V4/V4/A1/M4/_0_  (.A1(\V2/V4/V4/A1/M4/c1 ),
    .A2(\V2/V4/V4/A1/M4/c2 ),
    .ZN(\V2/V4/V4/c1 ));
 AND2_X1 \V2/V4/V4/A2/M1/M1/_0_  (.A1(\V2/V4/V4/s1 [0]),
    .A2(\V2/V4/V4/v1 [2]),
    .ZN(\V2/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M1/M1/_1_  (.A(\V2/V4/V4/s1 [0]),
    .B(\V2/V4/V4/v1 [2]),
    .Z(\V2/V4/V4/A2/M1/s1 ));
 AND2_X1 \V2/V4/V4/A2/M1/M2/_0_  (.A1(\V2/V4/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M1/M2/_1_  (.A(\V2/V4/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v4 [2]));
 OR2_X1 \V2/V4/V4/A2/M1/_0_  (.A1(\V2/V4/V4/A2/M1/c1 ),
    .A2(\V2/V4/V4/A2/M1/c2 ),
    .ZN(\V2/V4/V4/A2/c1 ));
 AND2_X1 \V2/V4/V4/A2/M2/M1/_0_  (.A1(\V2/V4/V4/s1 [1]),
    .A2(\V2/V4/V4/v1 [3]),
    .ZN(\V2/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M2/M1/_1_  (.A(\V2/V4/V4/s1 [1]),
    .B(\V2/V4/V4/v1 [3]),
    .Z(\V2/V4/V4/A2/M2/s1 ));
 AND2_X1 \V2/V4/V4/A2/M2/M2/_0_  (.A1(\V2/V4/V4/A2/M2/s1 ),
    .A2(\V2/V4/V4/A2/c1 ),
    .ZN(\V2/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M2/M2/_1_  (.A(\V2/V4/V4/A2/M2/s1 ),
    .B(\V2/V4/V4/A2/c1 ),
    .Z(\V2/V4/v4 [3]));
 OR2_X1 \V2/V4/V4/A2/M2/_0_  (.A1(\V2/V4/V4/A2/M2/c1 ),
    .A2(\V2/V4/V4/A2/M2/c2 ),
    .ZN(\V2/V4/V4/A2/c2 ));
 AND2_X1 \V2/V4/V4/A2/M3/M1/_0_  (.A1(\V2/V4/V4/s1 [2]),
    .A2(ground),
    .ZN(\V2/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M3/M1/_1_  (.A(\V2/V4/V4/s1 [2]),
    .B(ground),
    .Z(\V2/V4/V4/A2/M3/s1 ));
 AND2_X1 \V2/V4/V4/A2/M3/M2/_0_  (.A1(\V2/V4/V4/A2/M3/s1 ),
    .A2(\V2/V4/V4/A2/c2 ),
    .ZN(\V2/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M3/M2/_1_  (.A(\V2/V4/V4/A2/M3/s1 ),
    .B(\V2/V4/V4/A2/c2 ),
    .Z(\V2/V4/V4/s2 [2]));
 OR2_X1 \V2/V4/V4/A2/M3/_0_  (.A1(\V2/V4/V4/A2/M3/c1 ),
    .A2(\V2/V4/V4/A2/M3/c2 ),
    .ZN(\V2/V4/V4/A2/c3 ));
 AND2_X1 \V2/V4/V4/A2/M4/M1/_0_  (.A1(\V2/V4/V4/s1 [3]),
    .A2(ground),
    .ZN(\V2/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M4/M1/_1_  (.A(\V2/V4/V4/s1 [3]),
    .B(ground),
    .Z(\V2/V4/V4/A2/M4/s1 ));
 AND2_X1 \V2/V4/V4/A2/M4/M2/_0_  (.A1(\V2/V4/V4/A2/M4/s1 ),
    .A2(\V2/V4/V4/A2/c3 ),
    .ZN(\V2/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M4/M2/_1_  (.A(\V2/V4/V4/A2/M4/s1 ),
    .B(\V2/V4/V4/A2/c3 ),
    .Z(\V2/V4/V4/s2 [3]));
 OR2_X1 \V2/V4/V4/A2/M4/_0_  (.A1(\V2/V4/V4/A2/M4/c1 ),
    .A2(\V2/V4/V4/A2/M4/c2 ),
    .ZN(\V2/V4/V4/c2 ));
 AND2_X1 \V2/V4/V4/A3/M1/M1/_0_  (.A1(\V2/V4/V4/v4 [0]),
    .A2(\V2/V4/V4/s2 [2]),
    .ZN(\V2/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M1/M1/_1_  (.A(\V2/V4/V4/v4 [0]),
    .B(\V2/V4/V4/s2 [2]),
    .Z(\V2/V4/V4/A3/M1/s1 ));
 AND2_X1 \V2/V4/V4/A3/M1/M2/_0_  (.A1(\V2/V4/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V2/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M1/M2/_1_  (.A(\V2/V4/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V2/V4/v4 [4]));
 OR2_X1 \V2/V4/V4/A3/M1/_0_  (.A1(\V2/V4/V4/A3/M1/c1 ),
    .A2(\V2/V4/V4/A3/M1/c2 ),
    .ZN(\V2/V4/V4/A3/c1 ));
 AND2_X1 \V2/V4/V4/A3/M2/M1/_0_  (.A1(\V2/V4/V4/v4 [1]),
    .A2(\V2/V4/V4/s2 [3]),
    .ZN(\V2/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M2/M1/_1_  (.A(\V2/V4/V4/v4 [1]),
    .B(\V2/V4/V4/s2 [3]),
    .Z(\V2/V4/V4/A3/M2/s1 ));
 AND2_X1 \V2/V4/V4/A3/M2/M2/_0_  (.A1(\V2/V4/V4/A3/M2/s1 ),
    .A2(\V2/V4/V4/A3/c1 ),
    .ZN(\V2/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M2/M2/_1_  (.A(\V2/V4/V4/A3/M2/s1 ),
    .B(\V2/V4/V4/A3/c1 ),
    .Z(\V2/V4/v4 [5]));
 OR2_X1 \V2/V4/V4/A3/M2/_0_  (.A1(\V2/V4/V4/A3/M2/c1 ),
    .A2(\V2/V4/V4/A3/M2/c2 ),
    .ZN(\V2/V4/V4/A3/c2 ));
 AND2_X1 \V2/V4/V4/A3/M3/M1/_0_  (.A1(\V2/V4/V4/v4 [2]),
    .A2(\V2/V4/V4/c3 ),
    .ZN(\V2/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M3/M1/_1_  (.A(\V2/V4/V4/v4 [2]),
    .B(\V2/V4/V4/c3 ),
    .Z(\V2/V4/V4/A3/M3/s1 ));
 AND2_X1 \V2/V4/V4/A3/M3/M2/_0_  (.A1(\V2/V4/V4/A3/M3/s1 ),
    .A2(\V2/V4/V4/A3/c2 ),
    .ZN(\V2/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M3/M2/_1_  (.A(\V2/V4/V4/A3/M3/s1 ),
    .B(\V2/V4/V4/A3/c2 ),
    .Z(\V2/V4/v4 [6]));
 OR2_X1 \V2/V4/V4/A3/M3/_0_  (.A1(\V2/V4/V4/A3/M3/c1 ),
    .A2(\V2/V4/V4/A3/M3/c2 ),
    .ZN(\V2/V4/V4/A3/c3 ));
 AND2_X1 \V2/V4/V4/A3/M4/M1/_0_  (.A1(\V2/V4/V4/v4 [3]),
    .A2(ground),
    .ZN(\V2/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M4/M1/_1_  (.A(\V2/V4/V4/v4 [3]),
    .B(ground),
    .Z(\V2/V4/V4/A3/M4/s1 ));
 AND2_X1 \V2/V4/V4/A3/M4/M2/_0_  (.A1(\V2/V4/V4/A3/M4/s1 ),
    .A2(\V2/V4/V4/A3/c3 ),
    .ZN(\V2/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M4/M2/_1_  (.A(\V2/V4/V4/A3/M4/s1 ),
    .B(\V2/V4/V4/A3/c3 ),
    .Z(\V2/V4/v4 [7]));
 OR2_X1 \V2/V4/V4/A3/M4/_0_  (.A1(\V2/V4/V4/A3/M4/c1 ),
    .A2(\V2/V4/V4/A3/M4/c2 ),
    .ZN(\V2/V4/V4/overflow ));
 AND2_X1 \V2/V4/V4/V1/HA1/_0_  (.A1(\V2/V4/V4/V1/w2 ),
    .A2(\V2/V4/V4/V1/w1 ),
    .ZN(\V2/V4/V4/V1/w4 ));
 XOR2_X2 \V2/V4/V4/V1/HA1/_1_  (.A(\V2/V4/V4/V1/w2 ),
    .B(\V2/V4/V4/V1/w1 ),
    .Z(\V2/V4/v4 [1]));
 AND2_X1 \V2/V4/V4/V1/HA2/_0_  (.A1(\V2/V4/V4/V1/w4 ),
    .A2(\V2/V4/V4/V1/w3 ),
    .ZN(\V2/V4/V4/v1 [3]));
 XOR2_X2 \V2/V4/V4/V1/HA2/_1_  (.A(\V2/V4/V4/V1/w4 ),
    .B(\V2/V4/V4/V1/w3 ),
    .Z(\V2/V4/V4/v1 [2]));
 AND2_X1 \V2/V4/V4/V1/_0_  (.A1(A[28]),
    .A2(B[12]),
    .ZN(\V2/V4/v4 [0]));
 AND2_X1 \V2/V4/V4/V1/_1_  (.A1(A[28]),
    .A2(B[13]),
    .ZN(\V2/V4/V4/V1/w1 ));
 AND2_X1 \V2/V4/V4/V1/_2_  (.A1(B[12]),
    .A2(A[29]),
    .ZN(\V2/V4/V4/V1/w2 ));
 AND2_X1 \V2/V4/V4/V1/_3_  (.A1(B[13]),
    .A2(A[29]),
    .ZN(\V2/V4/V4/V1/w3 ));
 AND2_X1 \V2/V4/V4/V2/HA1/_0_  (.A1(\V2/V4/V4/V2/w2 ),
    .A2(\V2/V4/V4/V2/w1 ),
    .ZN(\V2/V4/V4/V2/w4 ));
 XOR2_X2 \V2/V4/V4/V2/HA1/_1_  (.A(\V2/V4/V4/V2/w2 ),
    .B(\V2/V4/V4/V2/w1 ),
    .Z(\V2/V4/V4/v2 [1]));
 AND2_X1 \V2/V4/V4/V2/HA2/_0_  (.A1(\V2/V4/V4/V2/w4 ),
    .A2(\V2/V4/V4/V2/w3 ),
    .ZN(\V2/V4/V4/v2 [3]));
 XOR2_X2 \V2/V4/V4/V2/HA2/_1_  (.A(\V2/V4/V4/V2/w4 ),
    .B(\V2/V4/V4/V2/w3 ),
    .Z(\V2/V4/V4/v2 [2]));
 AND2_X1 \V2/V4/V4/V2/_0_  (.A1(A[30]),
    .A2(B[12]),
    .ZN(\V2/V4/V4/v2 [0]));
 AND2_X1 \V2/V4/V4/V2/_1_  (.A1(A[30]),
    .A2(B[13]),
    .ZN(\V2/V4/V4/V2/w1 ));
 AND2_X1 \V2/V4/V4/V2/_2_  (.A1(B[12]),
    .A2(A[31]),
    .ZN(\V2/V4/V4/V2/w2 ));
 AND2_X1 \V2/V4/V4/V2/_3_  (.A1(B[13]),
    .A2(A[31]),
    .ZN(\V2/V4/V4/V2/w3 ));
 AND2_X1 \V2/V4/V4/V3/HA1/_0_  (.A1(\V2/V4/V4/V3/w2 ),
    .A2(\V2/V4/V4/V3/w1 ),
    .ZN(\V2/V4/V4/V3/w4 ));
 XOR2_X2 \V2/V4/V4/V3/HA1/_1_  (.A(\V2/V4/V4/V3/w2 ),
    .B(\V2/V4/V4/V3/w1 ),
    .Z(\V2/V4/V4/v3 [1]));
 AND2_X1 \V2/V4/V4/V3/HA2/_0_  (.A1(\V2/V4/V4/V3/w4 ),
    .A2(\V2/V4/V4/V3/w3 ),
    .ZN(\V2/V4/V4/v3 [3]));
 XOR2_X2 \V2/V4/V4/V3/HA2/_1_  (.A(\V2/V4/V4/V3/w4 ),
    .B(\V2/V4/V4/V3/w3 ),
    .Z(\V2/V4/V4/v3 [2]));
 AND2_X1 \V2/V4/V4/V3/_0_  (.A1(A[28]),
    .A2(B[14]),
    .ZN(\V2/V4/V4/v3 [0]));
 AND2_X1 \V2/V4/V4/V3/_1_  (.A1(A[28]),
    .A2(B[15]),
    .ZN(\V2/V4/V4/V3/w1 ));
 AND2_X1 \V2/V4/V4/V3/_2_  (.A1(B[14]),
    .A2(A[29]),
    .ZN(\V2/V4/V4/V3/w2 ));
 AND2_X1 \V2/V4/V4/V3/_3_  (.A1(B[15]),
    .A2(A[29]),
    .ZN(\V2/V4/V4/V3/w3 ));
 AND2_X1 \V2/V4/V4/V4/HA1/_0_  (.A1(\V2/V4/V4/V4/w2 ),
    .A2(\V2/V4/V4/V4/w1 ),
    .ZN(\V2/V4/V4/V4/w4 ));
 XOR2_X2 \V2/V4/V4/V4/HA1/_1_  (.A(\V2/V4/V4/V4/w2 ),
    .B(\V2/V4/V4/V4/w1 ),
    .Z(\V2/V4/V4/v4 [1]));
 AND2_X1 \V2/V4/V4/V4/HA2/_0_  (.A1(\V2/V4/V4/V4/w4 ),
    .A2(\V2/V4/V4/V4/w3 ),
    .ZN(\V2/V4/V4/v4 [3]));
 XOR2_X2 \V2/V4/V4/V4/HA2/_1_  (.A(\V2/V4/V4/V4/w4 ),
    .B(\V2/V4/V4/V4/w3 ),
    .Z(\V2/V4/V4/v4 [2]));
 AND2_X1 \V2/V4/V4/V4/_0_  (.A1(A[30]),
    .A2(B[14]),
    .ZN(\V2/V4/V4/v4 [0]));
 AND2_X1 \V2/V4/V4/V4/_1_  (.A1(A[30]),
    .A2(B[15]),
    .ZN(\V2/V4/V4/V4/w1 ));
 AND2_X1 \V2/V4/V4/V4/_2_  (.A1(B[14]),
    .A2(A[31]),
    .ZN(\V2/V4/V4/V4/w2 ));
 AND2_X1 \V2/V4/V4/V4/_3_  (.A1(B[15]),
    .A2(A[31]),
    .ZN(\V2/V4/V4/V4/w3 ));
 OR2_X1 \V2/V4/V4/_0_  (.A1(\V2/V4/V4/c1 ),
    .A2(\V2/V4/V4/c2 ),
    .ZN(\V2/V4/V4/c3 ));
 OR2_X1 \V2/V4/_0_  (.A1(\V2/V4/c1 ),
    .A2(\V2/V4/c2 ),
    .ZN(\V2/V4/c3 ));
 OR2_X1 \V2/_0_  (.A1(\V2/c1 ),
    .A2(\V2/c2 ),
    .ZN(\V2/c3 ));
 AND2_X1 \V3/A1/A1/A1/M1/M1/_0_  (.A1(\V3/v2 [0]),
    .A2(\V3/v3 [0]),
    .ZN(\V3/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M1/M1/_1_  (.A(\V3/v2 [0]),
    .B(\V3/v3 [0]),
    .Z(\V3/A1/A1/A1/M1/s1 ));
 AND2_X1 \V3/A1/A1/A1/M1/M2/_0_  (.A1(\V3/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M1/M2/_1_  (.A(\V3/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/s1 [0]));
 OR2_X1 \V3/A1/A1/A1/M1/_0_  (.A1(\V3/A1/A1/A1/M1/c1 ),
    .A2(\V3/A1/A1/A1/M1/c2 ),
    .ZN(\V3/A1/A1/A1/c1 ));
 AND2_X1 \V3/A1/A1/A1/M2/M1/_0_  (.A1(\V3/v2 [1]),
    .A2(\V3/v3 [1]),
    .ZN(\V3/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M2/M1/_1_  (.A(\V3/v2 [1]),
    .B(\V3/v3 [1]),
    .Z(\V3/A1/A1/A1/M2/s1 ));
 AND2_X1 \V3/A1/A1/A1/M2/M2/_0_  (.A1(\V3/A1/A1/A1/M2/s1 ),
    .A2(\V3/A1/A1/A1/c1 ),
    .ZN(\V3/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M2/M2/_1_  (.A(\V3/A1/A1/A1/M2/s1 ),
    .B(\V3/A1/A1/A1/c1 ),
    .Z(\V3/s1 [1]));
 OR2_X1 \V3/A1/A1/A1/M2/_0_  (.A1(\V3/A1/A1/A1/M2/c1 ),
    .A2(\V3/A1/A1/A1/M2/c2 ),
    .ZN(\V3/A1/A1/A1/c2 ));
 AND2_X1 \V3/A1/A1/A1/M3/M1/_0_  (.A1(\V3/v2 [2]),
    .A2(\V3/v3 [2]),
    .ZN(\V3/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M3/M1/_1_  (.A(\V3/v2 [2]),
    .B(\V3/v3 [2]),
    .Z(\V3/A1/A1/A1/M3/s1 ));
 AND2_X1 \V3/A1/A1/A1/M3/M2/_0_  (.A1(\V3/A1/A1/A1/M3/s1 ),
    .A2(\V3/A1/A1/A1/c2 ),
    .ZN(\V3/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M3/M2/_1_  (.A(\V3/A1/A1/A1/M3/s1 ),
    .B(\V3/A1/A1/A1/c2 ),
    .Z(\V3/s1 [2]));
 OR2_X1 \V3/A1/A1/A1/M3/_0_  (.A1(\V3/A1/A1/A1/M3/c1 ),
    .A2(\V3/A1/A1/A1/M3/c2 ),
    .ZN(\V3/A1/A1/A1/c3 ));
 AND2_X1 \V3/A1/A1/A1/M4/M1/_0_  (.A1(\V3/v2 [3]),
    .A2(\V3/v3 [3]),
    .ZN(\V3/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M4/M1/_1_  (.A(\V3/v2 [3]),
    .B(\V3/v3 [3]),
    .Z(\V3/A1/A1/A1/M4/s1 ));
 AND2_X1 \V3/A1/A1/A1/M4/M2/_0_  (.A1(\V3/A1/A1/A1/M4/s1 ),
    .A2(\V3/A1/A1/A1/c3 ),
    .ZN(\V3/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M4/M2/_1_  (.A(\V3/A1/A1/A1/M4/s1 ),
    .B(\V3/A1/A1/A1/c3 ),
    .Z(\V3/s1 [3]));
 OR2_X1 \V3/A1/A1/A1/M4/_0_  (.A1(\V3/A1/A1/A1/M4/c1 ),
    .A2(\V3/A1/A1/A1/M4/c2 ),
    .ZN(\V3/A1/A1/c1 ));
 AND2_X1 \V3/A1/A1/A2/M1/M1/_0_  (.A1(\V3/v2 [4]),
    .A2(\V3/v3 [4]),
    .ZN(\V3/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M1/M1/_1_  (.A(\V3/v2 [4]),
    .B(\V3/v3 [4]),
    .Z(\V3/A1/A1/A2/M1/s1 ));
 AND2_X1 \V3/A1/A1/A2/M1/M2/_0_  (.A1(\V3/A1/A1/A2/M1/s1 ),
    .A2(\V3/A1/A1/c1 ),
    .ZN(\V3/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M1/M2/_1_  (.A(\V3/A1/A1/A2/M1/s1 ),
    .B(\V3/A1/A1/c1 ),
    .Z(\V3/s1 [4]));
 OR2_X1 \V3/A1/A1/A2/M1/_0_  (.A1(\V3/A1/A1/A2/M1/c1 ),
    .A2(\V3/A1/A1/A2/M1/c2 ),
    .ZN(\V3/A1/A1/A2/c1 ));
 AND2_X1 \V3/A1/A1/A2/M2/M1/_0_  (.A1(\V3/v2 [5]),
    .A2(\V3/v3 [5]),
    .ZN(\V3/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M2/M1/_1_  (.A(\V3/v2 [5]),
    .B(\V3/v3 [5]),
    .Z(\V3/A1/A1/A2/M2/s1 ));
 AND2_X1 \V3/A1/A1/A2/M2/M2/_0_  (.A1(\V3/A1/A1/A2/M2/s1 ),
    .A2(\V3/A1/A1/A2/c1 ),
    .ZN(\V3/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M2/M2/_1_  (.A(\V3/A1/A1/A2/M2/s1 ),
    .B(\V3/A1/A1/A2/c1 ),
    .Z(\V3/s1 [5]));
 OR2_X1 \V3/A1/A1/A2/M2/_0_  (.A1(\V3/A1/A1/A2/M2/c1 ),
    .A2(\V3/A1/A1/A2/M2/c2 ),
    .ZN(\V3/A1/A1/A2/c2 ));
 AND2_X1 \V3/A1/A1/A2/M3/M1/_0_  (.A1(\V3/v2 [6]),
    .A2(\V3/v3 [6]),
    .ZN(\V3/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M3/M1/_1_  (.A(\V3/v2 [6]),
    .B(\V3/v3 [6]),
    .Z(\V3/A1/A1/A2/M3/s1 ));
 AND2_X1 \V3/A1/A1/A2/M3/M2/_0_  (.A1(\V3/A1/A1/A2/M3/s1 ),
    .A2(\V3/A1/A1/A2/c2 ),
    .ZN(\V3/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M3/M2/_1_  (.A(\V3/A1/A1/A2/M3/s1 ),
    .B(\V3/A1/A1/A2/c2 ),
    .Z(\V3/s1 [6]));
 OR2_X1 \V3/A1/A1/A2/M3/_0_  (.A1(\V3/A1/A1/A2/M3/c1 ),
    .A2(\V3/A1/A1/A2/M3/c2 ),
    .ZN(\V3/A1/A1/A2/c3 ));
 AND2_X1 \V3/A1/A1/A2/M4/M1/_0_  (.A1(\V3/v2 [7]),
    .A2(\V3/v3 [7]),
    .ZN(\V3/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M4/M1/_1_  (.A(\V3/v2 [7]),
    .B(\V3/v3 [7]),
    .Z(\V3/A1/A1/A2/M4/s1 ));
 AND2_X1 \V3/A1/A1/A2/M4/M2/_0_  (.A1(\V3/A1/A1/A2/M4/s1 ),
    .A2(\V3/A1/A1/A2/c3 ),
    .ZN(\V3/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M4/M2/_1_  (.A(\V3/A1/A1/A2/M4/s1 ),
    .B(\V3/A1/A1/A2/c3 ),
    .Z(\V3/s1 [7]));
 OR2_X1 \V3/A1/A1/A2/M4/_0_  (.A1(\V3/A1/A1/A2/M4/c1 ),
    .A2(\V3/A1/A1/A2/M4/c2 ),
    .ZN(\V3/A1/c1 ));
 AND2_X1 \V3/A1/A2/A1/M1/M1/_0_  (.A1(\V3/v2 [8]),
    .A2(\V3/v3 [8]),
    .ZN(\V3/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M1/M1/_1_  (.A(\V3/v2 [8]),
    .B(\V3/v3 [8]),
    .Z(\V3/A1/A2/A1/M1/s1 ));
 AND2_X1 \V3/A1/A2/A1/M1/M2/_0_  (.A1(\V3/A1/A2/A1/M1/s1 ),
    .A2(\V3/A1/c1 ),
    .ZN(\V3/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M1/M2/_1_  (.A(\V3/A1/A2/A1/M1/s1 ),
    .B(\V3/A1/c1 ),
    .Z(\V3/s1 [8]));
 OR2_X1 \V3/A1/A2/A1/M1/_0_  (.A1(\V3/A1/A2/A1/M1/c1 ),
    .A2(\V3/A1/A2/A1/M1/c2 ),
    .ZN(\V3/A1/A2/A1/c1 ));
 AND2_X1 \V3/A1/A2/A1/M2/M1/_0_  (.A1(\V3/v2 [9]),
    .A2(\V3/v3 [9]),
    .ZN(\V3/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M2/M1/_1_  (.A(\V3/v2 [9]),
    .B(\V3/v3 [9]),
    .Z(\V3/A1/A2/A1/M2/s1 ));
 AND2_X1 \V3/A1/A2/A1/M2/M2/_0_  (.A1(\V3/A1/A2/A1/M2/s1 ),
    .A2(\V3/A1/A2/A1/c1 ),
    .ZN(\V3/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M2/M2/_1_  (.A(\V3/A1/A2/A1/M2/s1 ),
    .B(\V3/A1/A2/A1/c1 ),
    .Z(\V3/s1 [9]));
 OR2_X1 \V3/A1/A2/A1/M2/_0_  (.A1(\V3/A1/A2/A1/M2/c1 ),
    .A2(\V3/A1/A2/A1/M2/c2 ),
    .ZN(\V3/A1/A2/A1/c2 ));
 AND2_X1 \V3/A1/A2/A1/M3/M1/_0_  (.A1(\V3/v2 [10]),
    .A2(\V3/v3 [10]),
    .ZN(\V3/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M3/M1/_1_  (.A(\V3/v2 [10]),
    .B(\V3/v3 [10]),
    .Z(\V3/A1/A2/A1/M3/s1 ));
 AND2_X1 \V3/A1/A2/A1/M3/M2/_0_  (.A1(\V3/A1/A2/A1/M3/s1 ),
    .A2(\V3/A1/A2/A1/c2 ),
    .ZN(\V3/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M3/M2/_1_  (.A(\V3/A1/A2/A1/M3/s1 ),
    .B(\V3/A1/A2/A1/c2 ),
    .Z(\V3/s1 [10]));
 OR2_X1 \V3/A1/A2/A1/M3/_0_  (.A1(\V3/A1/A2/A1/M3/c1 ),
    .A2(\V3/A1/A2/A1/M3/c2 ),
    .ZN(\V3/A1/A2/A1/c3 ));
 AND2_X1 \V3/A1/A2/A1/M4/M1/_0_  (.A1(\V3/v2 [11]),
    .A2(\V3/v3 [11]),
    .ZN(\V3/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M4/M1/_1_  (.A(\V3/v2 [11]),
    .B(\V3/v3 [11]),
    .Z(\V3/A1/A2/A1/M4/s1 ));
 AND2_X1 \V3/A1/A2/A1/M4/M2/_0_  (.A1(\V3/A1/A2/A1/M4/s1 ),
    .A2(\V3/A1/A2/A1/c3 ),
    .ZN(\V3/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M4/M2/_1_  (.A(\V3/A1/A2/A1/M4/s1 ),
    .B(\V3/A1/A2/A1/c3 ),
    .Z(\V3/s1 [11]));
 OR2_X1 \V3/A1/A2/A1/M4/_0_  (.A1(\V3/A1/A2/A1/M4/c1 ),
    .A2(\V3/A1/A2/A1/M4/c2 ),
    .ZN(\V3/A1/A2/c1 ));
 AND2_X1 \V3/A1/A2/A2/M1/M1/_0_  (.A1(\V3/v2 [12]),
    .A2(\V3/v3 [12]),
    .ZN(\V3/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M1/M1/_1_  (.A(\V3/v2 [12]),
    .B(\V3/v3 [12]),
    .Z(\V3/A1/A2/A2/M1/s1 ));
 AND2_X1 \V3/A1/A2/A2/M1/M2/_0_  (.A1(\V3/A1/A2/A2/M1/s1 ),
    .A2(\V3/A1/A2/c1 ),
    .ZN(\V3/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M1/M2/_1_  (.A(\V3/A1/A2/A2/M1/s1 ),
    .B(\V3/A1/A2/c1 ),
    .Z(\V3/s1 [12]));
 OR2_X1 \V3/A1/A2/A2/M1/_0_  (.A1(\V3/A1/A2/A2/M1/c1 ),
    .A2(\V3/A1/A2/A2/M1/c2 ),
    .ZN(\V3/A1/A2/A2/c1 ));
 AND2_X1 \V3/A1/A2/A2/M2/M1/_0_  (.A1(\V3/v2 [13]),
    .A2(\V3/v3 [13]),
    .ZN(\V3/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M2/M1/_1_  (.A(\V3/v2 [13]),
    .B(\V3/v3 [13]),
    .Z(\V3/A1/A2/A2/M2/s1 ));
 AND2_X1 \V3/A1/A2/A2/M2/M2/_0_  (.A1(\V3/A1/A2/A2/M2/s1 ),
    .A2(\V3/A1/A2/A2/c1 ),
    .ZN(\V3/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M2/M2/_1_  (.A(\V3/A1/A2/A2/M2/s1 ),
    .B(\V3/A1/A2/A2/c1 ),
    .Z(\V3/s1 [13]));
 OR2_X1 \V3/A1/A2/A2/M2/_0_  (.A1(\V3/A1/A2/A2/M2/c1 ),
    .A2(\V3/A1/A2/A2/M2/c2 ),
    .ZN(\V3/A1/A2/A2/c2 ));
 AND2_X1 \V3/A1/A2/A2/M3/M1/_0_  (.A1(\V3/v2 [14]),
    .A2(\V3/v3 [14]),
    .ZN(\V3/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M3/M1/_1_  (.A(\V3/v2 [14]),
    .B(\V3/v3 [14]),
    .Z(\V3/A1/A2/A2/M3/s1 ));
 AND2_X1 \V3/A1/A2/A2/M3/M2/_0_  (.A1(\V3/A1/A2/A2/M3/s1 ),
    .A2(\V3/A1/A2/A2/c2 ),
    .ZN(\V3/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M3/M2/_1_  (.A(\V3/A1/A2/A2/M3/s1 ),
    .B(\V3/A1/A2/A2/c2 ),
    .Z(\V3/s1 [14]));
 OR2_X1 \V3/A1/A2/A2/M3/_0_  (.A1(\V3/A1/A2/A2/M3/c1 ),
    .A2(\V3/A1/A2/A2/M3/c2 ),
    .ZN(\V3/A1/A2/A2/c3 ));
 AND2_X1 \V3/A1/A2/A2/M4/M1/_0_  (.A1(\V3/v2 [15]),
    .A2(\V3/v3 [15]),
    .ZN(\V3/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M4/M1/_1_  (.A(\V3/v2 [15]),
    .B(\V3/v3 [15]),
    .Z(\V3/A1/A2/A2/M4/s1 ));
 AND2_X1 \V3/A1/A2/A2/M4/M2/_0_  (.A1(\V3/A1/A2/A2/M4/s1 ),
    .A2(\V3/A1/A2/A2/c3 ),
    .ZN(\V3/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M4/M2/_1_  (.A(\V3/A1/A2/A2/M4/s1 ),
    .B(\V3/A1/A2/A2/c3 ),
    .Z(\V3/s1 [15]));
 OR2_X1 \V3/A1/A2/A2/M4/_0_  (.A1(\V3/A1/A2/A2/M4/c1 ),
    .A2(\V3/A1/A2/A2/M4/c2 ),
    .ZN(\V3/c1 ));
 AND2_X1 \V3/A2/A1/A1/M1/M1/_0_  (.A1(\V3/s1 [0]),
    .A2(\V3/v1 [8]),
    .ZN(\V3/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M1/M1/_1_  (.A(\V3/s1 [0]),
    .B(\V3/v1 [8]),
    .Z(\V3/A2/A1/A1/M1/s1 ));
 AND2_X1 \V3/A2/A1/A1/M1/M2/_0_  (.A1(\V3/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M1/M2/_1_  (.A(\V3/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v3[8]));
 OR2_X1 \V3/A2/A1/A1/M1/_0_  (.A1(\V3/A2/A1/A1/M1/c1 ),
    .A2(\V3/A2/A1/A1/M1/c2 ),
    .ZN(\V3/A2/A1/A1/c1 ));
 AND2_X1 \V3/A2/A1/A1/M2/M1/_0_  (.A1(\V3/s1 [1]),
    .A2(\V3/v1 [9]),
    .ZN(\V3/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M2/M1/_1_  (.A(\V3/s1 [1]),
    .B(\V3/v1 [9]),
    .Z(\V3/A2/A1/A1/M2/s1 ));
 AND2_X1 \V3/A2/A1/A1/M2/M2/_0_  (.A1(\V3/A2/A1/A1/M2/s1 ),
    .A2(\V3/A2/A1/A1/c1 ),
    .ZN(\V3/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M2/M2/_1_  (.A(\V3/A2/A1/A1/M2/s1 ),
    .B(\V3/A2/A1/A1/c1 ),
    .Z(v3[9]));
 OR2_X1 \V3/A2/A1/A1/M2/_0_  (.A1(\V3/A2/A1/A1/M2/c1 ),
    .A2(\V3/A2/A1/A1/M2/c2 ),
    .ZN(\V3/A2/A1/A1/c2 ));
 AND2_X1 \V3/A2/A1/A1/M3/M1/_0_  (.A1(\V3/s1 [2]),
    .A2(\V3/v1 [10]),
    .ZN(\V3/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M3/M1/_1_  (.A(\V3/s1 [2]),
    .B(\V3/v1 [10]),
    .Z(\V3/A2/A1/A1/M3/s1 ));
 AND2_X1 \V3/A2/A1/A1/M3/M2/_0_  (.A1(\V3/A2/A1/A1/M3/s1 ),
    .A2(\V3/A2/A1/A1/c2 ),
    .ZN(\V3/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M3/M2/_1_  (.A(\V3/A2/A1/A1/M3/s1 ),
    .B(\V3/A2/A1/A1/c2 ),
    .Z(v3[10]));
 OR2_X1 \V3/A2/A1/A1/M3/_0_  (.A1(\V3/A2/A1/A1/M3/c1 ),
    .A2(\V3/A2/A1/A1/M3/c2 ),
    .ZN(\V3/A2/A1/A1/c3 ));
 AND2_X1 \V3/A2/A1/A1/M4/M1/_0_  (.A1(\V3/s1 [3]),
    .A2(\V3/v1 [11]),
    .ZN(\V3/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M4/M1/_1_  (.A(\V3/s1 [3]),
    .B(\V3/v1 [11]),
    .Z(\V3/A2/A1/A1/M4/s1 ));
 AND2_X1 \V3/A2/A1/A1/M4/M2/_0_  (.A1(\V3/A2/A1/A1/M4/s1 ),
    .A2(\V3/A2/A1/A1/c3 ),
    .ZN(\V3/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M4/M2/_1_  (.A(\V3/A2/A1/A1/M4/s1 ),
    .B(\V3/A2/A1/A1/c3 ),
    .Z(v3[11]));
 OR2_X1 \V3/A2/A1/A1/M4/_0_  (.A1(\V3/A2/A1/A1/M4/c1 ),
    .A2(\V3/A2/A1/A1/M4/c2 ),
    .ZN(\V3/A2/A1/c1 ));
 AND2_X1 \V3/A2/A1/A2/M1/M1/_0_  (.A1(\V3/s1 [4]),
    .A2(\V3/v1 [12]),
    .ZN(\V3/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M1/M1/_1_  (.A(\V3/s1 [4]),
    .B(\V3/v1 [12]),
    .Z(\V3/A2/A1/A2/M1/s1 ));
 AND2_X1 \V3/A2/A1/A2/M1/M2/_0_  (.A1(\V3/A2/A1/A2/M1/s1 ),
    .A2(\V3/A2/A1/c1 ),
    .ZN(\V3/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M1/M2/_1_  (.A(\V3/A2/A1/A2/M1/s1 ),
    .B(\V3/A2/A1/c1 ),
    .Z(v3[12]));
 OR2_X1 \V3/A2/A1/A2/M1/_0_  (.A1(\V3/A2/A1/A2/M1/c1 ),
    .A2(\V3/A2/A1/A2/M1/c2 ),
    .ZN(\V3/A2/A1/A2/c1 ));
 AND2_X1 \V3/A2/A1/A2/M2/M1/_0_  (.A1(\V3/s1 [5]),
    .A2(\V3/v1 [13]),
    .ZN(\V3/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M2/M1/_1_  (.A(\V3/s1 [5]),
    .B(\V3/v1 [13]),
    .Z(\V3/A2/A1/A2/M2/s1 ));
 AND2_X1 \V3/A2/A1/A2/M2/M2/_0_  (.A1(\V3/A2/A1/A2/M2/s1 ),
    .A2(\V3/A2/A1/A2/c1 ),
    .ZN(\V3/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M2/M2/_1_  (.A(\V3/A2/A1/A2/M2/s1 ),
    .B(\V3/A2/A1/A2/c1 ),
    .Z(v3[13]));
 OR2_X1 \V3/A2/A1/A2/M2/_0_  (.A1(\V3/A2/A1/A2/M2/c1 ),
    .A2(\V3/A2/A1/A2/M2/c2 ),
    .ZN(\V3/A2/A1/A2/c2 ));
 AND2_X1 \V3/A2/A1/A2/M3/M1/_0_  (.A1(\V3/s1 [6]),
    .A2(\V3/v1 [14]),
    .ZN(\V3/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M3/M1/_1_  (.A(\V3/s1 [6]),
    .B(\V3/v1 [14]),
    .Z(\V3/A2/A1/A2/M3/s1 ));
 AND2_X1 \V3/A2/A1/A2/M3/M2/_0_  (.A1(\V3/A2/A1/A2/M3/s1 ),
    .A2(\V3/A2/A1/A2/c2 ),
    .ZN(\V3/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M3/M2/_1_  (.A(\V3/A2/A1/A2/M3/s1 ),
    .B(\V3/A2/A1/A2/c2 ),
    .Z(v3[14]));
 OR2_X1 \V3/A2/A1/A2/M3/_0_  (.A1(\V3/A2/A1/A2/M3/c1 ),
    .A2(\V3/A2/A1/A2/M3/c2 ),
    .ZN(\V3/A2/A1/A2/c3 ));
 AND2_X1 \V3/A2/A1/A2/M4/M1/_0_  (.A1(\V3/s1 [7]),
    .A2(\V3/v1 [15]),
    .ZN(\V3/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M4/M1/_1_  (.A(\V3/s1 [7]),
    .B(\V3/v1 [15]),
    .Z(\V3/A2/A1/A2/M4/s1 ));
 AND2_X1 \V3/A2/A1/A2/M4/M2/_0_  (.A1(\V3/A2/A1/A2/M4/s1 ),
    .A2(\V3/A2/A1/A2/c3 ),
    .ZN(\V3/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M4/M2/_1_  (.A(\V3/A2/A1/A2/M4/s1 ),
    .B(\V3/A2/A1/A2/c3 ),
    .Z(v3[15]));
 OR2_X2 \V3/A2/A1/A2/M4/_0_  (.A1(\V3/A2/A1/A2/M4/c1 ),
    .A2(\V3/A2/A1/A2/M4/c2 ),
    .ZN(\V3/A2/c1 ));
 AND2_X1 \V3/A2/A2/A1/M1/M1/_0_  (.A1(\V3/s1 [8]),
    .A2(ground),
    .ZN(\V3/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M1/M1/_1_  (.A(\V3/s1 [8]),
    .B(ground),
    .Z(\V3/A2/A2/A1/M1/s1 ));
 AND2_X1 \V3/A2/A2/A1/M1/M2/_0_  (.A1(\V3/A2/A2/A1/M1/s1 ),
    .A2(\V3/A2/c1 ),
    .ZN(\V3/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M1/M2/_1_  (.A(\V3/A2/A2/A1/M1/s1 ),
    .B(\V3/A2/c1 ),
    .Z(\V3/s2 [8]));
 OR2_X1 \V3/A2/A2/A1/M1/_0_  (.A1(\V3/A2/A2/A1/M1/c1 ),
    .A2(\V3/A2/A2/A1/M1/c2 ),
    .ZN(\V3/A2/A2/A1/c1 ));
 AND2_X1 \V3/A2/A2/A1/M2/M1/_0_  (.A1(\V3/s1 [9]),
    .A2(ground),
    .ZN(\V3/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M2/M1/_1_  (.A(\V3/s1 [9]),
    .B(ground),
    .Z(\V3/A2/A2/A1/M2/s1 ));
 AND2_X1 \V3/A2/A2/A1/M2/M2/_0_  (.A1(\V3/A2/A2/A1/M2/s1 ),
    .A2(\V3/A2/A2/A1/c1 ),
    .ZN(\V3/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M2/M2/_1_  (.A(\V3/A2/A2/A1/M2/s1 ),
    .B(\V3/A2/A2/A1/c1 ),
    .Z(\V3/s2 [9]));
 OR2_X1 \V3/A2/A2/A1/M2/_0_  (.A1(\V3/A2/A2/A1/M2/c1 ),
    .A2(\V3/A2/A2/A1/M2/c2 ),
    .ZN(\V3/A2/A2/A1/c2 ));
 AND2_X1 \V3/A2/A2/A1/M3/M1/_0_  (.A1(\V3/s1 [10]),
    .A2(ground),
    .ZN(\V3/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M3/M1/_1_  (.A(\V3/s1 [10]),
    .B(ground),
    .Z(\V3/A2/A2/A1/M3/s1 ));
 AND2_X1 \V3/A2/A2/A1/M3/M2/_0_  (.A1(\V3/A2/A2/A1/M3/s1 ),
    .A2(\V3/A2/A2/A1/c2 ),
    .ZN(\V3/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M3/M2/_1_  (.A(\V3/A2/A2/A1/M3/s1 ),
    .B(\V3/A2/A2/A1/c2 ),
    .Z(\V3/s2 [10]));
 OR2_X1 \V3/A2/A2/A1/M3/_0_  (.A1(\V3/A2/A2/A1/M3/c1 ),
    .A2(\V3/A2/A2/A1/M3/c2 ),
    .ZN(\V3/A2/A2/A1/c3 ));
 AND2_X1 \V3/A2/A2/A1/M4/M1/_0_  (.A1(\V3/s1 [11]),
    .A2(ground),
    .ZN(\V3/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M4/M1/_1_  (.A(\V3/s1 [11]),
    .B(ground),
    .Z(\V3/A2/A2/A1/M4/s1 ));
 AND2_X1 \V3/A2/A2/A1/M4/M2/_0_  (.A1(\V3/A2/A2/A1/M4/s1 ),
    .A2(\V3/A2/A2/A1/c3 ),
    .ZN(\V3/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M4/M2/_1_  (.A(\V3/A2/A2/A1/M4/s1 ),
    .B(\V3/A2/A2/A1/c3 ),
    .Z(\V3/s2 [11]));
 OR2_X1 \V3/A2/A2/A1/M4/_0_  (.A1(\V3/A2/A2/A1/M4/c1 ),
    .A2(\V3/A2/A2/A1/M4/c2 ),
    .ZN(\V3/A2/A2/c1 ));
 AND2_X1 \V3/A2/A2/A2/M1/M1/_0_  (.A1(\V3/s1 [12]),
    .A2(ground),
    .ZN(\V3/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M1/M1/_1_  (.A(\V3/s1 [12]),
    .B(ground),
    .Z(\V3/A2/A2/A2/M1/s1 ));
 AND2_X1 \V3/A2/A2/A2/M1/M2/_0_  (.A1(\V3/A2/A2/A2/M1/s1 ),
    .A2(\V3/A2/A2/c1 ),
    .ZN(\V3/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M1/M2/_1_  (.A(\V3/A2/A2/A2/M1/s1 ),
    .B(\V3/A2/A2/c1 ),
    .Z(\V3/s2 [12]));
 OR2_X1 \V3/A2/A2/A2/M1/_0_  (.A1(\V3/A2/A2/A2/M1/c1 ),
    .A2(\V3/A2/A2/A2/M1/c2 ),
    .ZN(\V3/A2/A2/A2/c1 ));
 AND2_X1 \V3/A2/A2/A2/M2/M1/_0_  (.A1(\V3/s1 [13]),
    .A2(ground),
    .ZN(\V3/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M2/M1/_1_  (.A(\V3/s1 [13]),
    .B(ground),
    .Z(\V3/A2/A2/A2/M2/s1 ));
 AND2_X1 \V3/A2/A2/A2/M2/M2/_0_  (.A1(\V3/A2/A2/A2/M2/s1 ),
    .A2(\V3/A2/A2/A2/c1 ),
    .ZN(\V3/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M2/M2/_1_  (.A(\V3/A2/A2/A2/M2/s1 ),
    .B(\V3/A2/A2/A2/c1 ),
    .Z(\V3/s2 [13]));
 OR2_X1 \V3/A2/A2/A2/M2/_0_  (.A1(\V3/A2/A2/A2/M2/c1 ),
    .A2(\V3/A2/A2/A2/M2/c2 ),
    .ZN(\V3/A2/A2/A2/c2 ));
 AND2_X1 \V3/A2/A2/A2/M3/M1/_0_  (.A1(\V3/s1 [14]),
    .A2(ground),
    .ZN(\V3/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M3/M1/_1_  (.A(\V3/s1 [14]),
    .B(ground),
    .Z(\V3/A2/A2/A2/M3/s1 ));
 AND2_X1 \V3/A2/A2/A2/M3/M2/_0_  (.A1(\V3/A2/A2/A2/M3/s1 ),
    .A2(\V3/A2/A2/A2/c2 ),
    .ZN(\V3/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M3/M2/_1_  (.A(\V3/A2/A2/A2/M3/s1 ),
    .B(\V3/A2/A2/A2/c2 ),
    .Z(\V3/s2 [14]));
 OR2_X1 \V3/A2/A2/A2/M3/_0_  (.A1(\V3/A2/A2/A2/M3/c1 ),
    .A2(\V3/A2/A2/A2/M3/c2 ),
    .ZN(\V3/A2/A2/A2/c3 ));
 AND2_X1 \V3/A2/A2/A2/M4/M1/_0_  (.A1(\V3/s1 [15]),
    .A2(ground),
    .ZN(\V3/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M4/M1/_1_  (.A(\V3/s1 [15]),
    .B(ground),
    .Z(\V3/A2/A2/A2/M4/s1 ));
 AND2_X1 \V3/A2/A2/A2/M4/M2/_0_  (.A1(\V3/A2/A2/A2/M4/s1 ),
    .A2(\V3/A2/A2/A2/c3 ),
    .ZN(\V3/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M4/M2/_1_  (.A(\V3/A2/A2/A2/M4/s1 ),
    .B(\V3/A2/A2/A2/c3 ),
    .Z(\V3/s2 [15]));
 OR2_X1 \V3/A2/A2/A2/M4/_0_  (.A1(\V3/A2/A2/A2/M4/c1 ),
    .A2(\V3/A2/A2/A2/M4/c2 ),
    .ZN(\V3/c2 ));
 AND2_X1 \V3/A3/A1/A1/M1/M1/_0_  (.A1(\V3/v4 [0]),
    .A2(\V3/s2 [8]),
    .ZN(\V3/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M1/M1/_1_  (.A(\V3/v4 [0]),
    .B(\V3/s2 [8]),
    .Z(\V3/A3/A1/A1/M1/s1 ));
 AND2_X1 \V3/A3/A1/A1/M1/M2/_0_  (.A1(\V3/A3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M1/M2/_1_  (.A(\V3/A3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v3[16]));
 OR2_X1 \V3/A3/A1/A1/M1/_0_  (.A1(\V3/A3/A1/A1/M1/c1 ),
    .A2(\V3/A3/A1/A1/M1/c2 ),
    .ZN(\V3/A3/A1/A1/c1 ));
 AND2_X1 \V3/A3/A1/A1/M2/M1/_0_  (.A1(\V3/v4 [1]),
    .A2(\V3/s2 [9]),
    .ZN(\V3/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M2/M1/_1_  (.A(\V3/v4 [1]),
    .B(\V3/s2 [9]),
    .Z(\V3/A3/A1/A1/M2/s1 ));
 AND2_X1 \V3/A3/A1/A1/M2/M2/_0_  (.A1(\V3/A3/A1/A1/M2/s1 ),
    .A2(\V3/A3/A1/A1/c1 ),
    .ZN(\V3/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M2/M2/_1_  (.A(\V3/A3/A1/A1/M2/s1 ),
    .B(\V3/A3/A1/A1/c1 ),
    .Z(v3[17]));
 OR2_X1 \V3/A3/A1/A1/M2/_0_  (.A1(\V3/A3/A1/A1/M2/c1 ),
    .A2(\V3/A3/A1/A1/M2/c2 ),
    .ZN(\V3/A3/A1/A1/c2 ));
 AND2_X1 \V3/A3/A1/A1/M3/M1/_0_  (.A1(\V3/v4 [2]),
    .A2(\V3/s2 [10]),
    .ZN(\V3/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M3/M1/_1_  (.A(\V3/v4 [2]),
    .B(\V3/s2 [10]),
    .Z(\V3/A3/A1/A1/M3/s1 ));
 AND2_X1 \V3/A3/A1/A1/M3/M2/_0_  (.A1(\V3/A3/A1/A1/M3/s1 ),
    .A2(\V3/A3/A1/A1/c2 ),
    .ZN(\V3/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M3/M2/_1_  (.A(\V3/A3/A1/A1/M3/s1 ),
    .B(\V3/A3/A1/A1/c2 ),
    .Z(v3[18]));
 OR2_X1 \V3/A3/A1/A1/M3/_0_  (.A1(\V3/A3/A1/A1/M3/c1 ),
    .A2(\V3/A3/A1/A1/M3/c2 ),
    .ZN(\V3/A3/A1/A1/c3 ));
 AND2_X1 \V3/A3/A1/A1/M4/M1/_0_  (.A1(\V3/v4 [3]),
    .A2(\V3/s2 [11]),
    .ZN(\V3/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M4/M1/_1_  (.A(\V3/v4 [3]),
    .B(\V3/s2 [11]),
    .Z(\V3/A3/A1/A1/M4/s1 ));
 AND2_X1 \V3/A3/A1/A1/M4/M2/_0_  (.A1(\V3/A3/A1/A1/M4/s1 ),
    .A2(\V3/A3/A1/A1/c3 ),
    .ZN(\V3/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M4/M2/_1_  (.A(\V3/A3/A1/A1/M4/s1 ),
    .B(\V3/A3/A1/A1/c3 ),
    .Z(v3[19]));
 OR2_X1 \V3/A3/A1/A1/M4/_0_  (.A1(\V3/A3/A1/A1/M4/c1 ),
    .A2(\V3/A3/A1/A1/M4/c2 ),
    .ZN(\V3/A3/A1/c1 ));
 AND2_X1 \V3/A3/A1/A2/M1/M1/_0_  (.A1(\V3/v4 [4]),
    .A2(\V3/s2 [12]),
    .ZN(\V3/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M1/M1/_1_  (.A(\V3/v4 [4]),
    .B(\V3/s2 [12]),
    .Z(\V3/A3/A1/A2/M1/s1 ));
 AND2_X1 \V3/A3/A1/A2/M1/M2/_0_  (.A1(\V3/A3/A1/A2/M1/s1 ),
    .A2(\V3/A3/A1/c1 ),
    .ZN(\V3/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M1/M2/_1_  (.A(\V3/A3/A1/A2/M1/s1 ),
    .B(\V3/A3/A1/c1 ),
    .Z(v3[20]));
 OR2_X1 \V3/A3/A1/A2/M1/_0_  (.A1(\V3/A3/A1/A2/M1/c1 ),
    .A2(\V3/A3/A1/A2/M1/c2 ),
    .ZN(\V3/A3/A1/A2/c1 ));
 AND2_X1 \V3/A3/A1/A2/M2/M1/_0_  (.A1(\V3/v4 [5]),
    .A2(\V3/s2 [13]),
    .ZN(\V3/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M2/M1/_1_  (.A(\V3/v4 [5]),
    .B(\V3/s2 [13]),
    .Z(\V3/A3/A1/A2/M2/s1 ));
 AND2_X1 \V3/A3/A1/A2/M2/M2/_0_  (.A1(\V3/A3/A1/A2/M2/s1 ),
    .A2(\V3/A3/A1/A2/c1 ),
    .ZN(\V3/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M2/M2/_1_  (.A(\V3/A3/A1/A2/M2/s1 ),
    .B(\V3/A3/A1/A2/c1 ),
    .Z(v3[21]));
 OR2_X1 \V3/A3/A1/A2/M2/_0_  (.A1(\V3/A3/A1/A2/M2/c1 ),
    .A2(\V3/A3/A1/A2/M2/c2 ),
    .ZN(\V3/A3/A1/A2/c2 ));
 AND2_X1 \V3/A3/A1/A2/M3/M1/_0_  (.A1(\V3/v4 [6]),
    .A2(\V3/s2 [14]),
    .ZN(\V3/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M3/M1/_1_  (.A(\V3/v4 [6]),
    .B(\V3/s2 [14]),
    .Z(\V3/A3/A1/A2/M3/s1 ));
 AND2_X1 \V3/A3/A1/A2/M3/M2/_0_  (.A1(\V3/A3/A1/A2/M3/s1 ),
    .A2(\V3/A3/A1/A2/c2 ),
    .ZN(\V3/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M3/M2/_1_  (.A(\V3/A3/A1/A2/M3/s1 ),
    .B(\V3/A3/A1/A2/c2 ),
    .Z(v3[22]));
 OR2_X1 \V3/A3/A1/A2/M3/_0_  (.A1(\V3/A3/A1/A2/M3/c1 ),
    .A2(\V3/A3/A1/A2/M3/c2 ),
    .ZN(\V3/A3/A1/A2/c3 ));
 AND2_X1 \V3/A3/A1/A2/M4/M1/_0_  (.A1(\V3/v4 [7]),
    .A2(\V3/s2 [15]),
    .ZN(\V3/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M4/M1/_1_  (.A(\V3/v4 [7]),
    .B(\V3/s2 [15]),
    .Z(\V3/A3/A1/A2/M4/s1 ));
 AND2_X1 \V3/A3/A1/A2/M4/M2/_0_  (.A1(\V3/A3/A1/A2/M4/s1 ),
    .A2(\V3/A3/A1/A2/c3 ),
    .ZN(\V3/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M4/M2/_1_  (.A(\V3/A3/A1/A2/M4/s1 ),
    .B(\V3/A3/A1/A2/c3 ),
    .Z(v3[23]));
 OR2_X1 \V3/A3/A1/A2/M4/_0_  (.A1(\V3/A3/A1/A2/M4/c1 ),
    .A2(\V3/A3/A1/A2/M4/c2 ),
    .ZN(\V3/A3/c1 ));
 AND2_X1 \V3/A3/A2/A1/M1/M1/_0_  (.A1(\V3/v4 [8]),
    .A2(\V3/c3 ),
    .ZN(\V3/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M1/M1/_1_  (.A(\V3/v4 [8]),
    .B(\V3/c3 ),
    .Z(\V3/A3/A2/A1/M1/s1 ));
 AND2_X1 \V3/A3/A2/A1/M1/M2/_0_  (.A1(\V3/A3/A2/A1/M1/s1 ),
    .A2(\V3/A3/c1 ),
    .ZN(\V3/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M1/M2/_1_  (.A(\V3/A3/A2/A1/M1/s1 ),
    .B(\V3/A3/c1 ),
    .Z(v3[24]));
 OR2_X1 \V3/A3/A2/A1/M1/_0_  (.A1(\V3/A3/A2/A1/M1/c1 ),
    .A2(\V3/A3/A2/A1/M1/c2 ),
    .ZN(\V3/A3/A2/A1/c1 ));
 AND2_X1 \V3/A3/A2/A1/M2/M1/_0_  (.A1(\V3/v4 [9]),
    .A2(ground),
    .ZN(\V3/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M2/M1/_1_  (.A(\V3/v4 [9]),
    .B(ground),
    .Z(\V3/A3/A2/A1/M2/s1 ));
 AND2_X1 \V3/A3/A2/A1/M2/M2/_0_  (.A1(\V3/A3/A2/A1/M2/s1 ),
    .A2(\V3/A3/A2/A1/c1 ),
    .ZN(\V3/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M2/M2/_1_  (.A(\V3/A3/A2/A1/M2/s1 ),
    .B(\V3/A3/A2/A1/c1 ),
    .Z(v3[25]));
 OR2_X1 \V3/A3/A2/A1/M2/_0_  (.A1(\V3/A3/A2/A1/M2/c1 ),
    .A2(\V3/A3/A2/A1/M2/c2 ),
    .ZN(\V3/A3/A2/A1/c2 ));
 AND2_X1 \V3/A3/A2/A1/M3/M1/_0_  (.A1(\V3/v4 [10]),
    .A2(ground),
    .ZN(\V3/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M3/M1/_1_  (.A(\V3/v4 [10]),
    .B(ground),
    .Z(\V3/A3/A2/A1/M3/s1 ));
 AND2_X1 \V3/A3/A2/A1/M3/M2/_0_  (.A1(\V3/A3/A2/A1/M3/s1 ),
    .A2(\V3/A3/A2/A1/c2 ),
    .ZN(\V3/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M3/M2/_1_  (.A(\V3/A3/A2/A1/M3/s1 ),
    .B(\V3/A3/A2/A1/c2 ),
    .Z(v3[26]));
 OR2_X1 \V3/A3/A2/A1/M3/_0_  (.A1(\V3/A3/A2/A1/M3/c1 ),
    .A2(\V3/A3/A2/A1/M3/c2 ),
    .ZN(\V3/A3/A2/A1/c3 ));
 AND2_X1 \V3/A3/A2/A1/M4/M1/_0_  (.A1(\V3/v4 [11]),
    .A2(ground),
    .ZN(\V3/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M4/M1/_1_  (.A(\V3/v4 [11]),
    .B(ground),
    .Z(\V3/A3/A2/A1/M4/s1 ));
 AND2_X1 \V3/A3/A2/A1/M4/M2/_0_  (.A1(\V3/A3/A2/A1/M4/s1 ),
    .A2(\V3/A3/A2/A1/c3 ),
    .ZN(\V3/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M4/M2/_1_  (.A(\V3/A3/A2/A1/M4/s1 ),
    .B(\V3/A3/A2/A1/c3 ),
    .Z(v3[27]));
 OR2_X1 \V3/A3/A2/A1/M4/_0_  (.A1(\V3/A3/A2/A1/M4/c1 ),
    .A2(\V3/A3/A2/A1/M4/c2 ),
    .ZN(\V3/A3/A2/c1 ));
 AND2_X1 \V3/A3/A2/A2/M1/M1/_0_  (.A1(\V3/v4 [12]),
    .A2(ground),
    .ZN(\V3/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M1/M1/_1_  (.A(\V3/v4 [12]),
    .B(ground),
    .Z(\V3/A3/A2/A2/M1/s1 ));
 AND2_X1 \V3/A3/A2/A2/M1/M2/_0_  (.A1(\V3/A3/A2/A2/M1/s1 ),
    .A2(\V3/A3/A2/c1 ),
    .ZN(\V3/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M1/M2/_1_  (.A(\V3/A3/A2/A2/M1/s1 ),
    .B(\V3/A3/A2/c1 ),
    .Z(v3[28]));
 OR2_X1 \V3/A3/A2/A2/M1/_0_  (.A1(\V3/A3/A2/A2/M1/c1 ),
    .A2(\V3/A3/A2/A2/M1/c2 ),
    .ZN(\V3/A3/A2/A2/c1 ));
 AND2_X1 \V3/A3/A2/A2/M2/M1/_0_  (.A1(\V3/v4 [13]),
    .A2(ground),
    .ZN(\V3/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M2/M1/_1_  (.A(\V3/v4 [13]),
    .B(ground),
    .Z(\V3/A3/A2/A2/M2/s1 ));
 AND2_X1 \V3/A3/A2/A2/M2/M2/_0_  (.A1(\V3/A3/A2/A2/M2/s1 ),
    .A2(\V3/A3/A2/A2/c1 ),
    .ZN(\V3/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M2/M2/_1_  (.A(\V3/A3/A2/A2/M2/s1 ),
    .B(\V3/A3/A2/A2/c1 ),
    .Z(v3[29]));
 OR2_X1 \V3/A3/A2/A2/M2/_0_  (.A1(\V3/A3/A2/A2/M2/c1 ),
    .A2(\V3/A3/A2/A2/M2/c2 ),
    .ZN(\V3/A3/A2/A2/c2 ));
 AND2_X1 \V3/A3/A2/A2/M3/M1/_0_  (.A1(\V3/v4 [14]),
    .A2(ground),
    .ZN(\V3/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M3/M1/_1_  (.A(\V3/v4 [14]),
    .B(ground),
    .Z(\V3/A3/A2/A2/M3/s1 ));
 AND2_X1 \V3/A3/A2/A2/M3/M2/_0_  (.A1(\V3/A3/A2/A2/M3/s1 ),
    .A2(\V3/A3/A2/A2/c2 ),
    .ZN(\V3/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M3/M2/_1_  (.A(\V3/A3/A2/A2/M3/s1 ),
    .B(\V3/A3/A2/A2/c2 ),
    .Z(v3[30]));
 OR2_X1 \V3/A3/A2/A2/M3/_0_  (.A1(\V3/A3/A2/A2/M3/c1 ),
    .A2(\V3/A3/A2/A2/M3/c2 ),
    .ZN(\V3/A3/A2/A2/c3 ));
 AND2_X1 \V3/A3/A2/A2/M4/M1/_0_  (.A1(\V3/v4 [15]),
    .A2(ground),
    .ZN(\V3/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M4/M1/_1_  (.A(\V3/v4 [15]),
    .B(ground),
    .Z(\V3/A3/A2/A2/M4/s1 ));
 AND2_X1 \V3/A3/A2/A2/M4/M2/_0_  (.A1(\V3/A3/A2/A2/M4/s1 ),
    .A2(\V3/A3/A2/A2/c3 ),
    .ZN(\V3/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M4/M2/_1_  (.A(\V3/A3/A2/A2/M4/s1 ),
    .B(\V3/A3/A2/A2/c3 ),
    .Z(v3[31]));
 OR2_X1 \V3/A3/A2/A2/M4/_0_  (.A1(\V3/A3/A2/A2/M4/c1 ),
    .A2(\V3/A3/A2/A2/M4/c2 ),
    .ZN(\V3/overflow ));
 AND2_X1 \V3/V1/A1/A1/M1/M1/_0_  (.A1(\V3/V1/v2 [0]),
    .A2(\V3/V1/v3 [0]),
    .ZN(\V3/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M1/M1/_1_  (.A(\V3/V1/v2 [0]),
    .B(\V3/V1/v3 [0]),
    .Z(\V3/V1/A1/A1/M1/s1 ));
 AND2_X1 \V3/V1/A1/A1/M1/M2/_0_  (.A1(\V3/V1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M1/M2/_1_  (.A(\V3/V1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/s1 [0]));
 OR2_X2 \V3/V1/A1/A1/M1/_0_  (.A1(\V3/V1/A1/A1/M1/c1 ),
    .A2(\V3/V1/A1/A1/M1/c2 ),
    .ZN(\V3/V1/A1/A1/c1 ));
 AND2_X1 \V3/V1/A1/A1/M2/M1/_0_  (.A1(\V3/V1/v2 [1]),
    .A2(\V3/V1/v3 [1]),
    .ZN(\V3/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M2/M1/_1_  (.A(\V3/V1/v2 [1]),
    .B(\V3/V1/v3 [1]),
    .Z(\V3/V1/A1/A1/M2/s1 ));
 AND2_X1 \V3/V1/A1/A1/M2/M2/_0_  (.A1(\V3/V1/A1/A1/M2/s1 ),
    .A2(\V3/V1/A1/A1/c1 ),
    .ZN(\V3/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M2/M2/_1_  (.A(\V3/V1/A1/A1/M2/s1 ),
    .B(\V3/V1/A1/A1/c1 ),
    .Z(\V3/V1/s1 [1]));
 OR2_X1 \V3/V1/A1/A1/M2/_0_  (.A1(\V3/V1/A1/A1/M2/c1 ),
    .A2(\V3/V1/A1/A1/M2/c2 ),
    .ZN(\V3/V1/A1/A1/c2 ));
 AND2_X1 \V3/V1/A1/A1/M3/M1/_0_  (.A1(\V3/V1/v2 [2]),
    .A2(\V3/V1/v3 [2]),
    .ZN(\V3/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M3/M1/_1_  (.A(\V3/V1/v2 [2]),
    .B(\V3/V1/v3 [2]),
    .Z(\V3/V1/A1/A1/M3/s1 ));
 AND2_X1 \V3/V1/A1/A1/M3/M2/_0_  (.A1(\V3/V1/A1/A1/M3/s1 ),
    .A2(\V3/V1/A1/A1/c2 ),
    .ZN(\V3/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M3/M2/_1_  (.A(\V3/V1/A1/A1/M3/s1 ),
    .B(\V3/V1/A1/A1/c2 ),
    .Z(\V3/V1/s1 [2]));
 OR2_X1 \V3/V1/A1/A1/M3/_0_  (.A1(\V3/V1/A1/A1/M3/c1 ),
    .A2(\V3/V1/A1/A1/M3/c2 ),
    .ZN(\V3/V1/A1/A1/c3 ));
 AND2_X1 \V3/V1/A1/A1/M4/M1/_0_  (.A1(\V3/V1/v2 [3]),
    .A2(\V3/V1/v3 [3]),
    .ZN(\V3/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M4/M1/_1_  (.A(\V3/V1/v2 [3]),
    .B(\V3/V1/v3 [3]),
    .Z(\V3/V1/A1/A1/M4/s1 ));
 AND2_X1 \V3/V1/A1/A1/M4/M2/_0_  (.A1(\V3/V1/A1/A1/M4/s1 ),
    .A2(\V3/V1/A1/A1/c3 ),
    .ZN(\V3/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M4/M2/_1_  (.A(\V3/V1/A1/A1/M4/s1 ),
    .B(\V3/V1/A1/A1/c3 ),
    .Z(\V3/V1/s1 [3]));
 OR2_X1 \V3/V1/A1/A1/M4/_0_  (.A1(\V3/V1/A1/A1/M4/c1 ),
    .A2(\V3/V1/A1/A1/M4/c2 ),
    .ZN(\V3/V1/A1/c1 ));
 AND2_X1 \V3/V1/A1/A2/M1/M1/_0_  (.A1(\V3/V1/v2 [4]),
    .A2(\V3/V1/v3 [4]),
    .ZN(\V3/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M1/M1/_1_  (.A(\V3/V1/v2 [4]),
    .B(\V3/V1/v3 [4]),
    .Z(\V3/V1/A1/A2/M1/s1 ));
 AND2_X1 \V3/V1/A1/A2/M1/M2/_0_  (.A1(\V3/V1/A1/A2/M1/s1 ),
    .A2(\V3/V1/A1/c1 ),
    .ZN(\V3/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M1/M2/_1_  (.A(\V3/V1/A1/A2/M1/s1 ),
    .B(\V3/V1/A1/c1 ),
    .Z(\V3/V1/s1 [4]));
 OR2_X1 \V3/V1/A1/A2/M1/_0_  (.A1(\V3/V1/A1/A2/M1/c1 ),
    .A2(\V3/V1/A1/A2/M1/c2 ),
    .ZN(\V3/V1/A1/A2/c1 ));
 AND2_X1 \V3/V1/A1/A2/M2/M1/_0_  (.A1(\V3/V1/v2 [5]),
    .A2(\V3/V1/v3 [5]),
    .ZN(\V3/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M2/M1/_1_  (.A(\V3/V1/v2 [5]),
    .B(\V3/V1/v3 [5]),
    .Z(\V3/V1/A1/A2/M2/s1 ));
 AND2_X1 \V3/V1/A1/A2/M2/M2/_0_  (.A1(\V3/V1/A1/A2/M2/s1 ),
    .A2(\V3/V1/A1/A2/c1 ),
    .ZN(\V3/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M2/M2/_1_  (.A(\V3/V1/A1/A2/M2/s1 ),
    .B(\V3/V1/A1/A2/c1 ),
    .Z(\V3/V1/s1 [5]));
 OR2_X1 \V3/V1/A1/A2/M2/_0_  (.A1(\V3/V1/A1/A2/M2/c1 ),
    .A2(\V3/V1/A1/A2/M2/c2 ),
    .ZN(\V3/V1/A1/A2/c2 ));
 AND2_X1 \V3/V1/A1/A2/M3/M1/_0_  (.A1(\V3/V1/v2 [6]),
    .A2(\V3/V1/v3 [6]),
    .ZN(\V3/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M3/M1/_1_  (.A(\V3/V1/v2 [6]),
    .B(\V3/V1/v3 [6]),
    .Z(\V3/V1/A1/A2/M3/s1 ));
 AND2_X1 \V3/V1/A1/A2/M3/M2/_0_  (.A1(\V3/V1/A1/A2/M3/s1 ),
    .A2(\V3/V1/A1/A2/c2 ),
    .ZN(\V3/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M3/M2/_1_  (.A(\V3/V1/A1/A2/M3/s1 ),
    .B(\V3/V1/A1/A2/c2 ),
    .Z(\V3/V1/s1 [6]));
 OR2_X1 \V3/V1/A1/A2/M3/_0_  (.A1(\V3/V1/A1/A2/M3/c1 ),
    .A2(\V3/V1/A1/A2/M3/c2 ),
    .ZN(\V3/V1/A1/A2/c3 ));
 AND2_X1 \V3/V1/A1/A2/M4/M1/_0_  (.A1(\V3/V1/v2 [7]),
    .A2(\V3/V1/v3 [7]),
    .ZN(\V3/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M4/M1/_1_  (.A(\V3/V1/v2 [7]),
    .B(\V3/V1/v3 [7]),
    .Z(\V3/V1/A1/A2/M4/s1 ));
 AND2_X1 \V3/V1/A1/A2/M4/M2/_0_  (.A1(\V3/V1/A1/A2/M4/s1 ),
    .A2(\V3/V1/A1/A2/c3 ),
    .ZN(\V3/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M4/M2/_1_  (.A(\V3/V1/A1/A2/M4/s1 ),
    .B(\V3/V1/A1/A2/c3 ),
    .Z(\V3/V1/s1 [7]));
 OR2_X1 \V3/V1/A1/A2/M4/_0_  (.A1(\V3/V1/A1/A2/M4/c1 ),
    .A2(\V3/V1/A1/A2/M4/c2 ),
    .ZN(\V3/V1/c1 ));
 AND2_X1 \V3/V1/A2/A1/M1/M1/_0_  (.A1(\V3/V1/s1 [0]),
    .A2(\V3/V1/v1 [4]),
    .ZN(\V3/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M1/M1/_1_  (.A(\V3/V1/s1 [0]),
    .B(\V3/V1/v1 [4]),
    .Z(\V3/V1/A2/A1/M1/s1 ));
 AND2_X1 \V3/V1/A2/A1/M1/M2/_0_  (.A1(\V3/V1/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M1/M2/_1_  (.A(\V3/V1/A2/A1/M1/s1 ),
    .B(ground),
    .Z(v3[4]));
 OR2_X1 \V3/V1/A2/A1/M1/_0_  (.A1(\V3/V1/A2/A1/M1/c1 ),
    .A2(\V3/V1/A2/A1/M1/c2 ),
    .ZN(\V3/V1/A2/A1/c1 ));
 AND2_X1 \V3/V1/A2/A1/M2/M1/_0_  (.A1(\V3/V1/s1 [1]),
    .A2(\V3/V1/v1 [5]),
    .ZN(\V3/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M2/M1/_1_  (.A(\V3/V1/s1 [1]),
    .B(\V3/V1/v1 [5]),
    .Z(\V3/V1/A2/A1/M2/s1 ));
 AND2_X1 \V3/V1/A2/A1/M2/M2/_0_  (.A1(\V3/V1/A2/A1/M2/s1 ),
    .A2(\V3/V1/A2/A1/c1 ),
    .ZN(\V3/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M2/M2/_1_  (.A(\V3/V1/A2/A1/M2/s1 ),
    .B(\V3/V1/A2/A1/c1 ),
    .Z(v3[5]));
 OR2_X1 \V3/V1/A2/A1/M2/_0_  (.A1(\V3/V1/A2/A1/M2/c1 ),
    .A2(\V3/V1/A2/A1/M2/c2 ),
    .ZN(\V3/V1/A2/A1/c2 ));
 AND2_X1 \V3/V1/A2/A1/M3/M1/_0_  (.A1(\V3/V1/s1 [2]),
    .A2(\V3/V1/v1 [6]),
    .ZN(\V3/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M3/M1/_1_  (.A(\V3/V1/s1 [2]),
    .B(\V3/V1/v1 [6]),
    .Z(\V3/V1/A2/A1/M3/s1 ));
 AND2_X1 \V3/V1/A2/A1/M3/M2/_0_  (.A1(\V3/V1/A2/A1/M3/s1 ),
    .A2(\V3/V1/A2/A1/c2 ),
    .ZN(\V3/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M3/M2/_1_  (.A(\V3/V1/A2/A1/M3/s1 ),
    .B(\V3/V1/A2/A1/c2 ),
    .Z(v3[6]));
 OR2_X1 \V3/V1/A2/A1/M3/_0_  (.A1(\V3/V1/A2/A1/M3/c1 ),
    .A2(\V3/V1/A2/A1/M3/c2 ),
    .ZN(\V3/V1/A2/A1/c3 ));
 AND2_X1 \V3/V1/A2/A1/M4/M1/_0_  (.A1(\V3/V1/s1 [3]),
    .A2(\V3/V1/v1 [7]),
    .ZN(\V3/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M4/M1/_1_  (.A(\V3/V1/s1 [3]),
    .B(\V3/V1/v1 [7]),
    .Z(\V3/V1/A2/A1/M4/s1 ));
 AND2_X1 \V3/V1/A2/A1/M4/M2/_0_  (.A1(\V3/V1/A2/A1/M4/s1 ),
    .A2(\V3/V1/A2/A1/c3 ),
    .ZN(\V3/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M4/M2/_1_  (.A(\V3/V1/A2/A1/M4/s1 ),
    .B(\V3/V1/A2/A1/c3 ),
    .Z(v3[7]));
 OR2_X2 \V3/V1/A2/A1/M4/_0_  (.A1(\V3/V1/A2/A1/M4/c1 ),
    .A2(\V3/V1/A2/A1/M4/c2 ),
    .ZN(\V3/V1/A2/c1 ));
 AND2_X1 \V3/V1/A2/A2/M1/M1/_0_  (.A1(\V3/V1/s1 [4]),
    .A2(ground),
    .ZN(\V3/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M1/M1/_1_  (.A(\V3/V1/s1 [4]),
    .B(ground),
    .Z(\V3/V1/A2/A2/M1/s1 ));
 AND2_X1 \V3/V1/A2/A2/M1/M2/_0_  (.A1(\V3/V1/A2/A2/M1/s1 ),
    .A2(\V3/V1/A2/c1 ),
    .ZN(\V3/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M1/M2/_1_  (.A(\V3/V1/A2/A2/M1/s1 ),
    .B(\V3/V1/A2/c1 ),
    .Z(\V3/V1/s2 [4]));
 OR2_X1 \V3/V1/A2/A2/M1/_0_  (.A1(\V3/V1/A2/A2/M1/c1 ),
    .A2(\V3/V1/A2/A2/M1/c2 ),
    .ZN(\V3/V1/A2/A2/c1 ));
 AND2_X1 \V3/V1/A2/A2/M2/M1/_0_  (.A1(\V3/V1/s1 [5]),
    .A2(ground),
    .ZN(\V3/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M2/M1/_1_  (.A(\V3/V1/s1 [5]),
    .B(ground),
    .Z(\V3/V1/A2/A2/M2/s1 ));
 AND2_X1 \V3/V1/A2/A2/M2/M2/_0_  (.A1(\V3/V1/A2/A2/M2/s1 ),
    .A2(\V3/V1/A2/A2/c1 ),
    .ZN(\V3/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M2/M2/_1_  (.A(\V3/V1/A2/A2/M2/s1 ),
    .B(\V3/V1/A2/A2/c1 ),
    .Z(\V3/V1/s2 [5]));
 OR2_X1 \V3/V1/A2/A2/M2/_0_  (.A1(\V3/V1/A2/A2/M2/c1 ),
    .A2(\V3/V1/A2/A2/M2/c2 ),
    .ZN(\V3/V1/A2/A2/c2 ));
 AND2_X1 \V3/V1/A2/A2/M3/M1/_0_  (.A1(\V3/V1/s1 [6]),
    .A2(ground),
    .ZN(\V3/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M3/M1/_1_  (.A(\V3/V1/s1 [6]),
    .B(ground),
    .Z(\V3/V1/A2/A2/M3/s1 ));
 AND2_X1 \V3/V1/A2/A2/M3/M2/_0_  (.A1(\V3/V1/A2/A2/M3/s1 ),
    .A2(\V3/V1/A2/A2/c2 ),
    .ZN(\V3/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M3/M2/_1_  (.A(\V3/V1/A2/A2/M3/s1 ),
    .B(\V3/V1/A2/A2/c2 ),
    .Z(\V3/V1/s2 [6]));
 OR2_X1 \V3/V1/A2/A2/M3/_0_  (.A1(\V3/V1/A2/A2/M3/c1 ),
    .A2(\V3/V1/A2/A2/M3/c2 ),
    .ZN(\V3/V1/A2/A2/c3 ));
 AND2_X1 \V3/V1/A2/A2/M4/M1/_0_  (.A1(\V3/V1/s1 [7]),
    .A2(ground),
    .ZN(\V3/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M4/M1/_1_  (.A(\V3/V1/s1 [7]),
    .B(ground),
    .Z(\V3/V1/A2/A2/M4/s1 ));
 AND2_X1 \V3/V1/A2/A2/M4/M2/_0_  (.A1(\V3/V1/A2/A2/M4/s1 ),
    .A2(\V3/V1/A2/A2/c3 ),
    .ZN(\V3/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M4/M2/_1_  (.A(\V3/V1/A2/A2/M4/s1 ),
    .B(\V3/V1/A2/A2/c3 ),
    .Z(\V3/V1/s2 [7]));
 OR2_X1 \V3/V1/A2/A2/M4/_0_  (.A1(\V3/V1/A2/A2/M4/c1 ),
    .A2(\V3/V1/A2/A2/M4/c2 ),
    .ZN(\V3/V1/c2 ));
 AND2_X1 \V3/V1/A3/A1/M1/M1/_0_  (.A1(\V3/V1/v4 [0]),
    .A2(\V3/V1/s2 [4]),
    .ZN(\V3/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M1/M1/_1_  (.A(\V3/V1/v4 [0]),
    .B(\V3/V1/s2 [4]),
    .Z(\V3/V1/A3/A1/M1/s1 ));
 AND2_X1 \V3/V1/A3/A1/M1/M2/_0_  (.A1(\V3/V1/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M1/M2/_1_  (.A(\V3/V1/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v1 [8]));
 OR2_X1 \V3/V1/A3/A1/M1/_0_  (.A1(\V3/V1/A3/A1/M1/c1 ),
    .A2(\V3/V1/A3/A1/M1/c2 ),
    .ZN(\V3/V1/A3/A1/c1 ));
 AND2_X1 \V3/V1/A3/A1/M2/M1/_0_  (.A1(\V3/V1/v4 [1]),
    .A2(\V3/V1/s2 [5]),
    .ZN(\V3/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M2/M1/_1_  (.A(\V3/V1/v4 [1]),
    .B(\V3/V1/s2 [5]),
    .Z(\V3/V1/A3/A1/M2/s1 ));
 AND2_X1 \V3/V1/A3/A1/M2/M2/_0_  (.A1(\V3/V1/A3/A1/M2/s1 ),
    .A2(\V3/V1/A3/A1/c1 ),
    .ZN(\V3/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M2/M2/_1_  (.A(\V3/V1/A3/A1/M2/s1 ),
    .B(\V3/V1/A3/A1/c1 ),
    .Z(\V3/v1 [9]));
 OR2_X1 \V3/V1/A3/A1/M2/_0_  (.A1(\V3/V1/A3/A1/M2/c1 ),
    .A2(\V3/V1/A3/A1/M2/c2 ),
    .ZN(\V3/V1/A3/A1/c2 ));
 AND2_X1 \V3/V1/A3/A1/M3/M1/_0_  (.A1(\V3/V1/v4 [2]),
    .A2(\V3/V1/s2 [6]),
    .ZN(\V3/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M3/M1/_1_  (.A(\V3/V1/v4 [2]),
    .B(\V3/V1/s2 [6]),
    .Z(\V3/V1/A3/A1/M3/s1 ));
 AND2_X1 \V3/V1/A3/A1/M3/M2/_0_  (.A1(\V3/V1/A3/A1/M3/s1 ),
    .A2(\V3/V1/A3/A1/c2 ),
    .ZN(\V3/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M3/M2/_1_  (.A(\V3/V1/A3/A1/M3/s1 ),
    .B(\V3/V1/A3/A1/c2 ),
    .Z(\V3/v1 [10]));
 OR2_X1 \V3/V1/A3/A1/M3/_0_  (.A1(\V3/V1/A3/A1/M3/c1 ),
    .A2(\V3/V1/A3/A1/M3/c2 ),
    .ZN(\V3/V1/A3/A1/c3 ));
 AND2_X1 \V3/V1/A3/A1/M4/M1/_0_  (.A1(\V3/V1/v4 [3]),
    .A2(\V3/V1/s2 [7]),
    .ZN(\V3/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M4/M1/_1_  (.A(\V3/V1/v4 [3]),
    .B(\V3/V1/s2 [7]),
    .Z(\V3/V1/A3/A1/M4/s1 ));
 AND2_X1 \V3/V1/A3/A1/M4/M2/_0_  (.A1(\V3/V1/A3/A1/M4/s1 ),
    .A2(\V3/V1/A3/A1/c3 ),
    .ZN(\V3/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M4/M2/_1_  (.A(\V3/V1/A3/A1/M4/s1 ),
    .B(\V3/V1/A3/A1/c3 ),
    .Z(\V3/v1 [11]));
 OR2_X1 \V3/V1/A3/A1/M4/_0_  (.A1(\V3/V1/A3/A1/M4/c1 ),
    .A2(\V3/V1/A3/A1/M4/c2 ),
    .ZN(\V3/V1/A3/c1 ));
 AND2_X1 \V3/V1/A3/A2/M1/M1/_0_  (.A1(\V3/V1/v4 [4]),
    .A2(\V3/V1/c3 ),
    .ZN(\V3/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M1/M1/_1_  (.A(\V3/V1/v4 [4]),
    .B(\V3/V1/c3 ),
    .Z(\V3/V1/A3/A2/M1/s1 ));
 AND2_X1 \V3/V1/A3/A2/M1/M2/_0_  (.A1(\V3/V1/A3/A2/M1/s1 ),
    .A2(\V3/V1/A3/c1 ),
    .ZN(\V3/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M1/M2/_1_  (.A(\V3/V1/A3/A2/M1/s1 ),
    .B(\V3/V1/A3/c1 ),
    .Z(\V3/v1 [12]));
 OR2_X1 \V3/V1/A3/A2/M1/_0_  (.A1(\V3/V1/A3/A2/M1/c1 ),
    .A2(\V3/V1/A3/A2/M1/c2 ),
    .ZN(\V3/V1/A3/A2/c1 ));
 AND2_X1 \V3/V1/A3/A2/M2/M1/_0_  (.A1(\V3/V1/v4 [5]),
    .A2(ground),
    .ZN(\V3/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M2/M1/_1_  (.A(\V3/V1/v4 [5]),
    .B(ground),
    .Z(\V3/V1/A3/A2/M2/s1 ));
 AND2_X1 \V3/V1/A3/A2/M2/M2/_0_  (.A1(\V3/V1/A3/A2/M2/s1 ),
    .A2(\V3/V1/A3/A2/c1 ),
    .ZN(\V3/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M2/M2/_1_  (.A(\V3/V1/A3/A2/M2/s1 ),
    .B(\V3/V1/A3/A2/c1 ),
    .Z(\V3/v1 [13]));
 OR2_X1 \V3/V1/A3/A2/M2/_0_  (.A1(\V3/V1/A3/A2/M2/c1 ),
    .A2(\V3/V1/A3/A2/M2/c2 ),
    .ZN(\V3/V1/A3/A2/c2 ));
 AND2_X1 \V3/V1/A3/A2/M3/M1/_0_  (.A1(\V3/V1/v4 [6]),
    .A2(ground),
    .ZN(\V3/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M3/M1/_1_  (.A(\V3/V1/v4 [6]),
    .B(ground),
    .Z(\V3/V1/A3/A2/M3/s1 ));
 AND2_X1 \V3/V1/A3/A2/M3/M2/_0_  (.A1(\V3/V1/A3/A2/M3/s1 ),
    .A2(\V3/V1/A3/A2/c2 ),
    .ZN(\V3/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M3/M2/_1_  (.A(\V3/V1/A3/A2/M3/s1 ),
    .B(\V3/V1/A3/A2/c2 ),
    .Z(\V3/v1 [14]));
 OR2_X1 \V3/V1/A3/A2/M3/_0_  (.A1(\V3/V1/A3/A2/M3/c1 ),
    .A2(\V3/V1/A3/A2/M3/c2 ),
    .ZN(\V3/V1/A3/A2/c3 ));
 AND2_X1 \V3/V1/A3/A2/M4/M1/_0_  (.A1(\V3/V1/v4 [7]),
    .A2(ground),
    .ZN(\V3/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M4/M1/_1_  (.A(\V3/V1/v4 [7]),
    .B(ground),
    .Z(\V3/V1/A3/A2/M4/s1 ));
 AND2_X1 \V3/V1/A3/A2/M4/M2/_0_  (.A1(\V3/V1/A3/A2/M4/s1 ),
    .A2(\V3/V1/A3/A2/c3 ),
    .ZN(\V3/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M4/M2/_1_  (.A(\V3/V1/A3/A2/M4/s1 ),
    .B(\V3/V1/A3/A2/c3 ),
    .Z(\V3/v1 [15]));
 OR2_X1 \V3/V1/A3/A2/M4/_0_  (.A1(\V3/V1/A3/A2/M4/c1 ),
    .A2(\V3/V1/A3/A2/M4/c2 ),
    .ZN(\V3/V1/overflow ));
 AND2_X1 \V3/V1/V1/A1/M1/M1/_0_  (.A1(\V3/V1/V1/v2 [0]),
    .A2(\V3/V1/V1/v3 [0]),
    .ZN(\V3/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M1/M1/_1_  (.A(\V3/V1/V1/v2 [0]),
    .B(\V3/V1/V1/v3 [0]),
    .Z(\V3/V1/V1/A1/M1/s1 ));
 AND2_X1 \V3/V1/V1/A1/M1/M2/_0_  (.A1(\V3/V1/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M1/M2/_1_  (.A(\V3/V1/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/V1/s1 [0]));
 OR2_X1 \V3/V1/V1/A1/M1/_0_  (.A1(\V3/V1/V1/A1/M1/c1 ),
    .A2(\V3/V1/V1/A1/M1/c2 ),
    .ZN(\V3/V1/V1/A1/c1 ));
 AND2_X1 \V3/V1/V1/A1/M2/M1/_0_  (.A1(\V3/V1/V1/v2 [1]),
    .A2(\V3/V1/V1/v3 [1]),
    .ZN(\V3/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M2/M1/_1_  (.A(\V3/V1/V1/v2 [1]),
    .B(\V3/V1/V1/v3 [1]),
    .Z(\V3/V1/V1/A1/M2/s1 ));
 AND2_X1 \V3/V1/V1/A1/M2/M2/_0_  (.A1(\V3/V1/V1/A1/M2/s1 ),
    .A2(\V3/V1/V1/A1/c1 ),
    .ZN(\V3/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M2/M2/_1_  (.A(\V3/V1/V1/A1/M2/s1 ),
    .B(\V3/V1/V1/A1/c1 ),
    .Z(\V3/V1/V1/s1 [1]));
 OR2_X1 \V3/V1/V1/A1/M2/_0_  (.A1(\V3/V1/V1/A1/M2/c1 ),
    .A2(\V3/V1/V1/A1/M2/c2 ),
    .ZN(\V3/V1/V1/A1/c2 ));
 AND2_X1 \V3/V1/V1/A1/M3/M1/_0_  (.A1(\V3/V1/V1/v2 [2]),
    .A2(\V3/V1/V1/v3 [2]),
    .ZN(\V3/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M3/M1/_1_  (.A(\V3/V1/V1/v2 [2]),
    .B(\V3/V1/V1/v3 [2]),
    .Z(\V3/V1/V1/A1/M3/s1 ));
 AND2_X1 \V3/V1/V1/A1/M3/M2/_0_  (.A1(\V3/V1/V1/A1/M3/s1 ),
    .A2(\V3/V1/V1/A1/c2 ),
    .ZN(\V3/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M3/M2/_1_  (.A(\V3/V1/V1/A1/M3/s1 ),
    .B(\V3/V1/V1/A1/c2 ),
    .Z(\V3/V1/V1/s1 [2]));
 OR2_X1 \V3/V1/V1/A1/M3/_0_  (.A1(\V3/V1/V1/A1/M3/c1 ),
    .A2(\V3/V1/V1/A1/M3/c2 ),
    .ZN(\V3/V1/V1/A1/c3 ));
 AND2_X1 \V3/V1/V1/A1/M4/M1/_0_  (.A1(\V3/V1/V1/v2 [3]),
    .A2(\V3/V1/V1/v3 [3]),
    .ZN(\V3/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M4/M1/_1_  (.A(\V3/V1/V1/v2 [3]),
    .B(\V3/V1/V1/v3 [3]),
    .Z(\V3/V1/V1/A1/M4/s1 ));
 AND2_X1 \V3/V1/V1/A1/M4/M2/_0_  (.A1(\V3/V1/V1/A1/M4/s1 ),
    .A2(\V3/V1/V1/A1/c3 ),
    .ZN(\V3/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M4/M2/_1_  (.A(\V3/V1/V1/A1/M4/s1 ),
    .B(\V3/V1/V1/A1/c3 ),
    .Z(\V3/V1/V1/s1 [3]));
 OR2_X1 \V3/V1/V1/A1/M4/_0_  (.A1(\V3/V1/V1/A1/M4/c1 ),
    .A2(\V3/V1/V1/A1/M4/c2 ),
    .ZN(\V3/V1/V1/c1 ));
 AND2_X1 \V3/V1/V1/A2/M1/M1/_0_  (.A1(\V3/V1/V1/s1 [0]),
    .A2(\V3/V1/V1/v1 [2]),
    .ZN(\V3/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M1/M1/_1_  (.A(\V3/V1/V1/s1 [0]),
    .B(\V3/V1/V1/v1 [2]),
    .Z(\V3/V1/V1/A2/M1/s1 ));
 AND2_X1 \V3/V1/V1/A2/M1/M2/_0_  (.A1(\V3/V1/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M1/M2/_1_  (.A(\V3/V1/V1/A2/M1/s1 ),
    .B(ground),
    .Z(v3[2]));
 OR2_X1 \V3/V1/V1/A2/M1/_0_  (.A1(\V3/V1/V1/A2/M1/c1 ),
    .A2(\V3/V1/V1/A2/M1/c2 ),
    .ZN(\V3/V1/V1/A2/c1 ));
 AND2_X1 \V3/V1/V1/A2/M2/M1/_0_  (.A1(\V3/V1/V1/s1 [1]),
    .A2(\V3/V1/V1/v1 [3]),
    .ZN(\V3/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M2/M1/_1_  (.A(\V3/V1/V1/s1 [1]),
    .B(\V3/V1/V1/v1 [3]),
    .Z(\V3/V1/V1/A2/M2/s1 ));
 AND2_X1 \V3/V1/V1/A2/M2/M2/_0_  (.A1(\V3/V1/V1/A2/M2/s1 ),
    .A2(\V3/V1/V1/A2/c1 ),
    .ZN(\V3/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M2/M2/_1_  (.A(\V3/V1/V1/A2/M2/s1 ),
    .B(\V3/V1/V1/A2/c1 ),
    .Z(v3[3]));
 OR2_X1 \V3/V1/V1/A2/M2/_0_  (.A1(\V3/V1/V1/A2/M2/c1 ),
    .A2(\V3/V1/V1/A2/M2/c2 ),
    .ZN(\V3/V1/V1/A2/c2 ));
 AND2_X1 \V3/V1/V1/A2/M3/M1/_0_  (.A1(\V3/V1/V1/s1 [2]),
    .A2(ground),
    .ZN(\V3/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M3/M1/_1_  (.A(\V3/V1/V1/s1 [2]),
    .B(ground),
    .Z(\V3/V1/V1/A2/M3/s1 ));
 AND2_X1 \V3/V1/V1/A2/M3/M2/_0_  (.A1(\V3/V1/V1/A2/M3/s1 ),
    .A2(\V3/V1/V1/A2/c2 ),
    .ZN(\V3/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M3/M2/_1_  (.A(\V3/V1/V1/A2/M3/s1 ),
    .B(\V3/V1/V1/A2/c2 ),
    .Z(\V3/V1/V1/s2 [2]));
 OR2_X1 \V3/V1/V1/A2/M3/_0_  (.A1(\V3/V1/V1/A2/M3/c1 ),
    .A2(\V3/V1/V1/A2/M3/c2 ),
    .ZN(\V3/V1/V1/A2/c3 ));
 AND2_X1 \V3/V1/V1/A2/M4/M1/_0_  (.A1(\V3/V1/V1/s1 [3]),
    .A2(ground),
    .ZN(\V3/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M4/M1/_1_  (.A(\V3/V1/V1/s1 [3]),
    .B(ground),
    .Z(\V3/V1/V1/A2/M4/s1 ));
 AND2_X1 \V3/V1/V1/A2/M4/M2/_0_  (.A1(\V3/V1/V1/A2/M4/s1 ),
    .A2(\V3/V1/V1/A2/c3 ),
    .ZN(\V3/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M4/M2/_1_  (.A(\V3/V1/V1/A2/M4/s1 ),
    .B(\V3/V1/V1/A2/c3 ),
    .Z(\V3/V1/V1/s2 [3]));
 OR2_X1 \V3/V1/V1/A2/M4/_0_  (.A1(\V3/V1/V1/A2/M4/c1 ),
    .A2(\V3/V1/V1/A2/M4/c2 ),
    .ZN(\V3/V1/V1/c2 ));
 AND2_X1 \V3/V1/V1/A3/M1/M1/_0_  (.A1(\V3/V1/V1/v4 [0]),
    .A2(\V3/V1/V1/s2 [2]),
    .ZN(\V3/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M1/M1/_1_  (.A(\V3/V1/V1/v4 [0]),
    .B(\V3/V1/V1/s2 [2]),
    .Z(\V3/V1/V1/A3/M1/s1 ));
 AND2_X1 \V3/V1/V1/A3/M1/M2/_0_  (.A1(\V3/V1/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M1/M2/_1_  (.A(\V3/V1/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v1 [4]));
 OR2_X1 \V3/V1/V1/A3/M1/_0_  (.A1(\V3/V1/V1/A3/M1/c1 ),
    .A2(\V3/V1/V1/A3/M1/c2 ),
    .ZN(\V3/V1/V1/A3/c1 ));
 AND2_X1 \V3/V1/V1/A3/M2/M1/_0_  (.A1(\V3/V1/V1/v4 [1]),
    .A2(\V3/V1/V1/s2 [3]),
    .ZN(\V3/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M2/M1/_1_  (.A(\V3/V1/V1/v4 [1]),
    .B(\V3/V1/V1/s2 [3]),
    .Z(\V3/V1/V1/A3/M2/s1 ));
 AND2_X1 \V3/V1/V1/A3/M2/M2/_0_  (.A1(\V3/V1/V1/A3/M2/s1 ),
    .A2(\V3/V1/V1/A3/c1 ),
    .ZN(\V3/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M2/M2/_1_  (.A(\V3/V1/V1/A3/M2/s1 ),
    .B(\V3/V1/V1/A3/c1 ),
    .Z(\V3/V1/v1 [5]));
 OR2_X1 \V3/V1/V1/A3/M2/_0_  (.A1(\V3/V1/V1/A3/M2/c1 ),
    .A2(\V3/V1/V1/A3/M2/c2 ),
    .ZN(\V3/V1/V1/A3/c2 ));
 AND2_X1 \V3/V1/V1/A3/M3/M1/_0_  (.A1(\V3/V1/V1/v4 [2]),
    .A2(\V3/V1/V1/c3 ),
    .ZN(\V3/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M3/M1/_1_  (.A(\V3/V1/V1/v4 [2]),
    .B(\V3/V1/V1/c3 ),
    .Z(\V3/V1/V1/A3/M3/s1 ));
 AND2_X1 \V3/V1/V1/A3/M3/M2/_0_  (.A1(\V3/V1/V1/A3/M3/s1 ),
    .A2(\V3/V1/V1/A3/c2 ),
    .ZN(\V3/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M3/M2/_1_  (.A(\V3/V1/V1/A3/M3/s1 ),
    .B(\V3/V1/V1/A3/c2 ),
    .Z(\V3/V1/v1 [6]));
 OR2_X1 \V3/V1/V1/A3/M3/_0_  (.A1(\V3/V1/V1/A3/M3/c1 ),
    .A2(\V3/V1/V1/A3/M3/c2 ),
    .ZN(\V3/V1/V1/A3/c3 ));
 AND2_X1 \V3/V1/V1/A3/M4/M1/_0_  (.A1(\V3/V1/V1/v4 [3]),
    .A2(ground),
    .ZN(\V3/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M4/M1/_1_  (.A(\V3/V1/V1/v4 [3]),
    .B(ground),
    .Z(\V3/V1/V1/A3/M4/s1 ));
 AND2_X1 \V3/V1/V1/A3/M4/M2/_0_  (.A1(\V3/V1/V1/A3/M4/s1 ),
    .A2(\V3/V1/V1/A3/c3 ),
    .ZN(\V3/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M4/M2/_1_  (.A(\V3/V1/V1/A3/M4/s1 ),
    .B(\V3/V1/V1/A3/c3 ),
    .Z(\V3/V1/v1 [7]));
 OR2_X1 \V3/V1/V1/A3/M4/_0_  (.A1(\V3/V1/V1/A3/M4/c1 ),
    .A2(\V3/V1/V1/A3/M4/c2 ),
    .ZN(\V3/V1/V1/overflow ));
 AND2_X1 \V3/V1/V1/V1/HA1/_0_  (.A1(\V3/V1/V1/V1/w2 ),
    .A2(\V3/V1/V1/V1/w1 ),
    .ZN(\V3/V1/V1/V1/w4 ));
 XOR2_X2 \V3/V1/V1/V1/HA1/_1_  (.A(\V3/V1/V1/V1/w2 ),
    .B(\V3/V1/V1/V1/w1 ),
    .Z(v3[1]));
 AND2_X1 \V3/V1/V1/V1/HA2/_0_  (.A1(\V3/V1/V1/V1/w4 ),
    .A2(\V3/V1/V1/V1/w3 ),
    .ZN(\V3/V1/V1/v1 [3]));
 XOR2_X2 \V3/V1/V1/V1/HA2/_1_  (.A(\V3/V1/V1/V1/w4 ),
    .B(\V3/V1/V1/V1/w3 ),
    .Z(\V3/V1/V1/v1 [2]));
 AND2_X1 \V3/V1/V1/V1/_0_  (.A1(A[0]),
    .A2(B[16]),
    .ZN(v3[0]));
 AND2_X1 \V3/V1/V1/V1/_1_  (.A1(A[0]),
    .A2(B[17]),
    .ZN(\V3/V1/V1/V1/w1 ));
 AND2_X1 \V3/V1/V1/V1/_2_  (.A1(B[16]),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V1/w2 ));
 AND2_X1 \V3/V1/V1/V1/_3_  (.A1(B[17]),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V1/w3 ));
 AND2_X1 \V3/V1/V1/V2/HA1/_0_  (.A1(\V3/V1/V1/V2/w2 ),
    .A2(\V3/V1/V1/V2/w1 ),
    .ZN(\V3/V1/V1/V2/w4 ));
 XOR2_X2 \V3/V1/V1/V2/HA1/_1_  (.A(\V3/V1/V1/V2/w2 ),
    .B(\V3/V1/V1/V2/w1 ),
    .Z(\V3/V1/V1/v2 [1]));
 AND2_X1 \V3/V1/V1/V2/HA2/_0_  (.A1(\V3/V1/V1/V2/w4 ),
    .A2(\V3/V1/V1/V2/w3 ),
    .ZN(\V3/V1/V1/v2 [3]));
 XOR2_X2 \V3/V1/V1/V2/HA2/_1_  (.A(\V3/V1/V1/V2/w4 ),
    .B(\V3/V1/V1/V2/w3 ),
    .Z(\V3/V1/V1/v2 [2]));
 AND2_X1 \V3/V1/V1/V2/_0_  (.A1(A[2]),
    .A2(B[16]),
    .ZN(\V3/V1/V1/v2 [0]));
 AND2_X1 \V3/V1/V1/V2/_1_  (.A1(A[2]),
    .A2(B[17]),
    .ZN(\V3/V1/V1/V2/w1 ));
 AND2_X1 \V3/V1/V1/V2/_2_  (.A1(B[16]),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V2/w2 ));
 AND2_X1 \V3/V1/V1/V2/_3_  (.A1(B[17]),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V2/w3 ));
 AND2_X1 \V3/V1/V1/V3/HA1/_0_  (.A1(\V3/V1/V1/V3/w2 ),
    .A2(\V3/V1/V1/V3/w1 ),
    .ZN(\V3/V1/V1/V3/w4 ));
 XOR2_X2 \V3/V1/V1/V3/HA1/_1_  (.A(\V3/V1/V1/V3/w2 ),
    .B(\V3/V1/V1/V3/w1 ),
    .Z(\V3/V1/V1/v3 [1]));
 AND2_X1 \V3/V1/V1/V3/HA2/_0_  (.A1(\V3/V1/V1/V3/w4 ),
    .A2(\V3/V1/V1/V3/w3 ),
    .ZN(\V3/V1/V1/v3 [3]));
 XOR2_X2 \V3/V1/V1/V3/HA2/_1_  (.A(\V3/V1/V1/V3/w4 ),
    .B(\V3/V1/V1/V3/w3 ),
    .Z(\V3/V1/V1/v3 [2]));
 AND2_X1 \V3/V1/V1/V3/_0_  (.A1(A[0]),
    .A2(B[18]),
    .ZN(\V3/V1/V1/v3 [0]));
 AND2_X1 \V3/V1/V1/V3/_1_  (.A1(A[0]),
    .A2(B[19]),
    .ZN(\V3/V1/V1/V3/w1 ));
 AND2_X1 \V3/V1/V1/V3/_2_  (.A1(B[18]),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V3/w2 ));
 AND2_X1 \V3/V1/V1/V3/_3_  (.A1(B[19]),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V3/w3 ));
 AND2_X1 \V3/V1/V1/V4/HA1/_0_  (.A1(\V3/V1/V1/V4/w2 ),
    .A2(\V3/V1/V1/V4/w1 ),
    .ZN(\V3/V1/V1/V4/w4 ));
 XOR2_X2 \V3/V1/V1/V4/HA1/_1_  (.A(\V3/V1/V1/V4/w2 ),
    .B(\V3/V1/V1/V4/w1 ),
    .Z(\V3/V1/V1/v4 [1]));
 AND2_X1 \V3/V1/V1/V4/HA2/_0_  (.A1(\V3/V1/V1/V4/w4 ),
    .A2(\V3/V1/V1/V4/w3 ),
    .ZN(\V3/V1/V1/v4 [3]));
 XOR2_X2 \V3/V1/V1/V4/HA2/_1_  (.A(\V3/V1/V1/V4/w4 ),
    .B(\V3/V1/V1/V4/w3 ),
    .Z(\V3/V1/V1/v4 [2]));
 AND2_X1 \V3/V1/V1/V4/_0_  (.A1(A[2]),
    .A2(B[18]),
    .ZN(\V3/V1/V1/v4 [0]));
 AND2_X1 \V3/V1/V1/V4/_1_  (.A1(A[2]),
    .A2(B[19]),
    .ZN(\V3/V1/V1/V4/w1 ));
 AND2_X1 \V3/V1/V1/V4/_2_  (.A1(B[18]),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V4/w2 ));
 AND2_X1 \V3/V1/V1/V4/_3_  (.A1(B[19]),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V4/w3 ));
 OR2_X1 \V3/V1/V1/_0_  (.A1(\V3/V1/V1/c1 ),
    .A2(\V3/V1/V1/c2 ),
    .ZN(\V3/V1/V1/c3 ));
 AND2_X1 \V3/V1/V2/A1/M1/M1/_0_  (.A1(\V3/V1/V2/v2 [0]),
    .A2(\V3/V1/V2/v3 [0]),
    .ZN(\V3/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M1/M1/_1_  (.A(\V3/V1/V2/v2 [0]),
    .B(\V3/V1/V2/v3 [0]),
    .Z(\V3/V1/V2/A1/M1/s1 ));
 AND2_X1 \V3/V1/V2/A1/M1/M2/_0_  (.A1(\V3/V1/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M1/M2/_1_  (.A(\V3/V1/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/V2/s1 [0]));
 OR2_X1 \V3/V1/V2/A1/M1/_0_  (.A1(\V3/V1/V2/A1/M1/c1 ),
    .A2(\V3/V1/V2/A1/M1/c2 ),
    .ZN(\V3/V1/V2/A1/c1 ));
 AND2_X1 \V3/V1/V2/A1/M2/M1/_0_  (.A1(\V3/V1/V2/v2 [1]),
    .A2(\V3/V1/V2/v3 [1]),
    .ZN(\V3/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M2/M1/_1_  (.A(\V3/V1/V2/v2 [1]),
    .B(\V3/V1/V2/v3 [1]),
    .Z(\V3/V1/V2/A1/M2/s1 ));
 AND2_X1 \V3/V1/V2/A1/M2/M2/_0_  (.A1(\V3/V1/V2/A1/M2/s1 ),
    .A2(\V3/V1/V2/A1/c1 ),
    .ZN(\V3/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M2/M2/_1_  (.A(\V3/V1/V2/A1/M2/s1 ),
    .B(\V3/V1/V2/A1/c1 ),
    .Z(\V3/V1/V2/s1 [1]));
 OR2_X1 \V3/V1/V2/A1/M2/_0_  (.A1(\V3/V1/V2/A1/M2/c1 ),
    .A2(\V3/V1/V2/A1/M2/c2 ),
    .ZN(\V3/V1/V2/A1/c2 ));
 AND2_X1 \V3/V1/V2/A1/M3/M1/_0_  (.A1(\V3/V1/V2/v2 [2]),
    .A2(\V3/V1/V2/v3 [2]),
    .ZN(\V3/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M3/M1/_1_  (.A(\V3/V1/V2/v2 [2]),
    .B(\V3/V1/V2/v3 [2]),
    .Z(\V3/V1/V2/A1/M3/s1 ));
 AND2_X1 \V3/V1/V2/A1/M3/M2/_0_  (.A1(\V3/V1/V2/A1/M3/s1 ),
    .A2(\V3/V1/V2/A1/c2 ),
    .ZN(\V3/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M3/M2/_1_  (.A(\V3/V1/V2/A1/M3/s1 ),
    .B(\V3/V1/V2/A1/c2 ),
    .Z(\V3/V1/V2/s1 [2]));
 OR2_X1 \V3/V1/V2/A1/M3/_0_  (.A1(\V3/V1/V2/A1/M3/c1 ),
    .A2(\V3/V1/V2/A1/M3/c2 ),
    .ZN(\V3/V1/V2/A1/c3 ));
 AND2_X1 \V3/V1/V2/A1/M4/M1/_0_  (.A1(\V3/V1/V2/v2 [3]),
    .A2(\V3/V1/V2/v3 [3]),
    .ZN(\V3/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M4/M1/_1_  (.A(\V3/V1/V2/v2 [3]),
    .B(\V3/V1/V2/v3 [3]),
    .Z(\V3/V1/V2/A1/M4/s1 ));
 AND2_X1 \V3/V1/V2/A1/M4/M2/_0_  (.A1(\V3/V1/V2/A1/M4/s1 ),
    .A2(\V3/V1/V2/A1/c3 ),
    .ZN(\V3/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M4/M2/_1_  (.A(\V3/V1/V2/A1/M4/s1 ),
    .B(\V3/V1/V2/A1/c3 ),
    .Z(\V3/V1/V2/s1 [3]));
 OR2_X1 \V3/V1/V2/A1/M4/_0_  (.A1(\V3/V1/V2/A1/M4/c1 ),
    .A2(\V3/V1/V2/A1/M4/c2 ),
    .ZN(\V3/V1/V2/c1 ));
 AND2_X1 \V3/V1/V2/A2/M1/M1/_0_  (.A1(\V3/V1/V2/s1 [0]),
    .A2(\V3/V1/V2/v1 [2]),
    .ZN(\V3/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M1/M1/_1_  (.A(\V3/V1/V2/s1 [0]),
    .B(\V3/V1/V2/v1 [2]),
    .Z(\V3/V1/V2/A2/M1/s1 ));
 AND2_X1 \V3/V1/V2/A2/M1/M2/_0_  (.A1(\V3/V1/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M1/M2/_1_  (.A(\V3/V1/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v2 [2]));
 OR2_X1 \V3/V1/V2/A2/M1/_0_  (.A1(\V3/V1/V2/A2/M1/c1 ),
    .A2(\V3/V1/V2/A2/M1/c2 ),
    .ZN(\V3/V1/V2/A2/c1 ));
 AND2_X1 \V3/V1/V2/A2/M2/M1/_0_  (.A1(\V3/V1/V2/s1 [1]),
    .A2(\V3/V1/V2/v1 [3]),
    .ZN(\V3/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M2/M1/_1_  (.A(\V3/V1/V2/s1 [1]),
    .B(\V3/V1/V2/v1 [3]),
    .Z(\V3/V1/V2/A2/M2/s1 ));
 AND2_X1 \V3/V1/V2/A2/M2/M2/_0_  (.A1(\V3/V1/V2/A2/M2/s1 ),
    .A2(\V3/V1/V2/A2/c1 ),
    .ZN(\V3/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M2/M2/_1_  (.A(\V3/V1/V2/A2/M2/s1 ),
    .B(\V3/V1/V2/A2/c1 ),
    .Z(\V3/V1/v2 [3]));
 OR2_X1 \V3/V1/V2/A2/M2/_0_  (.A1(\V3/V1/V2/A2/M2/c1 ),
    .A2(\V3/V1/V2/A2/M2/c2 ),
    .ZN(\V3/V1/V2/A2/c2 ));
 AND2_X1 \V3/V1/V2/A2/M3/M1/_0_  (.A1(\V3/V1/V2/s1 [2]),
    .A2(ground),
    .ZN(\V3/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M3/M1/_1_  (.A(\V3/V1/V2/s1 [2]),
    .B(ground),
    .Z(\V3/V1/V2/A2/M3/s1 ));
 AND2_X1 \V3/V1/V2/A2/M3/M2/_0_  (.A1(\V3/V1/V2/A2/M3/s1 ),
    .A2(\V3/V1/V2/A2/c2 ),
    .ZN(\V3/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M3/M2/_1_  (.A(\V3/V1/V2/A2/M3/s1 ),
    .B(\V3/V1/V2/A2/c2 ),
    .Z(\V3/V1/V2/s2 [2]));
 OR2_X1 \V3/V1/V2/A2/M3/_0_  (.A1(\V3/V1/V2/A2/M3/c1 ),
    .A2(\V3/V1/V2/A2/M3/c2 ),
    .ZN(\V3/V1/V2/A2/c3 ));
 AND2_X1 \V3/V1/V2/A2/M4/M1/_0_  (.A1(\V3/V1/V2/s1 [3]),
    .A2(ground),
    .ZN(\V3/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M4/M1/_1_  (.A(\V3/V1/V2/s1 [3]),
    .B(ground),
    .Z(\V3/V1/V2/A2/M4/s1 ));
 AND2_X1 \V3/V1/V2/A2/M4/M2/_0_  (.A1(\V3/V1/V2/A2/M4/s1 ),
    .A2(\V3/V1/V2/A2/c3 ),
    .ZN(\V3/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M4/M2/_1_  (.A(\V3/V1/V2/A2/M4/s1 ),
    .B(\V3/V1/V2/A2/c3 ),
    .Z(\V3/V1/V2/s2 [3]));
 OR2_X1 \V3/V1/V2/A2/M4/_0_  (.A1(\V3/V1/V2/A2/M4/c1 ),
    .A2(\V3/V1/V2/A2/M4/c2 ),
    .ZN(\V3/V1/V2/c2 ));
 AND2_X1 \V3/V1/V2/A3/M1/M1/_0_  (.A1(\V3/V1/V2/v4 [0]),
    .A2(\V3/V1/V2/s2 [2]),
    .ZN(\V3/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M1/M1/_1_  (.A(\V3/V1/V2/v4 [0]),
    .B(\V3/V1/V2/s2 [2]),
    .Z(\V3/V1/V2/A3/M1/s1 ));
 AND2_X1 \V3/V1/V2/A3/M1/M2/_0_  (.A1(\V3/V1/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M1/M2/_1_  (.A(\V3/V1/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v2 [4]));
 OR2_X1 \V3/V1/V2/A3/M1/_0_  (.A1(\V3/V1/V2/A3/M1/c1 ),
    .A2(\V3/V1/V2/A3/M1/c2 ),
    .ZN(\V3/V1/V2/A3/c1 ));
 AND2_X1 \V3/V1/V2/A3/M2/M1/_0_  (.A1(\V3/V1/V2/v4 [1]),
    .A2(\V3/V1/V2/s2 [3]),
    .ZN(\V3/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M2/M1/_1_  (.A(\V3/V1/V2/v4 [1]),
    .B(\V3/V1/V2/s2 [3]),
    .Z(\V3/V1/V2/A3/M2/s1 ));
 AND2_X1 \V3/V1/V2/A3/M2/M2/_0_  (.A1(\V3/V1/V2/A3/M2/s1 ),
    .A2(\V3/V1/V2/A3/c1 ),
    .ZN(\V3/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M2/M2/_1_  (.A(\V3/V1/V2/A3/M2/s1 ),
    .B(\V3/V1/V2/A3/c1 ),
    .Z(\V3/V1/v2 [5]));
 OR2_X1 \V3/V1/V2/A3/M2/_0_  (.A1(\V3/V1/V2/A3/M2/c1 ),
    .A2(\V3/V1/V2/A3/M2/c2 ),
    .ZN(\V3/V1/V2/A3/c2 ));
 AND2_X1 \V3/V1/V2/A3/M3/M1/_0_  (.A1(\V3/V1/V2/v4 [2]),
    .A2(\V3/V1/V2/c3 ),
    .ZN(\V3/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M3/M1/_1_  (.A(\V3/V1/V2/v4 [2]),
    .B(\V3/V1/V2/c3 ),
    .Z(\V3/V1/V2/A3/M3/s1 ));
 AND2_X1 \V3/V1/V2/A3/M3/M2/_0_  (.A1(\V3/V1/V2/A3/M3/s1 ),
    .A2(\V3/V1/V2/A3/c2 ),
    .ZN(\V3/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M3/M2/_1_  (.A(\V3/V1/V2/A3/M3/s1 ),
    .B(\V3/V1/V2/A3/c2 ),
    .Z(\V3/V1/v2 [6]));
 OR2_X1 \V3/V1/V2/A3/M3/_0_  (.A1(\V3/V1/V2/A3/M3/c1 ),
    .A2(\V3/V1/V2/A3/M3/c2 ),
    .ZN(\V3/V1/V2/A3/c3 ));
 AND2_X1 \V3/V1/V2/A3/M4/M1/_0_  (.A1(\V3/V1/V2/v4 [3]),
    .A2(ground),
    .ZN(\V3/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M4/M1/_1_  (.A(\V3/V1/V2/v4 [3]),
    .B(ground),
    .Z(\V3/V1/V2/A3/M4/s1 ));
 AND2_X1 \V3/V1/V2/A3/M4/M2/_0_  (.A1(\V3/V1/V2/A3/M4/s1 ),
    .A2(\V3/V1/V2/A3/c3 ),
    .ZN(\V3/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M4/M2/_1_  (.A(\V3/V1/V2/A3/M4/s1 ),
    .B(\V3/V1/V2/A3/c3 ),
    .Z(\V3/V1/v2 [7]));
 OR2_X1 \V3/V1/V2/A3/M4/_0_  (.A1(\V3/V1/V2/A3/M4/c1 ),
    .A2(\V3/V1/V2/A3/M4/c2 ),
    .ZN(\V3/V1/V2/overflow ));
 AND2_X1 \V3/V1/V2/V1/HA1/_0_  (.A1(\V3/V1/V2/V1/w2 ),
    .A2(\V3/V1/V2/V1/w1 ),
    .ZN(\V3/V1/V2/V1/w4 ));
 XOR2_X2 \V3/V1/V2/V1/HA1/_1_  (.A(\V3/V1/V2/V1/w2 ),
    .B(\V3/V1/V2/V1/w1 ),
    .Z(\V3/V1/v2 [1]));
 AND2_X1 \V3/V1/V2/V1/HA2/_0_  (.A1(\V3/V1/V2/V1/w4 ),
    .A2(\V3/V1/V2/V1/w3 ),
    .ZN(\V3/V1/V2/v1 [3]));
 XOR2_X2 \V3/V1/V2/V1/HA2/_1_  (.A(\V3/V1/V2/V1/w4 ),
    .B(\V3/V1/V2/V1/w3 ),
    .Z(\V3/V1/V2/v1 [2]));
 AND2_X1 \V3/V1/V2/V1/_0_  (.A1(A[4]),
    .A2(B[16]),
    .ZN(\V3/V1/v2 [0]));
 AND2_X1 \V3/V1/V2/V1/_1_  (.A1(A[4]),
    .A2(B[17]),
    .ZN(\V3/V1/V2/V1/w1 ));
 AND2_X1 \V3/V1/V2/V1/_2_  (.A1(B[16]),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V1/w2 ));
 AND2_X1 \V3/V1/V2/V1/_3_  (.A1(B[17]),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V1/w3 ));
 AND2_X1 \V3/V1/V2/V2/HA1/_0_  (.A1(\V3/V1/V2/V2/w2 ),
    .A2(\V3/V1/V2/V2/w1 ),
    .ZN(\V3/V1/V2/V2/w4 ));
 XOR2_X2 \V3/V1/V2/V2/HA1/_1_  (.A(\V3/V1/V2/V2/w2 ),
    .B(\V3/V1/V2/V2/w1 ),
    .Z(\V3/V1/V2/v2 [1]));
 AND2_X1 \V3/V1/V2/V2/HA2/_0_  (.A1(\V3/V1/V2/V2/w4 ),
    .A2(\V3/V1/V2/V2/w3 ),
    .ZN(\V3/V1/V2/v2 [3]));
 XOR2_X2 \V3/V1/V2/V2/HA2/_1_  (.A(\V3/V1/V2/V2/w4 ),
    .B(\V3/V1/V2/V2/w3 ),
    .Z(\V3/V1/V2/v2 [2]));
 AND2_X1 \V3/V1/V2/V2/_0_  (.A1(A[6]),
    .A2(B[16]),
    .ZN(\V3/V1/V2/v2 [0]));
 AND2_X1 \V3/V1/V2/V2/_1_  (.A1(A[6]),
    .A2(B[17]),
    .ZN(\V3/V1/V2/V2/w1 ));
 AND2_X1 \V3/V1/V2/V2/_2_  (.A1(B[16]),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V2/w2 ));
 AND2_X1 \V3/V1/V2/V2/_3_  (.A1(B[17]),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V2/w3 ));
 AND2_X1 \V3/V1/V2/V3/HA1/_0_  (.A1(\V3/V1/V2/V3/w2 ),
    .A2(\V3/V1/V2/V3/w1 ),
    .ZN(\V3/V1/V2/V3/w4 ));
 XOR2_X2 \V3/V1/V2/V3/HA1/_1_  (.A(\V3/V1/V2/V3/w2 ),
    .B(\V3/V1/V2/V3/w1 ),
    .Z(\V3/V1/V2/v3 [1]));
 AND2_X1 \V3/V1/V2/V3/HA2/_0_  (.A1(\V3/V1/V2/V3/w4 ),
    .A2(\V3/V1/V2/V3/w3 ),
    .ZN(\V3/V1/V2/v3 [3]));
 XOR2_X2 \V3/V1/V2/V3/HA2/_1_  (.A(\V3/V1/V2/V3/w4 ),
    .B(\V3/V1/V2/V3/w3 ),
    .Z(\V3/V1/V2/v3 [2]));
 AND2_X1 \V3/V1/V2/V3/_0_  (.A1(A[4]),
    .A2(B[18]),
    .ZN(\V3/V1/V2/v3 [0]));
 AND2_X1 \V3/V1/V2/V3/_1_  (.A1(A[4]),
    .A2(B[19]),
    .ZN(\V3/V1/V2/V3/w1 ));
 AND2_X1 \V3/V1/V2/V3/_2_  (.A1(B[18]),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V3/w2 ));
 AND2_X1 \V3/V1/V2/V3/_3_  (.A1(B[19]),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V3/w3 ));
 AND2_X1 \V3/V1/V2/V4/HA1/_0_  (.A1(\V3/V1/V2/V4/w2 ),
    .A2(\V3/V1/V2/V4/w1 ),
    .ZN(\V3/V1/V2/V4/w4 ));
 XOR2_X2 \V3/V1/V2/V4/HA1/_1_  (.A(\V3/V1/V2/V4/w2 ),
    .B(\V3/V1/V2/V4/w1 ),
    .Z(\V3/V1/V2/v4 [1]));
 AND2_X1 \V3/V1/V2/V4/HA2/_0_  (.A1(\V3/V1/V2/V4/w4 ),
    .A2(\V3/V1/V2/V4/w3 ),
    .ZN(\V3/V1/V2/v4 [3]));
 XOR2_X2 \V3/V1/V2/V4/HA2/_1_  (.A(\V3/V1/V2/V4/w4 ),
    .B(\V3/V1/V2/V4/w3 ),
    .Z(\V3/V1/V2/v4 [2]));
 AND2_X1 \V3/V1/V2/V4/_0_  (.A1(A[6]),
    .A2(B[18]),
    .ZN(\V3/V1/V2/v4 [0]));
 AND2_X1 \V3/V1/V2/V4/_1_  (.A1(A[6]),
    .A2(B[19]),
    .ZN(\V3/V1/V2/V4/w1 ));
 AND2_X1 \V3/V1/V2/V4/_2_  (.A1(B[18]),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V4/w2 ));
 AND2_X1 \V3/V1/V2/V4/_3_  (.A1(B[19]),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V4/w3 ));
 OR2_X1 \V3/V1/V2/_0_  (.A1(\V3/V1/V2/c1 ),
    .A2(\V3/V1/V2/c2 ),
    .ZN(\V3/V1/V2/c3 ));
 AND2_X1 \V3/V1/V3/A1/M1/M1/_0_  (.A1(\V3/V1/V3/v2 [0]),
    .A2(\V3/V1/V3/v3 [0]),
    .ZN(\V3/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M1/M1/_1_  (.A(\V3/V1/V3/v2 [0]),
    .B(\V3/V1/V3/v3 [0]),
    .Z(\V3/V1/V3/A1/M1/s1 ));
 AND2_X1 \V3/V1/V3/A1/M1/M2/_0_  (.A1(\V3/V1/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M1/M2/_1_  (.A(\V3/V1/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/V3/s1 [0]));
 OR2_X1 \V3/V1/V3/A1/M1/_0_  (.A1(\V3/V1/V3/A1/M1/c1 ),
    .A2(\V3/V1/V3/A1/M1/c2 ),
    .ZN(\V3/V1/V3/A1/c1 ));
 AND2_X1 \V3/V1/V3/A1/M2/M1/_0_  (.A1(\V3/V1/V3/v2 [1]),
    .A2(\V3/V1/V3/v3 [1]),
    .ZN(\V3/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M2/M1/_1_  (.A(\V3/V1/V3/v2 [1]),
    .B(\V3/V1/V3/v3 [1]),
    .Z(\V3/V1/V3/A1/M2/s1 ));
 AND2_X1 \V3/V1/V3/A1/M2/M2/_0_  (.A1(\V3/V1/V3/A1/M2/s1 ),
    .A2(\V3/V1/V3/A1/c1 ),
    .ZN(\V3/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M2/M2/_1_  (.A(\V3/V1/V3/A1/M2/s1 ),
    .B(\V3/V1/V3/A1/c1 ),
    .Z(\V3/V1/V3/s1 [1]));
 OR2_X1 \V3/V1/V3/A1/M2/_0_  (.A1(\V3/V1/V3/A1/M2/c1 ),
    .A2(\V3/V1/V3/A1/M2/c2 ),
    .ZN(\V3/V1/V3/A1/c2 ));
 AND2_X1 \V3/V1/V3/A1/M3/M1/_0_  (.A1(\V3/V1/V3/v2 [2]),
    .A2(\V3/V1/V3/v3 [2]),
    .ZN(\V3/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M3/M1/_1_  (.A(\V3/V1/V3/v2 [2]),
    .B(\V3/V1/V3/v3 [2]),
    .Z(\V3/V1/V3/A1/M3/s1 ));
 AND2_X1 \V3/V1/V3/A1/M3/M2/_0_  (.A1(\V3/V1/V3/A1/M3/s1 ),
    .A2(\V3/V1/V3/A1/c2 ),
    .ZN(\V3/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M3/M2/_1_  (.A(\V3/V1/V3/A1/M3/s1 ),
    .B(\V3/V1/V3/A1/c2 ),
    .Z(\V3/V1/V3/s1 [2]));
 OR2_X1 \V3/V1/V3/A1/M3/_0_  (.A1(\V3/V1/V3/A1/M3/c1 ),
    .A2(\V3/V1/V3/A1/M3/c2 ),
    .ZN(\V3/V1/V3/A1/c3 ));
 AND2_X1 \V3/V1/V3/A1/M4/M1/_0_  (.A1(\V3/V1/V3/v2 [3]),
    .A2(\V3/V1/V3/v3 [3]),
    .ZN(\V3/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M4/M1/_1_  (.A(\V3/V1/V3/v2 [3]),
    .B(\V3/V1/V3/v3 [3]),
    .Z(\V3/V1/V3/A1/M4/s1 ));
 AND2_X1 \V3/V1/V3/A1/M4/M2/_0_  (.A1(\V3/V1/V3/A1/M4/s1 ),
    .A2(\V3/V1/V3/A1/c3 ),
    .ZN(\V3/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M4/M2/_1_  (.A(\V3/V1/V3/A1/M4/s1 ),
    .B(\V3/V1/V3/A1/c3 ),
    .Z(\V3/V1/V3/s1 [3]));
 OR2_X1 \V3/V1/V3/A1/M4/_0_  (.A1(\V3/V1/V3/A1/M4/c1 ),
    .A2(\V3/V1/V3/A1/M4/c2 ),
    .ZN(\V3/V1/V3/c1 ));
 AND2_X1 \V3/V1/V3/A2/M1/M1/_0_  (.A1(\V3/V1/V3/s1 [0]),
    .A2(\V3/V1/V3/v1 [2]),
    .ZN(\V3/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M1/M1/_1_  (.A(\V3/V1/V3/s1 [0]),
    .B(\V3/V1/V3/v1 [2]),
    .Z(\V3/V1/V3/A2/M1/s1 ));
 AND2_X1 \V3/V1/V3/A2/M1/M2/_0_  (.A1(\V3/V1/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M1/M2/_1_  (.A(\V3/V1/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v3 [2]));
 OR2_X1 \V3/V1/V3/A2/M1/_0_  (.A1(\V3/V1/V3/A2/M1/c1 ),
    .A2(\V3/V1/V3/A2/M1/c2 ),
    .ZN(\V3/V1/V3/A2/c1 ));
 AND2_X1 \V3/V1/V3/A2/M2/M1/_0_  (.A1(\V3/V1/V3/s1 [1]),
    .A2(\V3/V1/V3/v1 [3]),
    .ZN(\V3/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M2/M1/_1_  (.A(\V3/V1/V3/s1 [1]),
    .B(\V3/V1/V3/v1 [3]),
    .Z(\V3/V1/V3/A2/M2/s1 ));
 AND2_X1 \V3/V1/V3/A2/M2/M2/_0_  (.A1(\V3/V1/V3/A2/M2/s1 ),
    .A2(\V3/V1/V3/A2/c1 ),
    .ZN(\V3/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M2/M2/_1_  (.A(\V3/V1/V3/A2/M2/s1 ),
    .B(\V3/V1/V3/A2/c1 ),
    .Z(\V3/V1/v3 [3]));
 OR2_X1 \V3/V1/V3/A2/M2/_0_  (.A1(\V3/V1/V3/A2/M2/c1 ),
    .A2(\V3/V1/V3/A2/M2/c2 ),
    .ZN(\V3/V1/V3/A2/c2 ));
 AND2_X1 \V3/V1/V3/A2/M3/M1/_0_  (.A1(\V3/V1/V3/s1 [2]),
    .A2(ground),
    .ZN(\V3/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M3/M1/_1_  (.A(\V3/V1/V3/s1 [2]),
    .B(ground),
    .Z(\V3/V1/V3/A2/M3/s1 ));
 AND2_X1 \V3/V1/V3/A2/M3/M2/_0_  (.A1(\V3/V1/V3/A2/M3/s1 ),
    .A2(\V3/V1/V3/A2/c2 ),
    .ZN(\V3/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M3/M2/_1_  (.A(\V3/V1/V3/A2/M3/s1 ),
    .B(\V3/V1/V3/A2/c2 ),
    .Z(\V3/V1/V3/s2 [2]));
 OR2_X1 \V3/V1/V3/A2/M3/_0_  (.A1(\V3/V1/V3/A2/M3/c1 ),
    .A2(\V3/V1/V3/A2/M3/c2 ),
    .ZN(\V3/V1/V3/A2/c3 ));
 AND2_X1 \V3/V1/V3/A2/M4/M1/_0_  (.A1(\V3/V1/V3/s1 [3]),
    .A2(ground),
    .ZN(\V3/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M4/M1/_1_  (.A(\V3/V1/V3/s1 [3]),
    .B(ground),
    .Z(\V3/V1/V3/A2/M4/s1 ));
 AND2_X1 \V3/V1/V3/A2/M4/M2/_0_  (.A1(\V3/V1/V3/A2/M4/s1 ),
    .A2(\V3/V1/V3/A2/c3 ),
    .ZN(\V3/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M4/M2/_1_  (.A(\V3/V1/V3/A2/M4/s1 ),
    .B(\V3/V1/V3/A2/c3 ),
    .Z(\V3/V1/V3/s2 [3]));
 OR2_X1 \V3/V1/V3/A2/M4/_0_  (.A1(\V3/V1/V3/A2/M4/c1 ),
    .A2(\V3/V1/V3/A2/M4/c2 ),
    .ZN(\V3/V1/V3/c2 ));
 AND2_X1 \V3/V1/V3/A3/M1/M1/_0_  (.A1(\V3/V1/V3/v4 [0]),
    .A2(\V3/V1/V3/s2 [2]),
    .ZN(\V3/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M1/M1/_1_  (.A(\V3/V1/V3/v4 [0]),
    .B(\V3/V1/V3/s2 [2]),
    .Z(\V3/V1/V3/A3/M1/s1 ));
 AND2_X1 \V3/V1/V3/A3/M1/M2/_0_  (.A1(\V3/V1/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M1/M2/_1_  (.A(\V3/V1/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v3 [4]));
 OR2_X1 \V3/V1/V3/A3/M1/_0_  (.A1(\V3/V1/V3/A3/M1/c1 ),
    .A2(\V3/V1/V3/A3/M1/c2 ),
    .ZN(\V3/V1/V3/A3/c1 ));
 AND2_X1 \V3/V1/V3/A3/M2/M1/_0_  (.A1(\V3/V1/V3/v4 [1]),
    .A2(\V3/V1/V3/s2 [3]),
    .ZN(\V3/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M2/M1/_1_  (.A(\V3/V1/V3/v4 [1]),
    .B(\V3/V1/V3/s2 [3]),
    .Z(\V3/V1/V3/A3/M2/s1 ));
 AND2_X1 \V3/V1/V3/A3/M2/M2/_0_  (.A1(\V3/V1/V3/A3/M2/s1 ),
    .A2(\V3/V1/V3/A3/c1 ),
    .ZN(\V3/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M2/M2/_1_  (.A(\V3/V1/V3/A3/M2/s1 ),
    .B(\V3/V1/V3/A3/c1 ),
    .Z(\V3/V1/v3 [5]));
 OR2_X1 \V3/V1/V3/A3/M2/_0_  (.A1(\V3/V1/V3/A3/M2/c1 ),
    .A2(\V3/V1/V3/A3/M2/c2 ),
    .ZN(\V3/V1/V3/A3/c2 ));
 AND2_X1 \V3/V1/V3/A3/M3/M1/_0_  (.A1(\V3/V1/V3/v4 [2]),
    .A2(\V3/V1/V3/c3 ),
    .ZN(\V3/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M3/M1/_1_  (.A(\V3/V1/V3/v4 [2]),
    .B(\V3/V1/V3/c3 ),
    .Z(\V3/V1/V3/A3/M3/s1 ));
 AND2_X1 \V3/V1/V3/A3/M3/M2/_0_  (.A1(\V3/V1/V3/A3/M3/s1 ),
    .A2(\V3/V1/V3/A3/c2 ),
    .ZN(\V3/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M3/M2/_1_  (.A(\V3/V1/V3/A3/M3/s1 ),
    .B(\V3/V1/V3/A3/c2 ),
    .Z(\V3/V1/v3 [6]));
 OR2_X1 \V3/V1/V3/A3/M3/_0_  (.A1(\V3/V1/V3/A3/M3/c1 ),
    .A2(\V3/V1/V3/A3/M3/c2 ),
    .ZN(\V3/V1/V3/A3/c3 ));
 AND2_X1 \V3/V1/V3/A3/M4/M1/_0_  (.A1(\V3/V1/V3/v4 [3]),
    .A2(ground),
    .ZN(\V3/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M4/M1/_1_  (.A(\V3/V1/V3/v4 [3]),
    .B(ground),
    .Z(\V3/V1/V3/A3/M4/s1 ));
 AND2_X1 \V3/V1/V3/A3/M4/M2/_0_  (.A1(\V3/V1/V3/A3/M4/s1 ),
    .A2(\V3/V1/V3/A3/c3 ),
    .ZN(\V3/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M4/M2/_1_  (.A(\V3/V1/V3/A3/M4/s1 ),
    .B(\V3/V1/V3/A3/c3 ),
    .Z(\V3/V1/v3 [7]));
 OR2_X1 \V3/V1/V3/A3/M4/_0_  (.A1(\V3/V1/V3/A3/M4/c1 ),
    .A2(\V3/V1/V3/A3/M4/c2 ),
    .ZN(\V3/V1/V3/overflow ));
 AND2_X1 \V3/V1/V3/V1/HA1/_0_  (.A1(\V3/V1/V3/V1/w2 ),
    .A2(\V3/V1/V3/V1/w1 ),
    .ZN(\V3/V1/V3/V1/w4 ));
 XOR2_X2 \V3/V1/V3/V1/HA1/_1_  (.A(\V3/V1/V3/V1/w2 ),
    .B(\V3/V1/V3/V1/w1 ),
    .Z(\V3/V1/v3 [1]));
 AND2_X1 \V3/V1/V3/V1/HA2/_0_  (.A1(\V3/V1/V3/V1/w4 ),
    .A2(\V3/V1/V3/V1/w3 ),
    .ZN(\V3/V1/V3/v1 [3]));
 XOR2_X2 \V3/V1/V3/V1/HA2/_1_  (.A(\V3/V1/V3/V1/w4 ),
    .B(\V3/V1/V3/V1/w3 ),
    .Z(\V3/V1/V3/v1 [2]));
 AND2_X1 \V3/V1/V3/V1/_0_  (.A1(A[0]),
    .A2(B[20]),
    .ZN(\V3/V1/v3 [0]));
 AND2_X1 \V3/V1/V3/V1/_1_  (.A1(A[0]),
    .A2(B[21]),
    .ZN(\V3/V1/V3/V1/w1 ));
 AND2_X1 \V3/V1/V3/V1/_2_  (.A1(B[20]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V1/w2 ));
 AND2_X1 \V3/V1/V3/V1/_3_  (.A1(B[21]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V1/w3 ));
 AND2_X1 \V3/V1/V3/V2/HA1/_0_  (.A1(\V3/V1/V3/V2/w2 ),
    .A2(\V3/V1/V3/V2/w1 ),
    .ZN(\V3/V1/V3/V2/w4 ));
 XOR2_X2 \V3/V1/V3/V2/HA1/_1_  (.A(\V3/V1/V3/V2/w2 ),
    .B(\V3/V1/V3/V2/w1 ),
    .Z(\V3/V1/V3/v2 [1]));
 AND2_X1 \V3/V1/V3/V2/HA2/_0_  (.A1(\V3/V1/V3/V2/w4 ),
    .A2(\V3/V1/V3/V2/w3 ),
    .ZN(\V3/V1/V3/v2 [3]));
 XOR2_X2 \V3/V1/V3/V2/HA2/_1_  (.A(\V3/V1/V3/V2/w4 ),
    .B(\V3/V1/V3/V2/w3 ),
    .Z(\V3/V1/V3/v2 [2]));
 AND2_X1 \V3/V1/V3/V2/_0_  (.A1(A[2]),
    .A2(B[20]),
    .ZN(\V3/V1/V3/v2 [0]));
 AND2_X1 \V3/V1/V3/V2/_1_  (.A1(A[2]),
    .A2(B[21]),
    .ZN(\V3/V1/V3/V2/w1 ));
 AND2_X1 \V3/V1/V3/V2/_2_  (.A1(B[20]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V2/w2 ));
 AND2_X1 \V3/V1/V3/V2/_3_  (.A1(B[21]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V2/w3 ));
 AND2_X1 \V3/V1/V3/V3/HA1/_0_  (.A1(\V3/V1/V3/V3/w2 ),
    .A2(\V3/V1/V3/V3/w1 ),
    .ZN(\V3/V1/V3/V3/w4 ));
 XOR2_X2 \V3/V1/V3/V3/HA1/_1_  (.A(\V3/V1/V3/V3/w2 ),
    .B(\V3/V1/V3/V3/w1 ),
    .Z(\V3/V1/V3/v3 [1]));
 AND2_X1 \V3/V1/V3/V3/HA2/_0_  (.A1(\V3/V1/V3/V3/w4 ),
    .A2(\V3/V1/V3/V3/w3 ),
    .ZN(\V3/V1/V3/v3 [3]));
 XOR2_X2 \V3/V1/V3/V3/HA2/_1_  (.A(\V3/V1/V3/V3/w4 ),
    .B(\V3/V1/V3/V3/w3 ),
    .Z(\V3/V1/V3/v3 [2]));
 AND2_X1 \V3/V1/V3/V3/_0_  (.A1(A[0]),
    .A2(B[22]),
    .ZN(\V3/V1/V3/v3 [0]));
 AND2_X1 \V3/V1/V3/V3/_1_  (.A1(A[0]),
    .A2(B[23]),
    .ZN(\V3/V1/V3/V3/w1 ));
 AND2_X1 \V3/V1/V3/V3/_2_  (.A1(B[22]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V3/w2 ));
 AND2_X1 \V3/V1/V3/V3/_3_  (.A1(B[23]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V3/w3 ));
 AND2_X1 \V3/V1/V3/V4/HA1/_0_  (.A1(\V3/V1/V3/V4/w2 ),
    .A2(\V3/V1/V3/V4/w1 ),
    .ZN(\V3/V1/V3/V4/w4 ));
 XOR2_X2 \V3/V1/V3/V4/HA1/_1_  (.A(\V3/V1/V3/V4/w2 ),
    .B(\V3/V1/V3/V4/w1 ),
    .Z(\V3/V1/V3/v4 [1]));
 AND2_X1 \V3/V1/V3/V4/HA2/_0_  (.A1(\V3/V1/V3/V4/w4 ),
    .A2(\V3/V1/V3/V4/w3 ),
    .ZN(\V3/V1/V3/v4 [3]));
 XOR2_X2 \V3/V1/V3/V4/HA2/_1_  (.A(\V3/V1/V3/V4/w4 ),
    .B(\V3/V1/V3/V4/w3 ),
    .Z(\V3/V1/V3/v4 [2]));
 AND2_X1 \V3/V1/V3/V4/_0_  (.A1(A[2]),
    .A2(B[22]),
    .ZN(\V3/V1/V3/v4 [0]));
 AND2_X1 \V3/V1/V3/V4/_1_  (.A1(A[2]),
    .A2(B[23]),
    .ZN(\V3/V1/V3/V4/w1 ));
 AND2_X1 \V3/V1/V3/V4/_2_  (.A1(B[22]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V4/w2 ));
 AND2_X1 \V3/V1/V3/V4/_3_  (.A1(B[23]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V4/w3 ));
 OR2_X1 \V3/V1/V3/_0_  (.A1(\V3/V1/V3/c1 ),
    .A2(\V3/V1/V3/c2 ),
    .ZN(\V3/V1/V3/c3 ));
 AND2_X1 \V3/V1/V4/A1/M1/M1/_0_  (.A1(\V3/V1/V4/v2 [0]),
    .A2(\V3/V1/V4/v3 [0]),
    .ZN(\V3/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M1/M1/_1_  (.A(\V3/V1/V4/v2 [0]),
    .B(\V3/V1/V4/v3 [0]),
    .Z(\V3/V1/V4/A1/M1/s1 ));
 AND2_X1 \V3/V1/V4/A1/M1/M2/_0_  (.A1(\V3/V1/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M1/M2/_1_  (.A(\V3/V1/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/V4/s1 [0]));
 OR2_X1 \V3/V1/V4/A1/M1/_0_  (.A1(\V3/V1/V4/A1/M1/c1 ),
    .A2(\V3/V1/V4/A1/M1/c2 ),
    .ZN(\V3/V1/V4/A1/c1 ));
 AND2_X1 \V3/V1/V4/A1/M2/M1/_0_  (.A1(\V3/V1/V4/v2 [1]),
    .A2(\V3/V1/V4/v3 [1]),
    .ZN(\V3/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M2/M1/_1_  (.A(\V3/V1/V4/v2 [1]),
    .B(\V3/V1/V4/v3 [1]),
    .Z(\V3/V1/V4/A1/M2/s1 ));
 AND2_X1 \V3/V1/V4/A1/M2/M2/_0_  (.A1(\V3/V1/V4/A1/M2/s1 ),
    .A2(\V3/V1/V4/A1/c1 ),
    .ZN(\V3/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M2/M2/_1_  (.A(\V3/V1/V4/A1/M2/s1 ),
    .B(\V3/V1/V4/A1/c1 ),
    .Z(\V3/V1/V4/s1 [1]));
 OR2_X1 \V3/V1/V4/A1/M2/_0_  (.A1(\V3/V1/V4/A1/M2/c1 ),
    .A2(\V3/V1/V4/A1/M2/c2 ),
    .ZN(\V3/V1/V4/A1/c2 ));
 AND2_X1 \V3/V1/V4/A1/M3/M1/_0_  (.A1(\V3/V1/V4/v2 [2]),
    .A2(\V3/V1/V4/v3 [2]),
    .ZN(\V3/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M3/M1/_1_  (.A(\V3/V1/V4/v2 [2]),
    .B(\V3/V1/V4/v3 [2]),
    .Z(\V3/V1/V4/A1/M3/s1 ));
 AND2_X1 \V3/V1/V4/A1/M3/M2/_0_  (.A1(\V3/V1/V4/A1/M3/s1 ),
    .A2(\V3/V1/V4/A1/c2 ),
    .ZN(\V3/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M3/M2/_1_  (.A(\V3/V1/V4/A1/M3/s1 ),
    .B(\V3/V1/V4/A1/c2 ),
    .Z(\V3/V1/V4/s1 [2]));
 OR2_X1 \V3/V1/V4/A1/M3/_0_  (.A1(\V3/V1/V4/A1/M3/c1 ),
    .A2(\V3/V1/V4/A1/M3/c2 ),
    .ZN(\V3/V1/V4/A1/c3 ));
 AND2_X1 \V3/V1/V4/A1/M4/M1/_0_  (.A1(\V3/V1/V4/v2 [3]),
    .A2(\V3/V1/V4/v3 [3]),
    .ZN(\V3/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M4/M1/_1_  (.A(\V3/V1/V4/v2 [3]),
    .B(\V3/V1/V4/v3 [3]),
    .Z(\V3/V1/V4/A1/M4/s1 ));
 AND2_X1 \V3/V1/V4/A1/M4/M2/_0_  (.A1(\V3/V1/V4/A1/M4/s1 ),
    .A2(\V3/V1/V4/A1/c3 ),
    .ZN(\V3/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M4/M2/_1_  (.A(\V3/V1/V4/A1/M4/s1 ),
    .B(\V3/V1/V4/A1/c3 ),
    .Z(\V3/V1/V4/s1 [3]));
 OR2_X1 \V3/V1/V4/A1/M4/_0_  (.A1(\V3/V1/V4/A1/M4/c1 ),
    .A2(\V3/V1/V4/A1/M4/c2 ),
    .ZN(\V3/V1/V4/c1 ));
 AND2_X1 \V3/V1/V4/A2/M1/M1/_0_  (.A1(\V3/V1/V4/s1 [0]),
    .A2(\V3/V1/V4/v1 [2]),
    .ZN(\V3/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M1/M1/_1_  (.A(\V3/V1/V4/s1 [0]),
    .B(\V3/V1/V4/v1 [2]),
    .Z(\V3/V1/V4/A2/M1/s1 ));
 AND2_X1 \V3/V1/V4/A2/M1/M2/_0_  (.A1(\V3/V1/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M1/M2/_1_  (.A(\V3/V1/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v4 [2]));
 OR2_X1 \V3/V1/V4/A2/M1/_0_  (.A1(\V3/V1/V4/A2/M1/c1 ),
    .A2(\V3/V1/V4/A2/M1/c2 ),
    .ZN(\V3/V1/V4/A2/c1 ));
 AND2_X1 \V3/V1/V4/A2/M2/M1/_0_  (.A1(\V3/V1/V4/s1 [1]),
    .A2(\V3/V1/V4/v1 [3]),
    .ZN(\V3/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M2/M1/_1_  (.A(\V3/V1/V4/s1 [1]),
    .B(\V3/V1/V4/v1 [3]),
    .Z(\V3/V1/V4/A2/M2/s1 ));
 AND2_X1 \V3/V1/V4/A2/M2/M2/_0_  (.A1(\V3/V1/V4/A2/M2/s1 ),
    .A2(\V3/V1/V4/A2/c1 ),
    .ZN(\V3/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M2/M2/_1_  (.A(\V3/V1/V4/A2/M2/s1 ),
    .B(\V3/V1/V4/A2/c1 ),
    .Z(\V3/V1/v4 [3]));
 OR2_X1 \V3/V1/V4/A2/M2/_0_  (.A1(\V3/V1/V4/A2/M2/c1 ),
    .A2(\V3/V1/V4/A2/M2/c2 ),
    .ZN(\V3/V1/V4/A2/c2 ));
 AND2_X1 \V3/V1/V4/A2/M3/M1/_0_  (.A1(\V3/V1/V4/s1 [2]),
    .A2(ground),
    .ZN(\V3/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M3/M1/_1_  (.A(\V3/V1/V4/s1 [2]),
    .B(ground),
    .Z(\V3/V1/V4/A2/M3/s1 ));
 AND2_X1 \V3/V1/V4/A2/M3/M2/_0_  (.A1(\V3/V1/V4/A2/M3/s1 ),
    .A2(\V3/V1/V4/A2/c2 ),
    .ZN(\V3/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M3/M2/_1_  (.A(\V3/V1/V4/A2/M3/s1 ),
    .B(\V3/V1/V4/A2/c2 ),
    .Z(\V3/V1/V4/s2 [2]));
 OR2_X1 \V3/V1/V4/A2/M3/_0_  (.A1(\V3/V1/V4/A2/M3/c1 ),
    .A2(\V3/V1/V4/A2/M3/c2 ),
    .ZN(\V3/V1/V4/A2/c3 ));
 AND2_X1 \V3/V1/V4/A2/M4/M1/_0_  (.A1(\V3/V1/V4/s1 [3]),
    .A2(ground),
    .ZN(\V3/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M4/M1/_1_  (.A(\V3/V1/V4/s1 [3]),
    .B(ground),
    .Z(\V3/V1/V4/A2/M4/s1 ));
 AND2_X1 \V3/V1/V4/A2/M4/M2/_0_  (.A1(\V3/V1/V4/A2/M4/s1 ),
    .A2(\V3/V1/V4/A2/c3 ),
    .ZN(\V3/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M4/M2/_1_  (.A(\V3/V1/V4/A2/M4/s1 ),
    .B(\V3/V1/V4/A2/c3 ),
    .Z(\V3/V1/V4/s2 [3]));
 OR2_X1 \V3/V1/V4/A2/M4/_0_  (.A1(\V3/V1/V4/A2/M4/c1 ),
    .A2(\V3/V1/V4/A2/M4/c2 ),
    .ZN(\V3/V1/V4/c2 ));
 AND2_X1 \V3/V1/V4/A3/M1/M1/_0_  (.A1(\V3/V1/V4/v4 [0]),
    .A2(\V3/V1/V4/s2 [2]),
    .ZN(\V3/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M1/M1/_1_  (.A(\V3/V1/V4/v4 [0]),
    .B(\V3/V1/V4/s2 [2]),
    .Z(\V3/V1/V4/A3/M1/s1 ));
 AND2_X1 \V3/V1/V4/A3/M1/M2/_0_  (.A1(\V3/V1/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M1/M2/_1_  (.A(\V3/V1/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V1/v4 [4]));
 OR2_X1 \V3/V1/V4/A3/M1/_0_  (.A1(\V3/V1/V4/A3/M1/c1 ),
    .A2(\V3/V1/V4/A3/M1/c2 ),
    .ZN(\V3/V1/V4/A3/c1 ));
 AND2_X1 \V3/V1/V4/A3/M2/M1/_0_  (.A1(\V3/V1/V4/v4 [1]),
    .A2(\V3/V1/V4/s2 [3]),
    .ZN(\V3/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M2/M1/_1_  (.A(\V3/V1/V4/v4 [1]),
    .B(\V3/V1/V4/s2 [3]),
    .Z(\V3/V1/V4/A3/M2/s1 ));
 AND2_X1 \V3/V1/V4/A3/M2/M2/_0_  (.A1(\V3/V1/V4/A3/M2/s1 ),
    .A2(\V3/V1/V4/A3/c1 ),
    .ZN(\V3/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M2/M2/_1_  (.A(\V3/V1/V4/A3/M2/s1 ),
    .B(\V3/V1/V4/A3/c1 ),
    .Z(\V3/V1/v4 [5]));
 OR2_X1 \V3/V1/V4/A3/M2/_0_  (.A1(\V3/V1/V4/A3/M2/c1 ),
    .A2(\V3/V1/V4/A3/M2/c2 ),
    .ZN(\V3/V1/V4/A3/c2 ));
 AND2_X1 \V3/V1/V4/A3/M3/M1/_0_  (.A1(\V3/V1/V4/v4 [2]),
    .A2(\V3/V1/V4/c3 ),
    .ZN(\V3/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M3/M1/_1_  (.A(\V3/V1/V4/v4 [2]),
    .B(\V3/V1/V4/c3 ),
    .Z(\V3/V1/V4/A3/M3/s1 ));
 AND2_X1 \V3/V1/V4/A3/M3/M2/_0_  (.A1(\V3/V1/V4/A3/M3/s1 ),
    .A2(\V3/V1/V4/A3/c2 ),
    .ZN(\V3/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M3/M2/_1_  (.A(\V3/V1/V4/A3/M3/s1 ),
    .B(\V3/V1/V4/A3/c2 ),
    .Z(\V3/V1/v4 [6]));
 OR2_X1 \V3/V1/V4/A3/M3/_0_  (.A1(\V3/V1/V4/A3/M3/c1 ),
    .A2(\V3/V1/V4/A3/M3/c2 ),
    .ZN(\V3/V1/V4/A3/c3 ));
 AND2_X1 \V3/V1/V4/A3/M4/M1/_0_  (.A1(\V3/V1/V4/v4 [3]),
    .A2(ground),
    .ZN(\V3/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M4/M1/_1_  (.A(\V3/V1/V4/v4 [3]),
    .B(ground),
    .Z(\V3/V1/V4/A3/M4/s1 ));
 AND2_X1 \V3/V1/V4/A3/M4/M2/_0_  (.A1(\V3/V1/V4/A3/M4/s1 ),
    .A2(\V3/V1/V4/A3/c3 ),
    .ZN(\V3/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M4/M2/_1_  (.A(\V3/V1/V4/A3/M4/s1 ),
    .B(\V3/V1/V4/A3/c3 ),
    .Z(\V3/V1/v4 [7]));
 OR2_X1 \V3/V1/V4/A3/M4/_0_  (.A1(\V3/V1/V4/A3/M4/c1 ),
    .A2(\V3/V1/V4/A3/M4/c2 ),
    .ZN(\V3/V1/V4/overflow ));
 AND2_X1 \V3/V1/V4/V1/HA1/_0_  (.A1(\V3/V1/V4/V1/w2 ),
    .A2(\V3/V1/V4/V1/w1 ),
    .ZN(\V3/V1/V4/V1/w4 ));
 XOR2_X2 \V3/V1/V4/V1/HA1/_1_  (.A(\V3/V1/V4/V1/w2 ),
    .B(\V3/V1/V4/V1/w1 ),
    .Z(\V3/V1/v4 [1]));
 AND2_X1 \V3/V1/V4/V1/HA2/_0_  (.A1(\V3/V1/V4/V1/w4 ),
    .A2(\V3/V1/V4/V1/w3 ),
    .ZN(\V3/V1/V4/v1 [3]));
 XOR2_X2 \V3/V1/V4/V1/HA2/_1_  (.A(\V3/V1/V4/V1/w4 ),
    .B(\V3/V1/V4/V1/w3 ),
    .Z(\V3/V1/V4/v1 [2]));
 AND2_X1 \V3/V1/V4/V1/_0_  (.A1(A[4]),
    .A2(B[20]),
    .ZN(\V3/V1/v4 [0]));
 AND2_X1 \V3/V1/V4/V1/_1_  (.A1(A[4]),
    .A2(B[21]),
    .ZN(\V3/V1/V4/V1/w1 ));
 AND2_X1 \V3/V1/V4/V1/_2_  (.A1(B[20]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V1/w2 ));
 AND2_X1 \V3/V1/V4/V1/_3_  (.A1(B[21]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V1/w3 ));
 AND2_X1 \V3/V1/V4/V2/HA1/_0_  (.A1(\V3/V1/V4/V2/w2 ),
    .A2(\V3/V1/V4/V2/w1 ),
    .ZN(\V3/V1/V4/V2/w4 ));
 XOR2_X2 \V3/V1/V4/V2/HA1/_1_  (.A(\V3/V1/V4/V2/w2 ),
    .B(\V3/V1/V4/V2/w1 ),
    .Z(\V3/V1/V4/v2 [1]));
 AND2_X1 \V3/V1/V4/V2/HA2/_0_  (.A1(\V3/V1/V4/V2/w4 ),
    .A2(\V3/V1/V4/V2/w3 ),
    .ZN(\V3/V1/V4/v2 [3]));
 XOR2_X2 \V3/V1/V4/V2/HA2/_1_  (.A(\V3/V1/V4/V2/w4 ),
    .B(\V3/V1/V4/V2/w3 ),
    .Z(\V3/V1/V4/v2 [2]));
 AND2_X1 \V3/V1/V4/V2/_0_  (.A1(A[6]),
    .A2(B[20]),
    .ZN(\V3/V1/V4/v2 [0]));
 AND2_X1 \V3/V1/V4/V2/_1_  (.A1(A[6]),
    .A2(B[21]),
    .ZN(\V3/V1/V4/V2/w1 ));
 AND2_X1 \V3/V1/V4/V2/_2_  (.A1(B[20]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V2/w2 ));
 AND2_X1 \V3/V1/V4/V2/_3_  (.A1(B[21]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V2/w3 ));
 AND2_X1 \V3/V1/V4/V3/HA1/_0_  (.A1(\V3/V1/V4/V3/w2 ),
    .A2(\V3/V1/V4/V3/w1 ),
    .ZN(\V3/V1/V4/V3/w4 ));
 XOR2_X2 \V3/V1/V4/V3/HA1/_1_  (.A(\V3/V1/V4/V3/w2 ),
    .B(\V3/V1/V4/V3/w1 ),
    .Z(\V3/V1/V4/v3 [1]));
 AND2_X1 \V3/V1/V4/V3/HA2/_0_  (.A1(\V3/V1/V4/V3/w4 ),
    .A2(\V3/V1/V4/V3/w3 ),
    .ZN(\V3/V1/V4/v3 [3]));
 XOR2_X2 \V3/V1/V4/V3/HA2/_1_  (.A(\V3/V1/V4/V3/w4 ),
    .B(\V3/V1/V4/V3/w3 ),
    .Z(\V3/V1/V4/v3 [2]));
 AND2_X1 \V3/V1/V4/V3/_0_  (.A1(A[4]),
    .A2(B[22]),
    .ZN(\V3/V1/V4/v3 [0]));
 AND2_X1 \V3/V1/V4/V3/_1_  (.A1(A[4]),
    .A2(B[23]),
    .ZN(\V3/V1/V4/V3/w1 ));
 AND2_X1 \V3/V1/V4/V3/_2_  (.A1(B[22]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V3/w2 ));
 AND2_X1 \V3/V1/V4/V3/_3_  (.A1(B[23]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V3/w3 ));
 AND2_X1 \V3/V1/V4/V4/HA1/_0_  (.A1(\V3/V1/V4/V4/w2 ),
    .A2(\V3/V1/V4/V4/w1 ),
    .ZN(\V3/V1/V4/V4/w4 ));
 XOR2_X2 \V3/V1/V4/V4/HA1/_1_  (.A(\V3/V1/V4/V4/w2 ),
    .B(\V3/V1/V4/V4/w1 ),
    .Z(\V3/V1/V4/v4 [1]));
 AND2_X1 \V3/V1/V4/V4/HA2/_0_  (.A1(\V3/V1/V4/V4/w4 ),
    .A2(\V3/V1/V4/V4/w3 ),
    .ZN(\V3/V1/V4/v4 [3]));
 XOR2_X2 \V3/V1/V4/V4/HA2/_1_  (.A(\V3/V1/V4/V4/w4 ),
    .B(\V3/V1/V4/V4/w3 ),
    .Z(\V3/V1/V4/v4 [2]));
 AND2_X1 \V3/V1/V4/V4/_0_  (.A1(A[6]),
    .A2(B[22]),
    .ZN(\V3/V1/V4/v4 [0]));
 AND2_X1 \V3/V1/V4/V4/_1_  (.A1(A[6]),
    .A2(B[23]),
    .ZN(\V3/V1/V4/V4/w1 ));
 AND2_X1 \V3/V1/V4/V4/_2_  (.A1(B[22]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V4/w2 ));
 AND2_X1 \V3/V1/V4/V4/_3_  (.A1(B[23]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V4/w3 ));
 OR2_X1 \V3/V1/V4/_0_  (.A1(\V3/V1/V4/c1 ),
    .A2(\V3/V1/V4/c2 ),
    .ZN(\V3/V1/V4/c3 ));
 OR2_X1 \V3/V1/_0_  (.A1(\V3/V1/c1 ),
    .A2(\V3/V1/c2 ),
    .ZN(\V3/V1/c3 ));
 AND2_X1 \V3/V2/A1/A1/M1/M1/_0_  (.A1(\V3/V2/v2 [0]),
    .A2(\V3/V2/v3 [0]),
    .ZN(\V3/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M1/M1/_1_  (.A(\V3/V2/v2 [0]),
    .B(\V3/V2/v3 [0]),
    .Z(\V3/V2/A1/A1/M1/s1 ));
 AND2_X1 \V3/V2/A1/A1/M1/M2/_0_  (.A1(\V3/V2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M1/M2/_1_  (.A(\V3/V2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/s1 [0]));
 OR2_X1 \V3/V2/A1/A1/M1/_0_  (.A1(\V3/V2/A1/A1/M1/c1 ),
    .A2(\V3/V2/A1/A1/M1/c2 ),
    .ZN(\V3/V2/A1/A1/c1 ));
 AND2_X1 \V3/V2/A1/A1/M2/M1/_0_  (.A1(\V3/V2/v2 [1]),
    .A2(\V3/V2/v3 [1]),
    .ZN(\V3/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M2/M1/_1_  (.A(\V3/V2/v2 [1]),
    .B(\V3/V2/v3 [1]),
    .Z(\V3/V2/A1/A1/M2/s1 ));
 AND2_X1 \V3/V2/A1/A1/M2/M2/_0_  (.A1(\V3/V2/A1/A1/M2/s1 ),
    .A2(\V3/V2/A1/A1/c1 ),
    .ZN(\V3/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M2/M2/_1_  (.A(\V3/V2/A1/A1/M2/s1 ),
    .B(\V3/V2/A1/A1/c1 ),
    .Z(\V3/V2/s1 [1]));
 OR2_X1 \V3/V2/A1/A1/M2/_0_  (.A1(\V3/V2/A1/A1/M2/c1 ),
    .A2(\V3/V2/A1/A1/M2/c2 ),
    .ZN(\V3/V2/A1/A1/c2 ));
 AND2_X1 \V3/V2/A1/A1/M3/M1/_0_  (.A1(\V3/V2/v2 [2]),
    .A2(\V3/V2/v3 [2]),
    .ZN(\V3/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M3/M1/_1_  (.A(\V3/V2/v2 [2]),
    .B(\V3/V2/v3 [2]),
    .Z(\V3/V2/A1/A1/M3/s1 ));
 AND2_X1 \V3/V2/A1/A1/M3/M2/_0_  (.A1(\V3/V2/A1/A1/M3/s1 ),
    .A2(\V3/V2/A1/A1/c2 ),
    .ZN(\V3/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M3/M2/_1_  (.A(\V3/V2/A1/A1/M3/s1 ),
    .B(\V3/V2/A1/A1/c2 ),
    .Z(\V3/V2/s1 [2]));
 OR2_X1 \V3/V2/A1/A1/M3/_0_  (.A1(\V3/V2/A1/A1/M3/c1 ),
    .A2(\V3/V2/A1/A1/M3/c2 ),
    .ZN(\V3/V2/A1/A1/c3 ));
 AND2_X1 \V3/V2/A1/A1/M4/M1/_0_  (.A1(\V3/V2/v2 [3]),
    .A2(\V3/V2/v3 [3]),
    .ZN(\V3/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M4/M1/_1_  (.A(\V3/V2/v2 [3]),
    .B(\V3/V2/v3 [3]),
    .Z(\V3/V2/A1/A1/M4/s1 ));
 AND2_X1 \V3/V2/A1/A1/M4/M2/_0_  (.A1(\V3/V2/A1/A1/M4/s1 ),
    .A2(\V3/V2/A1/A1/c3 ),
    .ZN(\V3/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M4/M2/_1_  (.A(\V3/V2/A1/A1/M4/s1 ),
    .B(\V3/V2/A1/A1/c3 ),
    .Z(\V3/V2/s1 [3]));
 OR2_X1 \V3/V2/A1/A1/M4/_0_  (.A1(\V3/V2/A1/A1/M4/c1 ),
    .A2(\V3/V2/A1/A1/M4/c2 ),
    .ZN(\V3/V2/A1/c1 ));
 AND2_X1 \V3/V2/A1/A2/M1/M1/_0_  (.A1(\V3/V2/v2 [4]),
    .A2(\V3/V2/v3 [4]),
    .ZN(\V3/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M1/M1/_1_  (.A(\V3/V2/v2 [4]),
    .B(\V3/V2/v3 [4]),
    .Z(\V3/V2/A1/A2/M1/s1 ));
 AND2_X1 \V3/V2/A1/A2/M1/M2/_0_  (.A1(\V3/V2/A1/A2/M1/s1 ),
    .A2(\V3/V2/A1/c1 ),
    .ZN(\V3/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M1/M2/_1_  (.A(\V3/V2/A1/A2/M1/s1 ),
    .B(\V3/V2/A1/c1 ),
    .Z(\V3/V2/s1 [4]));
 OR2_X1 \V3/V2/A1/A2/M1/_0_  (.A1(\V3/V2/A1/A2/M1/c1 ),
    .A2(\V3/V2/A1/A2/M1/c2 ),
    .ZN(\V3/V2/A1/A2/c1 ));
 AND2_X1 \V3/V2/A1/A2/M2/M1/_0_  (.A1(\V3/V2/v2 [5]),
    .A2(\V3/V2/v3 [5]),
    .ZN(\V3/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M2/M1/_1_  (.A(\V3/V2/v2 [5]),
    .B(\V3/V2/v3 [5]),
    .Z(\V3/V2/A1/A2/M2/s1 ));
 AND2_X1 \V3/V2/A1/A2/M2/M2/_0_  (.A1(\V3/V2/A1/A2/M2/s1 ),
    .A2(\V3/V2/A1/A2/c1 ),
    .ZN(\V3/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M2/M2/_1_  (.A(\V3/V2/A1/A2/M2/s1 ),
    .B(\V3/V2/A1/A2/c1 ),
    .Z(\V3/V2/s1 [5]));
 OR2_X1 \V3/V2/A1/A2/M2/_0_  (.A1(\V3/V2/A1/A2/M2/c1 ),
    .A2(\V3/V2/A1/A2/M2/c2 ),
    .ZN(\V3/V2/A1/A2/c2 ));
 AND2_X1 \V3/V2/A1/A2/M3/M1/_0_  (.A1(\V3/V2/v2 [6]),
    .A2(\V3/V2/v3 [6]),
    .ZN(\V3/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M3/M1/_1_  (.A(\V3/V2/v2 [6]),
    .B(\V3/V2/v3 [6]),
    .Z(\V3/V2/A1/A2/M3/s1 ));
 AND2_X1 \V3/V2/A1/A2/M3/M2/_0_  (.A1(\V3/V2/A1/A2/M3/s1 ),
    .A2(\V3/V2/A1/A2/c2 ),
    .ZN(\V3/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M3/M2/_1_  (.A(\V3/V2/A1/A2/M3/s1 ),
    .B(\V3/V2/A1/A2/c2 ),
    .Z(\V3/V2/s1 [6]));
 OR2_X1 \V3/V2/A1/A2/M3/_0_  (.A1(\V3/V2/A1/A2/M3/c1 ),
    .A2(\V3/V2/A1/A2/M3/c2 ),
    .ZN(\V3/V2/A1/A2/c3 ));
 AND2_X1 \V3/V2/A1/A2/M4/M1/_0_  (.A1(\V3/V2/v2 [7]),
    .A2(\V3/V2/v3 [7]),
    .ZN(\V3/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M4/M1/_1_  (.A(\V3/V2/v2 [7]),
    .B(\V3/V2/v3 [7]),
    .Z(\V3/V2/A1/A2/M4/s1 ));
 AND2_X1 \V3/V2/A1/A2/M4/M2/_0_  (.A1(\V3/V2/A1/A2/M4/s1 ),
    .A2(\V3/V2/A1/A2/c3 ),
    .ZN(\V3/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M4/M2/_1_  (.A(\V3/V2/A1/A2/M4/s1 ),
    .B(\V3/V2/A1/A2/c3 ),
    .Z(\V3/V2/s1 [7]));
 OR2_X1 \V3/V2/A1/A2/M4/_0_  (.A1(\V3/V2/A1/A2/M4/c1 ),
    .A2(\V3/V2/A1/A2/M4/c2 ),
    .ZN(\V3/V2/c1 ));
 AND2_X1 \V3/V2/A2/A1/M1/M1/_0_  (.A1(\V3/V2/s1 [0]),
    .A2(\V3/V2/v1 [4]),
    .ZN(\V3/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M1/M1/_1_  (.A(\V3/V2/s1 [0]),
    .B(\V3/V2/v1 [4]),
    .Z(\V3/V2/A2/A1/M1/s1 ));
 AND2_X1 \V3/V2/A2/A1/M1/M2/_0_  (.A1(\V3/V2/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M1/M2/_1_  (.A(\V3/V2/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v2 [4]));
 OR2_X1 \V3/V2/A2/A1/M1/_0_  (.A1(\V3/V2/A2/A1/M1/c1 ),
    .A2(\V3/V2/A2/A1/M1/c2 ),
    .ZN(\V3/V2/A2/A1/c1 ));
 AND2_X1 \V3/V2/A2/A1/M2/M1/_0_  (.A1(\V3/V2/s1 [1]),
    .A2(\V3/V2/v1 [5]),
    .ZN(\V3/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M2/M1/_1_  (.A(\V3/V2/s1 [1]),
    .B(\V3/V2/v1 [5]),
    .Z(\V3/V2/A2/A1/M2/s1 ));
 AND2_X1 \V3/V2/A2/A1/M2/M2/_0_  (.A1(\V3/V2/A2/A1/M2/s1 ),
    .A2(\V3/V2/A2/A1/c1 ),
    .ZN(\V3/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M2/M2/_1_  (.A(\V3/V2/A2/A1/M2/s1 ),
    .B(\V3/V2/A2/A1/c1 ),
    .Z(\V3/v2 [5]));
 OR2_X1 \V3/V2/A2/A1/M2/_0_  (.A1(\V3/V2/A2/A1/M2/c1 ),
    .A2(\V3/V2/A2/A1/M2/c2 ),
    .ZN(\V3/V2/A2/A1/c2 ));
 AND2_X1 \V3/V2/A2/A1/M3/M1/_0_  (.A1(\V3/V2/s1 [2]),
    .A2(\V3/V2/v1 [6]),
    .ZN(\V3/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M3/M1/_1_  (.A(\V3/V2/s1 [2]),
    .B(\V3/V2/v1 [6]),
    .Z(\V3/V2/A2/A1/M3/s1 ));
 AND2_X1 \V3/V2/A2/A1/M3/M2/_0_  (.A1(\V3/V2/A2/A1/M3/s1 ),
    .A2(\V3/V2/A2/A1/c2 ),
    .ZN(\V3/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M3/M2/_1_  (.A(\V3/V2/A2/A1/M3/s1 ),
    .B(\V3/V2/A2/A1/c2 ),
    .Z(\V3/v2 [6]));
 OR2_X1 \V3/V2/A2/A1/M3/_0_  (.A1(\V3/V2/A2/A1/M3/c1 ),
    .A2(\V3/V2/A2/A1/M3/c2 ),
    .ZN(\V3/V2/A2/A1/c3 ));
 AND2_X1 \V3/V2/A2/A1/M4/M1/_0_  (.A1(\V3/V2/s1 [3]),
    .A2(\V3/V2/v1 [7]),
    .ZN(\V3/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M4/M1/_1_  (.A(\V3/V2/s1 [3]),
    .B(\V3/V2/v1 [7]),
    .Z(\V3/V2/A2/A1/M4/s1 ));
 AND2_X1 \V3/V2/A2/A1/M4/M2/_0_  (.A1(\V3/V2/A2/A1/M4/s1 ),
    .A2(\V3/V2/A2/A1/c3 ),
    .ZN(\V3/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M4/M2/_1_  (.A(\V3/V2/A2/A1/M4/s1 ),
    .B(\V3/V2/A2/A1/c3 ),
    .Z(\V3/v2 [7]));
 OR2_X1 \V3/V2/A2/A1/M4/_0_  (.A1(\V3/V2/A2/A1/M4/c1 ),
    .A2(\V3/V2/A2/A1/M4/c2 ),
    .ZN(\V3/V2/A2/c1 ));
 AND2_X1 \V3/V2/A2/A2/M1/M1/_0_  (.A1(\V3/V2/s1 [4]),
    .A2(ground),
    .ZN(\V3/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M1/M1/_1_  (.A(\V3/V2/s1 [4]),
    .B(ground),
    .Z(\V3/V2/A2/A2/M1/s1 ));
 AND2_X1 \V3/V2/A2/A2/M1/M2/_0_  (.A1(\V3/V2/A2/A2/M1/s1 ),
    .A2(\V3/V2/A2/c1 ),
    .ZN(\V3/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M1/M2/_1_  (.A(\V3/V2/A2/A2/M1/s1 ),
    .B(\V3/V2/A2/c1 ),
    .Z(\V3/V2/s2 [4]));
 OR2_X1 \V3/V2/A2/A2/M1/_0_  (.A1(\V3/V2/A2/A2/M1/c1 ),
    .A2(\V3/V2/A2/A2/M1/c2 ),
    .ZN(\V3/V2/A2/A2/c1 ));
 AND2_X1 \V3/V2/A2/A2/M2/M1/_0_  (.A1(\V3/V2/s1 [5]),
    .A2(ground),
    .ZN(\V3/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M2/M1/_1_  (.A(\V3/V2/s1 [5]),
    .B(ground),
    .Z(\V3/V2/A2/A2/M2/s1 ));
 AND2_X1 \V3/V2/A2/A2/M2/M2/_0_  (.A1(\V3/V2/A2/A2/M2/s1 ),
    .A2(\V3/V2/A2/A2/c1 ),
    .ZN(\V3/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M2/M2/_1_  (.A(\V3/V2/A2/A2/M2/s1 ),
    .B(\V3/V2/A2/A2/c1 ),
    .Z(\V3/V2/s2 [5]));
 OR2_X1 \V3/V2/A2/A2/M2/_0_  (.A1(\V3/V2/A2/A2/M2/c1 ),
    .A2(\V3/V2/A2/A2/M2/c2 ),
    .ZN(\V3/V2/A2/A2/c2 ));
 AND2_X1 \V3/V2/A2/A2/M3/M1/_0_  (.A1(\V3/V2/s1 [6]),
    .A2(ground),
    .ZN(\V3/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M3/M1/_1_  (.A(\V3/V2/s1 [6]),
    .B(ground),
    .Z(\V3/V2/A2/A2/M3/s1 ));
 AND2_X1 \V3/V2/A2/A2/M3/M2/_0_  (.A1(\V3/V2/A2/A2/M3/s1 ),
    .A2(\V3/V2/A2/A2/c2 ),
    .ZN(\V3/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M3/M2/_1_  (.A(\V3/V2/A2/A2/M3/s1 ),
    .B(\V3/V2/A2/A2/c2 ),
    .Z(\V3/V2/s2 [6]));
 OR2_X1 \V3/V2/A2/A2/M3/_0_  (.A1(\V3/V2/A2/A2/M3/c1 ),
    .A2(\V3/V2/A2/A2/M3/c2 ),
    .ZN(\V3/V2/A2/A2/c3 ));
 AND2_X1 \V3/V2/A2/A2/M4/M1/_0_  (.A1(\V3/V2/s1 [7]),
    .A2(ground),
    .ZN(\V3/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M4/M1/_1_  (.A(\V3/V2/s1 [7]),
    .B(ground),
    .Z(\V3/V2/A2/A2/M4/s1 ));
 AND2_X1 \V3/V2/A2/A2/M4/M2/_0_  (.A1(\V3/V2/A2/A2/M4/s1 ),
    .A2(\V3/V2/A2/A2/c3 ),
    .ZN(\V3/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M4/M2/_1_  (.A(\V3/V2/A2/A2/M4/s1 ),
    .B(\V3/V2/A2/A2/c3 ),
    .Z(\V3/V2/s2 [7]));
 OR2_X1 \V3/V2/A2/A2/M4/_0_  (.A1(\V3/V2/A2/A2/M4/c1 ),
    .A2(\V3/V2/A2/A2/M4/c2 ),
    .ZN(\V3/V2/c2 ));
 AND2_X1 \V3/V2/A3/A1/M1/M1/_0_  (.A1(\V3/V2/v4 [0]),
    .A2(\V3/V2/s2 [4]),
    .ZN(\V3/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M1/M1/_1_  (.A(\V3/V2/v4 [0]),
    .B(\V3/V2/s2 [4]),
    .Z(\V3/V2/A3/A1/M1/s1 ));
 AND2_X1 \V3/V2/A3/A1/M1/M2/_0_  (.A1(\V3/V2/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M1/M2/_1_  (.A(\V3/V2/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v2 [8]));
 OR2_X1 \V3/V2/A3/A1/M1/_0_  (.A1(\V3/V2/A3/A1/M1/c1 ),
    .A2(\V3/V2/A3/A1/M1/c2 ),
    .ZN(\V3/V2/A3/A1/c1 ));
 AND2_X1 \V3/V2/A3/A1/M2/M1/_0_  (.A1(\V3/V2/v4 [1]),
    .A2(\V3/V2/s2 [5]),
    .ZN(\V3/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M2/M1/_1_  (.A(\V3/V2/v4 [1]),
    .B(\V3/V2/s2 [5]),
    .Z(\V3/V2/A3/A1/M2/s1 ));
 AND2_X1 \V3/V2/A3/A1/M2/M2/_0_  (.A1(\V3/V2/A3/A1/M2/s1 ),
    .A2(\V3/V2/A3/A1/c1 ),
    .ZN(\V3/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M2/M2/_1_  (.A(\V3/V2/A3/A1/M2/s1 ),
    .B(\V3/V2/A3/A1/c1 ),
    .Z(\V3/v2 [9]));
 OR2_X1 \V3/V2/A3/A1/M2/_0_  (.A1(\V3/V2/A3/A1/M2/c1 ),
    .A2(\V3/V2/A3/A1/M2/c2 ),
    .ZN(\V3/V2/A3/A1/c2 ));
 AND2_X1 \V3/V2/A3/A1/M3/M1/_0_  (.A1(\V3/V2/v4 [2]),
    .A2(\V3/V2/s2 [6]),
    .ZN(\V3/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M3/M1/_1_  (.A(\V3/V2/v4 [2]),
    .B(\V3/V2/s2 [6]),
    .Z(\V3/V2/A3/A1/M3/s1 ));
 AND2_X1 \V3/V2/A3/A1/M3/M2/_0_  (.A1(\V3/V2/A3/A1/M3/s1 ),
    .A2(\V3/V2/A3/A1/c2 ),
    .ZN(\V3/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M3/M2/_1_  (.A(\V3/V2/A3/A1/M3/s1 ),
    .B(\V3/V2/A3/A1/c2 ),
    .Z(\V3/v2 [10]));
 OR2_X1 \V3/V2/A3/A1/M3/_0_  (.A1(\V3/V2/A3/A1/M3/c1 ),
    .A2(\V3/V2/A3/A1/M3/c2 ),
    .ZN(\V3/V2/A3/A1/c3 ));
 AND2_X1 \V3/V2/A3/A1/M4/M1/_0_  (.A1(\V3/V2/v4 [3]),
    .A2(\V3/V2/s2 [7]),
    .ZN(\V3/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M4/M1/_1_  (.A(\V3/V2/v4 [3]),
    .B(\V3/V2/s2 [7]),
    .Z(\V3/V2/A3/A1/M4/s1 ));
 AND2_X1 \V3/V2/A3/A1/M4/M2/_0_  (.A1(\V3/V2/A3/A1/M4/s1 ),
    .A2(\V3/V2/A3/A1/c3 ),
    .ZN(\V3/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M4/M2/_1_  (.A(\V3/V2/A3/A1/M4/s1 ),
    .B(\V3/V2/A3/A1/c3 ),
    .Z(\V3/v2 [11]));
 OR2_X1 \V3/V2/A3/A1/M4/_0_  (.A1(\V3/V2/A3/A1/M4/c1 ),
    .A2(\V3/V2/A3/A1/M4/c2 ),
    .ZN(\V3/V2/A3/c1 ));
 AND2_X1 \V3/V2/A3/A2/M1/M1/_0_  (.A1(\V3/V2/v4 [4]),
    .A2(\V3/V2/c3 ),
    .ZN(\V3/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M1/M1/_1_  (.A(\V3/V2/v4 [4]),
    .B(\V3/V2/c3 ),
    .Z(\V3/V2/A3/A2/M1/s1 ));
 AND2_X1 \V3/V2/A3/A2/M1/M2/_0_  (.A1(\V3/V2/A3/A2/M1/s1 ),
    .A2(\V3/V2/A3/c1 ),
    .ZN(\V3/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M1/M2/_1_  (.A(\V3/V2/A3/A2/M1/s1 ),
    .B(\V3/V2/A3/c1 ),
    .Z(\V3/v2 [12]));
 OR2_X1 \V3/V2/A3/A2/M1/_0_  (.A1(\V3/V2/A3/A2/M1/c1 ),
    .A2(\V3/V2/A3/A2/M1/c2 ),
    .ZN(\V3/V2/A3/A2/c1 ));
 AND2_X1 \V3/V2/A3/A2/M2/M1/_0_  (.A1(\V3/V2/v4 [5]),
    .A2(ground),
    .ZN(\V3/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M2/M1/_1_  (.A(\V3/V2/v4 [5]),
    .B(ground),
    .Z(\V3/V2/A3/A2/M2/s1 ));
 AND2_X1 \V3/V2/A3/A2/M2/M2/_0_  (.A1(\V3/V2/A3/A2/M2/s1 ),
    .A2(\V3/V2/A3/A2/c1 ),
    .ZN(\V3/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M2/M2/_1_  (.A(\V3/V2/A3/A2/M2/s1 ),
    .B(\V3/V2/A3/A2/c1 ),
    .Z(\V3/v2 [13]));
 OR2_X1 \V3/V2/A3/A2/M2/_0_  (.A1(\V3/V2/A3/A2/M2/c1 ),
    .A2(\V3/V2/A3/A2/M2/c2 ),
    .ZN(\V3/V2/A3/A2/c2 ));
 AND2_X1 \V3/V2/A3/A2/M3/M1/_0_  (.A1(\V3/V2/v4 [6]),
    .A2(ground),
    .ZN(\V3/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M3/M1/_1_  (.A(\V3/V2/v4 [6]),
    .B(ground),
    .Z(\V3/V2/A3/A2/M3/s1 ));
 AND2_X1 \V3/V2/A3/A2/M3/M2/_0_  (.A1(\V3/V2/A3/A2/M3/s1 ),
    .A2(\V3/V2/A3/A2/c2 ),
    .ZN(\V3/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M3/M2/_1_  (.A(\V3/V2/A3/A2/M3/s1 ),
    .B(\V3/V2/A3/A2/c2 ),
    .Z(\V3/v2 [14]));
 OR2_X1 \V3/V2/A3/A2/M3/_0_  (.A1(\V3/V2/A3/A2/M3/c1 ),
    .A2(\V3/V2/A3/A2/M3/c2 ),
    .ZN(\V3/V2/A3/A2/c3 ));
 AND2_X1 \V3/V2/A3/A2/M4/M1/_0_  (.A1(\V3/V2/v4 [7]),
    .A2(ground),
    .ZN(\V3/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M4/M1/_1_  (.A(\V3/V2/v4 [7]),
    .B(ground),
    .Z(\V3/V2/A3/A2/M4/s1 ));
 AND2_X1 \V3/V2/A3/A2/M4/M2/_0_  (.A1(\V3/V2/A3/A2/M4/s1 ),
    .A2(\V3/V2/A3/A2/c3 ),
    .ZN(\V3/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M4/M2/_1_  (.A(\V3/V2/A3/A2/M4/s1 ),
    .B(\V3/V2/A3/A2/c3 ),
    .Z(\V3/v2 [15]));
 OR2_X1 \V3/V2/A3/A2/M4/_0_  (.A1(\V3/V2/A3/A2/M4/c1 ),
    .A2(\V3/V2/A3/A2/M4/c2 ),
    .ZN(\V3/V2/overflow ));
 AND2_X1 \V3/V2/V1/A1/M1/M1/_0_  (.A1(\V3/V2/V1/v2 [0]),
    .A2(\V3/V2/V1/v3 [0]),
    .ZN(\V3/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M1/M1/_1_  (.A(\V3/V2/V1/v2 [0]),
    .B(\V3/V2/V1/v3 [0]),
    .Z(\V3/V2/V1/A1/M1/s1 ));
 AND2_X1 \V3/V2/V1/A1/M1/M2/_0_  (.A1(\V3/V2/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M1/M2/_1_  (.A(\V3/V2/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/V1/s1 [0]));
 OR2_X1 \V3/V2/V1/A1/M1/_0_  (.A1(\V3/V2/V1/A1/M1/c1 ),
    .A2(\V3/V2/V1/A1/M1/c2 ),
    .ZN(\V3/V2/V1/A1/c1 ));
 AND2_X1 \V3/V2/V1/A1/M2/M1/_0_  (.A1(\V3/V2/V1/v2 [1]),
    .A2(\V3/V2/V1/v3 [1]),
    .ZN(\V3/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M2/M1/_1_  (.A(\V3/V2/V1/v2 [1]),
    .B(\V3/V2/V1/v3 [1]),
    .Z(\V3/V2/V1/A1/M2/s1 ));
 AND2_X1 \V3/V2/V1/A1/M2/M2/_0_  (.A1(\V3/V2/V1/A1/M2/s1 ),
    .A2(\V3/V2/V1/A1/c1 ),
    .ZN(\V3/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M2/M2/_1_  (.A(\V3/V2/V1/A1/M2/s1 ),
    .B(\V3/V2/V1/A1/c1 ),
    .Z(\V3/V2/V1/s1 [1]));
 OR2_X1 \V3/V2/V1/A1/M2/_0_  (.A1(\V3/V2/V1/A1/M2/c1 ),
    .A2(\V3/V2/V1/A1/M2/c2 ),
    .ZN(\V3/V2/V1/A1/c2 ));
 AND2_X1 \V3/V2/V1/A1/M3/M1/_0_  (.A1(\V3/V2/V1/v2 [2]),
    .A2(\V3/V2/V1/v3 [2]),
    .ZN(\V3/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M3/M1/_1_  (.A(\V3/V2/V1/v2 [2]),
    .B(\V3/V2/V1/v3 [2]),
    .Z(\V3/V2/V1/A1/M3/s1 ));
 AND2_X1 \V3/V2/V1/A1/M3/M2/_0_  (.A1(\V3/V2/V1/A1/M3/s1 ),
    .A2(\V3/V2/V1/A1/c2 ),
    .ZN(\V3/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M3/M2/_1_  (.A(\V3/V2/V1/A1/M3/s1 ),
    .B(\V3/V2/V1/A1/c2 ),
    .Z(\V3/V2/V1/s1 [2]));
 OR2_X1 \V3/V2/V1/A1/M3/_0_  (.A1(\V3/V2/V1/A1/M3/c1 ),
    .A2(\V3/V2/V1/A1/M3/c2 ),
    .ZN(\V3/V2/V1/A1/c3 ));
 AND2_X1 \V3/V2/V1/A1/M4/M1/_0_  (.A1(\V3/V2/V1/v2 [3]),
    .A2(\V3/V2/V1/v3 [3]),
    .ZN(\V3/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M4/M1/_1_  (.A(\V3/V2/V1/v2 [3]),
    .B(\V3/V2/V1/v3 [3]),
    .Z(\V3/V2/V1/A1/M4/s1 ));
 AND2_X1 \V3/V2/V1/A1/M4/M2/_0_  (.A1(\V3/V2/V1/A1/M4/s1 ),
    .A2(\V3/V2/V1/A1/c3 ),
    .ZN(\V3/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M4/M2/_1_  (.A(\V3/V2/V1/A1/M4/s1 ),
    .B(\V3/V2/V1/A1/c3 ),
    .Z(\V3/V2/V1/s1 [3]));
 OR2_X1 \V3/V2/V1/A1/M4/_0_  (.A1(\V3/V2/V1/A1/M4/c1 ),
    .A2(\V3/V2/V1/A1/M4/c2 ),
    .ZN(\V3/V2/V1/c1 ));
 AND2_X1 \V3/V2/V1/A2/M1/M1/_0_  (.A1(\V3/V2/V1/s1 [0]),
    .A2(\V3/V2/V1/v1 [2]),
    .ZN(\V3/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M1/M1/_1_  (.A(\V3/V2/V1/s1 [0]),
    .B(\V3/V2/V1/v1 [2]),
    .Z(\V3/V2/V1/A2/M1/s1 ));
 AND2_X1 \V3/V2/V1/A2/M1/M2/_0_  (.A1(\V3/V2/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M1/M2/_1_  (.A(\V3/V2/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/v2 [2]));
 OR2_X1 \V3/V2/V1/A2/M1/_0_  (.A1(\V3/V2/V1/A2/M1/c1 ),
    .A2(\V3/V2/V1/A2/M1/c2 ),
    .ZN(\V3/V2/V1/A2/c1 ));
 AND2_X1 \V3/V2/V1/A2/M2/M1/_0_  (.A1(\V3/V2/V1/s1 [1]),
    .A2(\V3/V2/V1/v1 [3]),
    .ZN(\V3/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M2/M1/_1_  (.A(\V3/V2/V1/s1 [1]),
    .B(\V3/V2/V1/v1 [3]),
    .Z(\V3/V2/V1/A2/M2/s1 ));
 AND2_X1 \V3/V2/V1/A2/M2/M2/_0_  (.A1(\V3/V2/V1/A2/M2/s1 ),
    .A2(\V3/V2/V1/A2/c1 ),
    .ZN(\V3/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M2/M2/_1_  (.A(\V3/V2/V1/A2/M2/s1 ),
    .B(\V3/V2/V1/A2/c1 ),
    .Z(\V3/v2 [3]));
 OR2_X1 \V3/V2/V1/A2/M2/_0_  (.A1(\V3/V2/V1/A2/M2/c1 ),
    .A2(\V3/V2/V1/A2/M2/c2 ),
    .ZN(\V3/V2/V1/A2/c2 ));
 AND2_X1 \V3/V2/V1/A2/M3/M1/_0_  (.A1(\V3/V2/V1/s1 [2]),
    .A2(ground),
    .ZN(\V3/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M3/M1/_1_  (.A(\V3/V2/V1/s1 [2]),
    .B(ground),
    .Z(\V3/V2/V1/A2/M3/s1 ));
 AND2_X1 \V3/V2/V1/A2/M3/M2/_0_  (.A1(\V3/V2/V1/A2/M3/s1 ),
    .A2(\V3/V2/V1/A2/c2 ),
    .ZN(\V3/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M3/M2/_1_  (.A(\V3/V2/V1/A2/M3/s1 ),
    .B(\V3/V2/V1/A2/c2 ),
    .Z(\V3/V2/V1/s2 [2]));
 OR2_X1 \V3/V2/V1/A2/M3/_0_  (.A1(\V3/V2/V1/A2/M3/c1 ),
    .A2(\V3/V2/V1/A2/M3/c2 ),
    .ZN(\V3/V2/V1/A2/c3 ));
 AND2_X1 \V3/V2/V1/A2/M4/M1/_0_  (.A1(\V3/V2/V1/s1 [3]),
    .A2(ground),
    .ZN(\V3/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M4/M1/_1_  (.A(\V3/V2/V1/s1 [3]),
    .B(ground),
    .Z(\V3/V2/V1/A2/M4/s1 ));
 AND2_X1 \V3/V2/V1/A2/M4/M2/_0_  (.A1(\V3/V2/V1/A2/M4/s1 ),
    .A2(\V3/V2/V1/A2/c3 ),
    .ZN(\V3/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M4/M2/_1_  (.A(\V3/V2/V1/A2/M4/s1 ),
    .B(\V3/V2/V1/A2/c3 ),
    .Z(\V3/V2/V1/s2 [3]));
 OR2_X1 \V3/V2/V1/A2/M4/_0_  (.A1(\V3/V2/V1/A2/M4/c1 ),
    .A2(\V3/V2/V1/A2/M4/c2 ),
    .ZN(\V3/V2/V1/c2 ));
 AND2_X1 \V3/V2/V1/A3/M1/M1/_0_  (.A1(\V3/V2/V1/v4 [0]),
    .A2(\V3/V2/V1/s2 [2]),
    .ZN(\V3/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M1/M1/_1_  (.A(\V3/V2/V1/v4 [0]),
    .B(\V3/V2/V1/s2 [2]),
    .Z(\V3/V2/V1/A3/M1/s1 ));
 AND2_X1 \V3/V2/V1/A3/M1/M2/_0_  (.A1(\V3/V2/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M1/M2/_1_  (.A(\V3/V2/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v1 [4]));
 OR2_X1 \V3/V2/V1/A3/M1/_0_  (.A1(\V3/V2/V1/A3/M1/c1 ),
    .A2(\V3/V2/V1/A3/M1/c2 ),
    .ZN(\V3/V2/V1/A3/c1 ));
 AND2_X1 \V3/V2/V1/A3/M2/M1/_0_  (.A1(\V3/V2/V1/v4 [1]),
    .A2(\V3/V2/V1/s2 [3]),
    .ZN(\V3/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M2/M1/_1_  (.A(\V3/V2/V1/v4 [1]),
    .B(\V3/V2/V1/s2 [3]),
    .Z(\V3/V2/V1/A3/M2/s1 ));
 AND2_X1 \V3/V2/V1/A3/M2/M2/_0_  (.A1(\V3/V2/V1/A3/M2/s1 ),
    .A2(\V3/V2/V1/A3/c1 ),
    .ZN(\V3/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M2/M2/_1_  (.A(\V3/V2/V1/A3/M2/s1 ),
    .B(\V3/V2/V1/A3/c1 ),
    .Z(\V3/V2/v1 [5]));
 OR2_X1 \V3/V2/V1/A3/M2/_0_  (.A1(\V3/V2/V1/A3/M2/c1 ),
    .A2(\V3/V2/V1/A3/M2/c2 ),
    .ZN(\V3/V2/V1/A3/c2 ));
 AND2_X1 \V3/V2/V1/A3/M3/M1/_0_  (.A1(\V3/V2/V1/v4 [2]),
    .A2(\V3/V2/V1/c3 ),
    .ZN(\V3/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M3/M1/_1_  (.A(\V3/V2/V1/v4 [2]),
    .B(\V3/V2/V1/c3 ),
    .Z(\V3/V2/V1/A3/M3/s1 ));
 AND2_X1 \V3/V2/V1/A3/M3/M2/_0_  (.A1(\V3/V2/V1/A3/M3/s1 ),
    .A2(\V3/V2/V1/A3/c2 ),
    .ZN(\V3/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M3/M2/_1_  (.A(\V3/V2/V1/A3/M3/s1 ),
    .B(\V3/V2/V1/A3/c2 ),
    .Z(\V3/V2/v1 [6]));
 OR2_X1 \V3/V2/V1/A3/M3/_0_  (.A1(\V3/V2/V1/A3/M3/c1 ),
    .A2(\V3/V2/V1/A3/M3/c2 ),
    .ZN(\V3/V2/V1/A3/c3 ));
 AND2_X1 \V3/V2/V1/A3/M4/M1/_0_  (.A1(\V3/V2/V1/v4 [3]),
    .A2(ground),
    .ZN(\V3/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M4/M1/_1_  (.A(\V3/V2/V1/v4 [3]),
    .B(ground),
    .Z(\V3/V2/V1/A3/M4/s1 ));
 AND2_X1 \V3/V2/V1/A3/M4/M2/_0_  (.A1(\V3/V2/V1/A3/M4/s1 ),
    .A2(\V3/V2/V1/A3/c3 ),
    .ZN(\V3/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M4/M2/_1_  (.A(\V3/V2/V1/A3/M4/s1 ),
    .B(\V3/V2/V1/A3/c3 ),
    .Z(\V3/V2/v1 [7]));
 OR2_X1 \V3/V2/V1/A3/M4/_0_  (.A1(\V3/V2/V1/A3/M4/c1 ),
    .A2(\V3/V2/V1/A3/M4/c2 ),
    .ZN(\V3/V2/V1/overflow ));
 AND2_X1 \V3/V2/V1/V1/HA1/_0_  (.A1(\V3/V2/V1/V1/w2 ),
    .A2(\V3/V2/V1/V1/w1 ),
    .ZN(\V3/V2/V1/V1/w4 ));
 XOR2_X2 \V3/V2/V1/V1/HA1/_1_  (.A(\V3/V2/V1/V1/w2 ),
    .B(\V3/V2/V1/V1/w1 ),
    .Z(\V3/v2 [1]));
 AND2_X1 \V3/V2/V1/V1/HA2/_0_  (.A1(\V3/V2/V1/V1/w4 ),
    .A2(\V3/V2/V1/V1/w3 ),
    .ZN(\V3/V2/V1/v1 [3]));
 XOR2_X2 \V3/V2/V1/V1/HA2/_1_  (.A(\V3/V2/V1/V1/w4 ),
    .B(\V3/V2/V1/V1/w3 ),
    .Z(\V3/V2/V1/v1 [2]));
 AND2_X1 \V3/V2/V1/V1/_0_  (.A1(A[8]),
    .A2(B[16]),
    .ZN(\V3/v2 [0]));
 AND2_X1 \V3/V2/V1/V1/_1_  (.A1(A[8]),
    .A2(B[17]),
    .ZN(\V3/V2/V1/V1/w1 ));
 AND2_X1 \V3/V2/V1/V1/_2_  (.A1(B[16]),
    .A2(A[9]),
    .ZN(\V3/V2/V1/V1/w2 ));
 AND2_X1 \V3/V2/V1/V1/_3_  (.A1(B[17]),
    .A2(A[9]),
    .ZN(\V3/V2/V1/V1/w3 ));
 AND2_X1 \V3/V2/V1/V2/HA1/_0_  (.A1(\V3/V2/V1/V2/w2 ),
    .A2(\V3/V2/V1/V2/w1 ),
    .ZN(\V3/V2/V1/V2/w4 ));
 XOR2_X2 \V3/V2/V1/V2/HA1/_1_  (.A(\V3/V2/V1/V2/w2 ),
    .B(\V3/V2/V1/V2/w1 ),
    .Z(\V3/V2/V1/v2 [1]));
 AND2_X1 \V3/V2/V1/V2/HA2/_0_  (.A1(\V3/V2/V1/V2/w4 ),
    .A2(\V3/V2/V1/V2/w3 ),
    .ZN(\V3/V2/V1/v2 [3]));
 XOR2_X2 \V3/V2/V1/V2/HA2/_1_  (.A(\V3/V2/V1/V2/w4 ),
    .B(\V3/V2/V1/V2/w3 ),
    .Z(\V3/V2/V1/v2 [2]));
 AND2_X1 \V3/V2/V1/V2/_0_  (.A1(A[10]),
    .A2(B[16]),
    .ZN(\V3/V2/V1/v2 [0]));
 AND2_X1 \V3/V2/V1/V2/_1_  (.A1(A[10]),
    .A2(B[17]),
    .ZN(\V3/V2/V1/V2/w1 ));
 AND2_X1 \V3/V2/V1/V2/_2_  (.A1(B[16]),
    .A2(A[11]),
    .ZN(\V3/V2/V1/V2/w2 ));
 AND2_X1 \V3/V2/V1/V2/_3_  (.A1(B[17]),
    .A2(A[11]),
    .ZN(\V3/V2/V1/V2/w3 ));
 AND2_X1 \V3/V2/V1/V3/HA1/_0_  (.A1(\V3/V2/V1/V3/w2 ),
    .A2(\V3/V2/V1/V3/w1 ),
    .ZN(\V3/V2/V1/V3/w4 ));
 XOR2_X2 \V3/V2/V1/V3/HA1/_1_  (.A(\V3/V2/V1/V3/w2 ),
    .B(\V3/V2/V1/V3/w1 ),
    .Z(\V3/V2/V1/v3 [1]));
 AND2_X1 \V3/V2/V1/V3/HA2/_0_  (.A1(\V3/V2/V1/V3/w4 ),
    .A2(\V3/V2/V1/V3/w3 ),
    .ZN(\V3/V2/V1/v3 [3]));
 XOR2_X2 \V3/V2/V1/V3/HA2/_1_  (.A(\V3/V2/V1/V3/w4 ),
    .B(\V3/V2/V1/V3/w3 ),
    .Z(\V3/V2/V1/v3 [2]));
 AND2_X1 \V3/V2/V1/V3/_0_  (.A1(A[8]),
    .A2(B[18]),
    .ZN(\V3/V2/V1/v3 [0]));
 AND2_X1 \V3/V2/V1/V3/_1_  (.A1(A[8]),
    .A2(B[19]),
    .ZN(\V3/V2/V1/V3/w1 ));
 AND2_X1 \V3/V2/V1/V3/_2_  (.A1(B[18]),
    .A2(A[9]),
    .ZN(\V3/V2/V1/V3/w2 ));
 AND2_X1 \V3/V2/V1/V3/_3_  (.A1(B[19]),
    .A2(A[9]),
    .ZN(\V3/V2/V1/V3/w3 ));
 AND2_X1 \V3/V2/V1/V4/HA1/_0_  (.A1(\V3/V2/V1/V4/w2 ),
    .A2(\V3/V2/V1/V4/w1 ),
    .ZN(\V3/V2/V1/V4/w4 ));
 XOR2_X2 \V3/V2/V1/V4/HA1/_1_  (.A(\V3/V2/V1/V4/w2 ),
    .B(\V3/V2/V1/V4/w1 ),
    .Z(\V3/V2/V1/v4 [1]));
 AND2_X1 \V3/V2/V1/V4/HA2/_0_  (.A1(\V3/V2/V1/V4/w4 ),
    .A2(\V3/V2/V1/V4/w3 ),
    .ZN(\V3/V2/V1/v4 [3]));
 XOR2_X2 \V3/V2/V1/V4/HA2/_1_  (.A(\V3/V2/V1/V4/w4 ),
    .B(\V3/V2/V1/V4/w3 ),
    .Z(\V3/V2/V1/v4 [2]));
 AND2_X1 \V3/V2/V1/V4/_0_  (.A1(A[10]),
    .A2(B[18]),
    .ZN(\V3/V2/V1/v4 [0]));
 AND2_X1 \V3/V2/V1/V4/_1_  (.A1(A[10]),
    .A2(B[19]),
    .ZN(\V3/V2/V1/V4/w1 ));
 AND2_X1 \V3/V2/V1/V4/_2_  (.A1(B[18]),
    .A2(A[11]),
    .ZN(\V3/V2/V1/V4/w2 ));
 AND2_X1 \V3/V2/V1/V4/_3_  (.A1(B[19]),
    .A2(A[11]),
    .ZN(\V3/V2/V1/V4/w3 ));
 OR2_X1 \V3/V2/V1/_0_  (.A1(\V3/V2/V1/c1 ),
    .A2(\V3/V2/V1/c2 ),
    .ZN(\V3/V2/V1/c3 ));
 AND2_X1 \V3/V2/V2/A1/M1/M1/_0_  (.A1(\V3/V2/V2/v2 [0]),
    .A2(\V3/V2/V2/v3 [0]),
    .ZN(\V3/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M1/M1/_1_  (.A(\V3/V2/V2/v2 [0]),
    .B(\V3/V2/V2/v3 [0]),
    .Z(\V3/V2/V2/A1/M1/s1 ));
 AND2_X1 \V3/V2/V2/A1/M1/M2/_0_  (.A1(\V3/V2/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M1/M2/_1_  (.A(\V3/V2/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/V2/s1 [0]));
 OR2_X1 \V3/V2/V2/A1/M1/_0_  (.A1(\V3/V2/V2/A1/M1/c1 ),
    .A2(\V3/V2/V2/A1/M1/c2 ),
    .ZN(\V3/V2/V2/A1/c1 ));
 AND2_X1 \V3/V2/V2/A1/M2/M1/_0_  (.A1(\V3/V2/V2/v2 [1]),
    .A2(\V3/V2/V2/v3 [1]),
    .ZN(\V3/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M2/M1/_1_  (.A(\V3/V2/V2/v2 [1]),
    .B(\V3/V2/V2/v3 [1]),
    .Z(\V3/V2/V2/A1/M2/s1 ));
 AND2_X1 \V3/V2/V2/A1/M2/M2/_0_  (.A1(\V3/V2/V2/A1/M2/s1 ),
    .A2(\V3/V2/V2/A1/c1 ),
    .ZN(\V3/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M2/M2/_1_  (.A(\V3/V2/V2/A1/M2/s1 ),
    .B(\V3/V2/V2/A1/c1 ),
    .Z(\V3/V2/V2/s1 [1]));
 OR2_X1 \V3/V2/V2/A1/M2/_0_  (.A1(\V3/V2/V2/A1/M2/c1 ),
    .A2(\V3/V2/V2/A1/M2/c2 ),
    .ZN(\V3/V2/V2/A1/c2 ));
 AND2_X1 \V3/V2/V2/A1/M3/M1/_0_  (.A1(\V3/V2/V2/v2 [2]),
    .A2(\V3/V2/V2/v3 [2]),
    .ZN(\V3/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M3/M1/_1_  (.A(\V3/V2/V2/v2 [2]),
    .B(\V3/V2/V2/v3 [2]),
    .Z(\V3/V2/V2/A1/M3/s1 ));
 AND2_X1 \V3/V2/V2/A1/M3/M2/_0_  (.A1(\V3/V2/V2/A1/M3/s1 ),
    .A2(\V3/V2/V2/A1/c2 ),
    .ZN(\V3/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M3/M2/_1_  (.A(\V3/V2/V2/A1/M3/s1 ),
    .B(\V3/V2/V2/A1/c2 ),
    .Z(\V3/V2/V2/s1 [2]));
 OR2_X1 \V3/V2/V2/A1/M3/_0_  (.A1(\V3/V2/V2/A1/M3/c1 ),
    .A2(\V3/V2/V2/A1/M3/c2 ),
    .ZN(\V3/V2/V2/A1/c3 ));
 AND2_X1 \V3/V2/V2/A1/M4/M1/_0_  (.A1(\V3/V2/V2/v2 [3]),
    .A2(\V3/V2/V2/v3 [3]),
    .ZN(\V3/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M4/M1/_1_  (.A(\V3/V2/V2/v2 [3]),
    .B(\V3/V2/V2/v3 [3]),
    .Z(\V3/V2/V2/A1/M4/s1 ));
 AND2_X1 \V3/V2/V2/A1/M4/M2/_0_  (.A1(\V3/V2/V2/A1/M4/s1 ),
    .A2(\V3/V2/V2/A1/c3 ),
    .ZN(\V3/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M4/M2/_1_  (.A(\V3/V2/V2/A1/M4/s1 ),
    .B(\V3/V2/V2/A1/c3 ),
    .Z(\V3/V2/V2/s1 [3]));
 OR2_X1 \V3/V2/V2/A1/M4/_0_  (.A1(\V3/V2/V2/A1/M4/c1 ),
    .A2(\V3/V2/V2/A1/M4/c2 ),
    .ZN(\V3/V2/V2/c1 ));
 AND2_X1 \V3/V2/V2/A2/M1/M1/_0_  (.A1(\V3/V2/V2/s1 [0]),
    .A2(\V3/V2/V2/v1 [2]),
    .ZN(\V3/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M1/M1/_1_  (.A(\V3/V2/V2/s1 [0]),
    .B(\V3/V2/V2/v1 [2]),
    .Z(\V3/V2/V2/A2/M1/s1 ));
 AND2_X1 \V3/V2/V2/A2/M1/M2/_0_  (.A1(\V3/V2/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M1/M2/_1_  (.A(\V3/V2/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v2 [2]));
 OR2_X1 \V3/V2/V2/A2/M1/_0_  (.A1(\V3/V2/V2/A2/M1/c1 ),
    .A2(\V3/V2/V2/A2/M1/c2 ),
    .ZN(\V3/V2/V2/A2/c1 ));
 AND2_X1 \V3/V2/V2/A2/M2/M1/_0_  (.A1(\V3/V2/V2/s1 [1]),
    .A2(\V3/V2/V2/v1 [3]),
    .ZN(\V3/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M2/M1/_1_  (.A(\V3/V2/V2/s1 [1]),
    .B(\V3/V2/V2/v1 [3]),
    .Z(\V3/V2/V2/A2/M2/s1 ));
 AND2_X1 \V3/V2/V2/A2/M2/M2/_0_  (.A1(\V3/V2/V2/A2/M2/s1 ),
    .A2(\V3/V2/V2/A2/c1 ),
    .ZN(\V3/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M2/M2/_1_  (.A(\V3/V2/V2/A2/M2/s1 ),
    .B(\V3/V2/V2/A2/c1 ),
    .Z(\V3/V2/v2 [3]));
 OR2_X1 \V3/V2/V2/A2/M2/_0_  (.A1(\V3/V2/V2/A2/M2/c1 ),
    .A2(\V3/V2/V2/A2/M2/c2 ),
    .ZN(\V3/V2/V2/A2/c2 ));
 AND2_X1 \V3/V2/V2/A2/M3/M1/_0_  (.A1(\V3/V2/V2/s1 [2]),
    .A2(ground),
    .ZN(\V3/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M3/M1/_1_  (.A(\V3/V2/V2/s1 [2]),
    .B(ground),
    .Z(\V3/V2/V2/A2/M3/s1 ));
 AND2_X1 \V3/V2/V2/A2/M3/M2/_0_  (.A1(\V3/V2/V2/A2/M3/s1 ),
    .A2(\V3/V2/V2/A2/c2 ),
    .ZN(\V3/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M3/M2/_1_  (.A(\V3/V2/V2/A2/M3/s1 ),
    .B(\V3/V2/V2/A2/c2 ),
    .Z(\V3/V2/V2/s2 [2]));
 OR2_X1 \V3/V2/V2/A2/M3/_0_  (.A1(\V3/V2/V2/A2/M3/c1 ),
    .A2(\V3/V2/V2/A2/M3/c2 ),
    .ZN(\V3/V2/V2/A2/c3 ));
 AND2_X1 \V3/V2/V2/A2/M4/M1/_0_  (.A1(\V3/V2/V2/s1 [3]),
    .A2(ground),
    .ZN(\V3/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M4/M1/_1_  (.A(\V3/V2/V2/s1 [3]),
    .B(ground),
    .Z(\V3/V2/V2/A2/M4/s1 ));
 AND2_X1 \V3/V2/V2/A2/M4/M2/_0_  (.A1(\V3/V2/V2/A2/M4/s1 ),
    .A2(\V3/V2/V2/A2/c3 ),
    .ZN(\V3/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M4/M2/_1_  (.A(\V3/V2/V2/A2/M4/s1 ),
    .B(\V3/V2/V2/A2/c3 ),
    .Z(\V3/V2/V2/s2 [3]));
 OR2_X1 \V3/V2/V2/A2/M4/_0_  (.A1(\V3/V2/V2/A2/M4/c1 ),
    .A2(\V3/V2/V2/A2/M4/c2 ),
    .ZN(\V3/V2/V2/c2 ));
 AND2_X1 \V3/V2/V2/A3/M1/M1/_0_  (.A1(\V3/V2/V2/v4 [0]),
    .A2(\V3/V2/V2/s2 [2]),
    .ZN(\V3/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M1/M1/_1_  (.A(\V3/V2/V2/v4 [0]),
    .B(\V3/V2/V2/s2 [2]),
    .Z(\V3/V2/V2/A3/M1/s1 ));
 AND2_X1 \V3/V2/V2/A3/M1/M2/_0_  (.A1(\V3/V2/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M1/M2/_1_  (.A(\V3/V2/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v2 [4]));
 OR2_X1 \V3/V2/V2/A3/M1/_0_  (.A1(\V3/V2/V2/A3/M1/c1 ),
    .A2(\V3/V2/V2/A3/M1/c2 ),
    .ZN(\V3/V2/V2/A3/c1 ));
 AND2_X1 \V3/V2/V2/A3/M2/M1/_0_  (.A1(\V3/V2/V2/v4 [1]),
    .A2(\V3/V2/V2/s2 [3]),
    .ZN(\V3/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M2/M1/_1_  (.A(\V3/V2/V2/v4 [1]),
    .B(\V3/V2/V2/s2 [3]),
    .Z(\V3/V2/V2/A3/M2/s1 ));
 AND2_X1 \V3/V2/V2/A3/M2/M2/_0_  (.A1(\V3/V2/V2/A3/M2/s1 ),
    .A2(\V3/V2/V2/A3/c1 ),
    .ZN(\V3/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M2/M2/_1_  (.A(\V3/V2/V2/A3/M2/s1 ),
    .B(\V3/V2/V2/A3/c1 ),
    .Z(\V3/V2/v2 [5]));
 OR2_X1 \V3/V2/V2/A3/M2/_0_  (.A1(\V3/V2/V2/A3/M2/c1 ),
    .A2(\V3/V2/V2/A3/M2/c2 ),
    .ZN(\V3/V2/V2/A3/c2 ));
 AND2_X1 \V3/V2/V2/A3/M3/M1/_0_  (.A1(\V3/V2/V2/v4 [2]),
    .A2(\V3/V2/V2/c3 ),
    .ZN(\V3/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M3/M1/_1_  (.A(\V3/V2/V2/v4 [2]),
    .B(\V3/V2/V2/c3 ),
    .Z(\V3/V2/V2/A3/M3/s1 ));
 AND2_X1 \V3/V2/V2/A3/M3/M2/_0_  (.A1(\V3/V2/V2/A3/M3/s1 ),
    .A2(\V3/V2/V2/A3/c2 ),
    .ZN(\V3/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M3/M2/_1_  (.A(\V3/V2/V2/A3/M3/s1 ),
    .B(\V3/V2/V2/A3/c2 ),
    .Z(\V3/V2/v2 [6]));
 OR2_X1 \V3/V2/V2/A3/M3/_0_  (.A1(\V3/V2/V2/A3/M3/c1 ),
    .A2(\V3/V2/V2/A3/M3/c2 ),
    .ZN(\V3/V2/V2/A3/c3 ));
 AND2_X1 \V3/V2/V2/A3/M4/M1/_0_  (.A1(\V3/V2/V2/v4 [3]),
    .A2(ground),
    .ZN(\V3/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M4/M1/_1_  (.A(\V3/V2/V2/v4 [3]),
    .B(ground),
    .Z(\V3/V2/V2/A3/M4/s1 ));
 AND2_X1 \V3/V2/V2/A3/M4/M2/_0_  (.A1(\V3/V2/V2/A3/M4/s1 ),
    .A2(\V3/V2/V2/A3/c3 ),
    .ZN(\V3/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M4/M2/_1_  (.A(\V3/V2/V2/A3/M4/s1 ),
    .B(\V3/V2/V2/A3/c3 ),
    .Z(\V3/V2/v2 [7]));
 OR2_X1 \V3/V2/V2/A3/M4/_0_  (.A1(\V3/V2/V2/A3/M4/c1 ),
    .A2(\V3/V2/V2/A3/M4/c2 ),
    .ZN(\V3/V2/V2/overflow ));
 AND2_X1 \V3/V2/V2/V1/HA1/_0_  (.A1(\V3/V2/V2/V1/w2 ),
    .A2(\V3/V2/V2/V1/w1 ),
    .ZN(\V3/V2/V2/V1/w4 ));
 XOR2_X2 \V3/V2/V2/V1/HA1/_1_  (.A(\V3/V2/V2/V1/w2 ),
    .B(\V3/V2/V2/V1/w1 ),
    .Z(\V3/V2/v2 [1]));
 AND2_X1 \V3/V2/V2/V1/HA2/_0_  (.A1(\V3/V2/V2/V1/w4 ),
    .A2(\V3/V2/V2/V1/w3 ),
    .ZN(\V3/V2/V2/v1 [3]));
 XOR2_X2 \V3/V2/V2/V1/HA2/_1_  (.A(\V3/V2/V2/V1/w4 ),
    .B(\V3/V2/V2/V1/w3 ),
    .Z(\V3/V2/V2/v1 [2]));
 AND2_X1 \V3/V2/V2/V1/_0_  (.A1(A[12]),
    .A2(B[16]),
    .ZN(\V3/V2/v2 [0]));
 AND2_X1 \V3/V2/V2/V1/_1_  (.A1(A[12]),
    .A2(B[17]),
    .ZN(\V3/V2/V2/V1/w1 ));
 AND2_X1 \V3/V2/V2/V1/_2_  (.A1(B[16]),
    .A2(A[13]),
    .ZN(\V3/V2/V2/V1/w2 ));
 AND2_X1 \V3/V2/V2/V1/_3_  (.A1(B[17]),
    .A2(A[13]),
    .ZN(\V3/V2/V2/V1/w3 ));
 AND2_X1 \V3/V2/V2/V2/HA1/_0_  (.A1(\V3/V2/V2/V2/w2 ),
    .A2(\V3/V2/V2/V2/w1 ),
    .ZN(\V3/V2/V2/V2/w4 ));
 XOR2_X2 \V3/V2/V2/V2/HA1/_1_  (.A(\V3/V2/V2/V2/w2 ),
    .B(\V3/V2/V2/V2/w1 ),
    .Z(\V3/V2/V2/v2 [1]));
 AND2_X1 \V3/V2/V2/V2/HA2/_0_  (.A1(\V3/V2/V2/V2/w4 ),
    .A2(\V3/V2/V2/V2/w3 ),
    .ZN(\V3/V2/V2/v2 [3]));
 XOR2_X2 \V3/V2/V2/V2/HA2/_1_  (.A(\V3/V2/V2/V2/w4 ),
    .B(\V3/V2/V2/V2/w3 ),
    .Z(\V3/V2/V2/v2 [2]));
 AND2_X1 \V3/V2/V2/V2/_0_  (.A1(A[14]),
    .A2(B[16]),
    .ZN(\V3/V2/V2/v2 [0]));
 AND2_X1 \V3/V2/V2/V2/_1_  (.A1(A[14]),
    .A2(B[17]),
    .ZN(\V3/V2/V2/V2/w1 ));
 AND2_X1 \V3/V2/V2/V2/_2_  (.A1(B[16]),
    .A2(A[15]),
    .ZN(\V3/V2/V2/V2/w2 ));
 AND2_X1 \V3/V2/V2/V2/_3_  (.A1(B[17]),
    .A2(A[15]),
    .ZN(\V3/V2/V2/V2/w3 ));
 AND2_X1 \V3/V2/V2/V3/HA1/_0_  (.A1(\V3/V2/V2/V3/w2 ),
    .A2(\V3/V2/V2/V3/w1 ),
    .ZN(\V3/V2/V2/V3/w4 ));
 XOR2_X2 \V3/V2/V2/V3/HA1/_1_  (.A(\V3/V2/V2/V3/w2 ),
    .B(\V3/V2/V2/V3/w1 ),
    .Z(\V3/V2/V2/v3 [1]));
 AND2_X1 \V3/V2/V2/V3/HA2/_0_  (.A1(\V3/V2/V2/V3/w4 ),
    .A2(\V3/V2/V2/V3/w3 ),
    .ZN(\V3/V2/V2/v3 [3]));
 XOR2_X2 \V3/V2/V2/V3/HA2/_1_  (.A(\V3/V2/V2/V3/w4 ),
    .B(\V3/V2/V2/V3/w3 ),
    .Z(\V3/V2/V2/v3 [2]));
 AND2_X1 \V3/V2/V2/V3/_0_  (.A1(A[12]),
    .A2(B[18]),
    .ZN(\V3/V2/V2/v3 [0]));
 AND2_X1 \V3/V2/V2/V3/_1_  (.A1(A[12]),
    .A2(B[19]),
    .ZN(\V3/V2/V2/V3/w1 ));
 AND2_X1 \V3/V2/V2/V3/_2_  (.A1(B[18]),
    .A2(A[13]),
    .ZN(\V3/V2/V2/V3/w2 ));
 AND2_X1 \V3/V2/V2/V3/_3_  (.A1(B[19]),
    .A2(A[13]),
    .ZN(\V3/V2/V2/V3/w3 ));
 AND2_X1 \V3/V2/V2/V4/HA1/_0_  (.A1(\V3/V2/V2/V4/w2 ),
    .A2(\V3/V2/V2/V4/w1 ),
    .ZN(\V3/V2/V2/V4/w4 ));
 XOR2_X2 \V3/V2/V2/V4/HA1/_1_  (.A(\V3/V2/V2/V4/w2 ),
    .B(\V3/V2/V2/V4/w1 ),
    .Z(\V3/V2/V2/v4 [1]));
 AND2_X1 \V3/V2/V2/V4/HA2/_0_  (.A1(\V3/V2/V2/V4/w4 ),
    .A2(\V3/V2/V2/V4/w3 ),
    .ZN(\V3/V2/V2/v4 [3]));
 XOR2_X2 \V3/V2/V2/V4/HA2/_1_  (.A(\V3/V2/V2/V4/w4 ),
    .B(\V3/V2/V2/V4/w3 ),
    .Z(\V3/V2/V2/v4 [2]));
 AND2_X1 \V3/V2/V2/V4/_0_  (.A1(A[14]),
    .A2(B[18]),
    .ZN(\V3/V2/V2/v4 [0]));
 AND2_X1 \V3/V2/V2/V4/_1_  (.A1(A[14]),
    .A2(B[19]),
    .ZN(\V3/V2/V2/V4/w1 ));
 AND2_X1 \V3/V2/V2/V4/_2_  (.A1(B[18]),
    .A2(A[15]),
    .ZN(\V3/V2/V2/V4/w2 ));
 AND2_X1 \V3/V2/V2/V4/_3_  (.A1(B[19]),
    .A2(A[15]),
    .ZN(\V3/V2/V2/V4/w3 ));
 OR2_X1 \V3/V2/V2/_0_  (.A1(\V3/V2/V2/c1 ),
    .A2(\V3/V2/V2/c2 ),
    .ZN(\V3/V2/V2/c3 ));
 AND2_X1 \V3/V2/V3/A1/M1/M1/_0_  (.A1(\V3/V2/V3/v2 [0]),
    .A2(\V3/V2/V3/v3 [0]),
    .ZN(\V3/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M1/M1/_1_  (.A(\V3/V2/V3/v2 [0]),
    .B(\V3/V2/V3/v3 [0]),
    .Z(\V3/V2/V3/A1/M1/s1 ));
 AND2_X1 \V3/V2/V3/A1/M1/M2/_0_  (.A1(\V3/V2/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M1/M2/_1_  (.A(\V3/V2/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/V3/s1 [0]));
 OR2_X1 \V3/V2/V3/A1/M1/_0_  (.A1(\V3/V2/V3/A1/M1/c1 ),
    .A2(\V3/V2/V3/A1/M1/c2 ),
    .ZN(\V3/V2/V3/A1/c1 ));
 AND2_X1 \V3/V2/V3/A1/M2/M1/_0_  (.A1(\V3/V2/V3/v2 [1]),
    .A2(\V3/V2/V3/v3 [1]),
    .ZN(\V3/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M2/M1/_1_  (.A(\V3/V2/V3/v2 [1]),
    .B(\V3/V2/V3/v3 [1]),
    .Z(\V3/V2/V3/A1/M2/s1 ));
 AND2_X1 \V3/V2/V3/A1/M2/M2/_0_  (.A1(\V3/V2/V3/A1/M2/s1 ),
    .A2(\V3/V2/V3/A1/c1 ),
    .ZN(\V3/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M2/M2/_1_  (.A(\V3/V2/V3/A1/M2/s1 ),
    .B(\V3/V2/V3/A1/c1 ),
    .Z(\V3/V2/V3/s1 [1]));
 OR2_X1 \V3/V2/V3/A1/M2/_0_  (.A1(\V3/V2/V3/A1/M2/c1 ),
    .A2(\V3/V2/V3/A1/M2/c2 ),
    .ZN(\V3/V2/V3/A1/c2 ));
 AND2_X1 \V3/V2/V3/A1/M3/M1/_0_  (.A1(\V3/V2/V3/v2 [2]),
    .A2(\V3/V2/V3/v3 [2]),
    .ZN(\V3/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M3/M1/_1_  (.A(\V3/V2/V3/v2 [2]),
    .B(\V3/V2/V3/v3 [2]),
    .Z(\V3/V2/V3/A1/M3/s1 ));
 AND2_X1 \V3/V2/V3/A1/M3/M2/_0_  (.A1(\V3/V2/V3/A1/M3/s1 ),
    .A2(\V3/V2/V3/A1/c2 ),
    .ZN(\V3/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M3/M2/_1_  (.A(\V3/V2/V3/A1/M3/s1 ),
    .B(\V3/V2/V3/A1/c2 ),
    .Z(\V3/V2/V3/s1 [2]));
 OR2_X1 \V3/V2/V3/A1/M3/_0_  (.A1(\V3/V2/V3/A1/M3/c1 ),
    .A2(\V3/V2/V3/A1/M3/c2 ),
    .ZN(\V3/V2/V3/A1/c3 ));
 AND2_X1 \V3/V2/V3/A1/M4/M1/_0_  (.A1(\V3/V2/V3/v2 [3]),
    .A2(\V3/V2/V3/v3 [3]),
    .ZN(\V3/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M4/M1/_1_  (.A(\V3/V2/V3/v2 [3]),
    .B(\V3/V2/V3/v3 [3]),
    .Z(\V3/V2/V3/A1/M4/s1 ));
 AND2_X1 \V3/V2/V3/A1/M4/M2/_0_  (.A1(\V3/V2/V3/A1/M4/s1 ),
    .A2(\V3/V2/V3/A1/c3 ),
    .ZN(\V3/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M4/M2/_1_  (.A(\V3/V2/V3/A1/M4/s1 ),
    .B(\V3/V2/V3/A1/c3 ),
    .Z(\V3/V2/V3/s1 [3]));
 OR2_X1 \V3/V2/V3/A1/M4/_0_  (.A1(\V3/V2/V3/A1/M4/c1 ),
    .A2(\V3/V2/V3/A1/M4/c2 ),
    .ZN(\V3/V2/V3/c1 ));
 AND2_X1 \V3/V2/V3/A2/M1/M1/_0_  (.A1(\V3/V2/V3/s1 [0]),
    .A2(\V3/V2/V3/v1 [2]),
    .ZN(\V3/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M1/M1/_1_  (.A(\V3/V2/V3/s1 [0]),
    .B(\V3/V2/V3/v1 [2]),
    .Z(\V3/V2/V3/A2/M1/s1 ));
 AND2_X1 \V3/V2/V3/A2/M1/M2/_0_  (.A1(\V3/V2/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M1/M2/_1_  (.A(\V3/V2/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v3 [2]));
 OR2_X1 \V3/V2/V3/A2/M1/_0_  (.A1(\V3/V2/V3/A2/M1/c1 ),
    .A2(\V3/V2/V3/A2/M1/c2 ),
    .ZN(\V3/V2/V3/A2/c1 ));
 AND2_X1 \V3/V2/V3/A2/M2/M1/_0_  (.A1(\V3/V2/V3/s1 [1]),
    .A2(\V3/V2/V3/v1 [3]),
    .ZN(\V3/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M2/M1/_1_  (.A(\V3/V2/V3/s1 [1]),
    .B(\V3/V2/V3/v1 [3]),
    .Z(\V3/V2/V3/A2/M2/s1 ));
 AND2_X1 \V3/V2/V3/A2/M2/M2/_0_  (.A1(\V3/V2/V3/A2/M2/s1 ),
    .A2(\V3/V2/V3/A2/c1 ),
    .ZN(\V3/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M2/M2/_1_  (.A(\V3/V2/V3/A2/M2/s1 ),
    .B(\V3/V2/V3/A2/c1 ),
    .Z(\V3/V2/v3 [3]));
 OR2_X1 \V3/V2/V3/A2/M2/_0_  (.A1(\V3/V2/V3/A2/M2/c1 ),
    .A2(\V3/V2/V3/A2/M2/c2 ),
    .ZN(\V3/V2/V3/A2/c2 ));
 AND2_X1 \V3/V2/V3/A2/M3/M1/_0_  (.A1(\V3/V2/V3/s1 [2]),
    .A2(ground),
    .ZN(\V3/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M3/M1/_1_  (.A(\V3/V2/V3/s1 [2]),
    .B(ground),
    .Z(\V3/V2/V3/A2/M3/s1 ));
 AND2_X1 \V3/V2/V3/A2/M3/M2/_0_  (.A1(\V3/V2/V3/A2/M3/s1 ),
    .A2(\V3/V2/V3/A2/c2 ),
    .ZN(\V3/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M3/M2/_1_  (.A(\V3/V2/V3/A2/M3/s1 ),
    .B(\V3/V2/V3/A2/c2 ),
    .Z(\V3/V2/V3/s2 [2]));
 OR2_X1 \V3/V2/V3/A2/M3/_0_  (.A1(\V3/V2/V3/A2/M3/c1 ),
    .A2(\V3/V2/V3/A2/M3/c2 ),
    .ZN(\V3/V2/V3/A2/c3 ));
 AND2_X1 \V3/V2/V3/A2/M4/M1/_0_  (.A1(\V3/V2/V3/s1 [3]),
    .A2(ground),
    .ZN(\V3/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M4/M1/_1_  (.A(\V3/V2/V3/s1 [3]),
    .B(ground),
    .Z(\V3/V2/V3/A2/M4/s1 ));
 AND2_X1 \V3/V2/V3/A2/M4/M2/_0_  (.A1(\V3/V2/V3/A2/M4/s1 ),
    .A2(\V3/V2/V3/A2/c3 ),
    .ZN(\V3/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M4/M2/_1_  (.A(\V3/V2/V3/A2/M4/s1 ),
    .B(\V3/V2/V3/A2/c3 ),
    .Z(\V3/V2/V3/s2 [3]));
 OR2_X1 \V3/V2/V3/A2/M4/_0_  (.A1(\V3/V2/V3/A2/M4/c1 ),
    .A2(\V3/V2/V3/A2/M4/c2 ),
    .ZN(\V3/V2/V3/c2 ));
 AND2_X1 \V3/V2/V3/A3/M1/M1/_0_  (.A1(\V3/V2/V3/v4 [0]),
    .A2(\V3/V2/V3/s2 [2]),
    .ZN(\V3/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M1/M1/_1_  (.A(\V3/V2/V3/v4 [0]),
    .B(\V3/V2/V3/s2 [2]),
    .Z(\V3/V2/V3/A3/M1/s1 ));
 AND2_X1 \V3/V2/V3/A3/M1/M2/_0_  (.A1(\V3/V2/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M1/M2/_1_  (.A(\V3/V2/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v3 [4]));
 OR2_X1 \V3/V2/V3/A3/M1/_0_  (.A1(\V3/V2/V3/A3/M1/c1 ),
    .A2(\V3/V2/V3/A3/M1/c2 ),
    .ZN(\V3/V2/V3/A3/c1 ));
 AND2_X1 \V3/V2/V3/A3/M2/M1/_0_  (.A1(\V3/V2/V3/v4 [1]),
    .A2(\V3/V2/V3/s2 [3]),
    .ZN(\V3/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M2/M1/_1_  (.A(\V3/V2/V3/v4 [1]),
    .B(\V3/V2/V3/s2 [3]),
    .Z(\V3/V2/V3/A3/M2/s1 ));
 AND2_X1 \V3/V2/V3/A3/M2/M2/_0_  (.A1(\V3/V2/V3/A3/M2/s1 ),
    .A2(\V3/V2/V3/A3/c1 ),
    .ZN(\V3/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M2/M2/_1_  (.A(\V3/V2/V3/A3/M2/s1 ),
    .B(\V3/V2/V3/A3/c1 ),
    .Z(\V3/V2/v3 [5]));
 OR2_X1 \V3/V2/V3/A3/M2/_0_  (.A1(\V3/V2/V3/A3/M2/c1 ),
    .A2(\V3/V2/V3/A3/M2/c2 ),
    .ZN(\V3/V2/V3/A3/c2 ));
 AND2_X1 \V3/V2/V3/A3/M3/M1/_0_  (.A1(\V3/V2/V3/v4 [2]),
    .A2(\V3/V2/V3/c3 ),
    .ZN(\V3/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M3/M1/_1_  (.A(\V3/V2/V3/v4 [2]),
    .B(\V3/V2/V3/c3 ),
    .Z(\V3/V2/V3/A3/M3/s1 ));
 AND2_X1 \V3/V2/V3/A3/M3/M2/_0_  (.A1(\V3/V2/V3/A3/M3/s1 ),
    .A2(\V3/V2/V3/A3/c2 ),
    .ZN(\V3/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M3/M2/_1_  (.A(\V3/V2/V3/A3/M3/s1 ),
    .B(\V3/V2/V3/A3/c2 ),
    .Z(\V3/V2/v3 [6]));
 OR2_X1 \V3/V2/V3/A3/M3/_0_  (.A1(\V3/V2/V3/A3/M3/c1 ),
    .A2(\V3/V2/V3/A3/M3/c2 ),
    .ZN(\V3/V2/V3/A3/c3 ));
 AND2_X1 \V3/V2/V3/A3/M4/M1/_0_  (.A1(\V3/V2/V3/v4 [3]),
    .A2(ground),
    .ZN(\V3/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M4/M1/_1_  (.A(\V3/V2/V3/v4 [3]),
    .B(ground),
    .Z(\V3/V2/V3/A3/M4/s1 ));
 AND2_X1 \V3/V2/V3/A3/M4/M2/_0_  (.A1(\V3/V2/V3/A3/M4/s1 ),
    .A2(\V3/V2/V3/A3/c3 ),
    .ZN(\V3/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M4/M2/_1_  (.A(\V3/V2/V3/A3/M4/s1 ),
    .B(\V3/V2/V3/A3/c3 ),
    .Z(\V3/V2/v3 [7]));
 OR2_X1 \V3/V2/V3/A3/M4/_0_  (.A1(\V3/V2/V3/A3/M4/c1 ),
    .A2(\V3/V2/V3/A3/M4/c2 ),
    .ZN(\V3/V2/V3/overflow ));
 AND2_X1 \V3/V2/V3/V1/HA1/_0_  (.A1(\V3/V2/V3/V1/w2 ),
    .A2(\V3/V2/V3/V1/w1 ),
    .ZN(\V3/V2/V3/V1/w4 ));
 XOR2_X2 \V3/V2/V3/V1/HA1/_1_  (.A(\V3/V2/V3/V1/w2 ),
    .B(\V3/V2/V3/V1/w1 ),
    .Z(\V3/V2/v3 [1]));
 AND2_X1 \V3/V2/V3/V1/HA2/_0_  (.A1(\V3/V2/V3/V1/w4 ),
    .A2(\V3/V2/V3/V1/w3 ),
    .ZN(\V3/V2/V3/v1 [3]));
 XOR2_X2 \V3/V2/V3/V1/HA2/_1_  (.A(\V3/V2/V3/V1/w4 ),
    .B(\V3/V2/V3/V1/w3 ),
    .Z(\V3/V2/V3/v1 [2]));
 AND2_X1 \V3/V2/V3/V1/_0_  (.A1(A[8]),
    .A2(B[20]),
    .ZN(\V3/V2/v3 [0]));
 AND2_X1 \V3/V2/V3/V1/_1_  (.A1(A[8]),
    .A2(B[21]),
    .ZN(\V3/V2/V3/V1/w1 ));
 AND2_X1 \V3/V2/V3/V1/_2_  (.A1(B[20]),
    .A2(A[9]),
    .ZN(\V3/V2/V3/V1/w2 ));
 AND2_X1 \V3/V2/V3/V1/_3_  (.A1(B[21]),
    .A2(A[9]),
    .ZN(\V3/V2/V3/V1/w3 ));
 AND2_X1 \V3/V2/V3/V2/HA1/_0_  (.A1(\V3/V2/V3/V2/w2 ),
    .A2(\V3/V2/V3/V2/w1 ),
    .ZN(\V3/V2/V3/V2/w4 ));
 XOR2_X2 \V3/V2/V3/V2/HA1/_1_  (.A(\V3/V2/V3/V2/w2 ),
    .B(\V3/V2/V3/V2/w1 ),
    .Z(\V3/V2/V3/v2 [1]));
 AND2_X1 \V3/V2/V3/V2/HA2/_0_  (.A1(\V3/V2/V3/V2/w4 ),
    .A2(\V3/V2/V3/V2/w3 ),
    .ZN(\V3/V2/V3/v2 [3]));
 XOR2_X2 \V3/V2/V3/V2/HA2/_1_  (.A(\V3/V2/V3/V2/w4 ),
    .B(\V3/V2/V3/V2/w3 ),
    .Z(\V3/V2/V3/v2 [2]));
 AND2_X1 \V3/V2/V3/V2/_0_  (.A1(A[10]),
    .A2(B[20]),
    .ZN(\V3/V2/V3/v2 [0]));
 AND2_X1 \V3/V2/V3/V2/_1_  (.A1(A[10]),
    .A2(B[21]),
    .ZN(\V3/V2/V3/V2/w1 ));
 AND2_X1 \V3/V2/V3/V2/_2_  (.A1(B[20]),
    .A2(A[11]),
    .ZN(\V3/V2/V3/V2/w2 ));
 AND2_X1 \V3/V2/V3/V2/_3_  (.A1(B[21]),
    .A2(A[11]),
    .ZN(\V3/V2/V3/V2/w3 ));
 AND2_X1 \V3/V2/V3/V3/HA1/_0_  (.A1(\V3/V2/V3/V3/w2 ),
    .A2(\V3/V2/V3/V3/w1 ),
    .ZN(\V3/V2/V3/V3/w4 ));
 XOR2_X2 \V3/V2/V3/V3/HA1/_1_  (.A(\V3/V2/V3/V3/w2 ),
    .B(\V3/V2/V3/V3/w1 ),
    .Z(\V3/V2/V3/v3 [1]));
 AND2_X1 \V3/V2/V3/V3/HA2/_0_  (.A1(\V3/V2/V3/V3/w4 ),
    .A2(\V3/V2/V3/V3/w3 ),
    .ZN(\V3/V2/V3/v3 [3]));
 XOR2_X2 \V3/V2/V3/V3/HA2/_1_  (.A(\V3/V2/V3/V3/w4 ),
    .B(\V3/V2/V3/V3/w3 ),
    .Z(\V3/V2/V3/v3 [2]));
 AND2_X1 \V3/V2/V3/V3/_0_  (.A1(A[8]),
    .A2(B[22]),
    .ZN(\V3/V2/V3/v3 [0]));
 AND2_X1 \V3/V2/V3/V3/_1_  (.A1(A[8]),
    .A2(B[23]),
    .ZN(\V3/V2/V3/V3/w1 ));
 AND2_X1 \V3/V2/V3/V3/_2_  (.A1(B[22]),
    .A2(A[9]),
    .ZN(\V3/V2/V3/V3/w2 ));
 AND2_X1 \V3/V2/V3/V3/_3_  (.A1(B[23]),
    .A2(A[9]),
    .ZN(\V3/V2/V3/V3/w3 ));
 AND2_X1 \V3/V2/V3/V4/HA1/_0_  (.A1(\V3/V2/V3/V4/w2 ),
    .A2(\V3/V2/V3/V4/w1 ),
    .ZN(\V3/V2/V3/V4/w4 ));
 XOR2_X2 \V3/V2/V3/V4/HA1/_1_  (.A(\V3/V2/V3/V4/w2 ),
    .B(\V3/V2/V3/V4/w1 ),
    .Z(\V3/V2/V3/v4 [1]));
 AND2_X1 \V3/V2/V3/V4/HA2/_0_  (.A1(\V3/V2/V3/V4/w4 ),
    .A2(\V3/V2/V3/V4/w3 ),
    .ZN(\V3/V2/V3/v4 [3]));
 XOR2_X2 \V3/V2/V3/V4/HA2/_1_  (.A(\V3/V2/V3/V4/w4 ),
    .B(\V3/V2/V3/V4/w3 ),
    .Z(\V3/V2/V3/v4 [2]));
 AND2_X1 \V3/V2/V3/V4/_0_  (.A1(A[10]),
    .A2(B[22]),
    .ZN(\V3/V2/V3/v4 [0]));
 AND2_X1 \V3/V2/V3/V4/_1_  (.A1(A[10]),
    .A2(B[23]),
    .ZN(\V3/V2/V3/V4/w1 ));
 AND2_X1 \V3/V2/V3/V4/_2_  (.A1(B[22]),
    .A2(A[11]),
    .ZN(\V3/V2/V3/V4/w2 ));
 AND2_X1 \V3/V2/V3/V4/_3_  (.A1(B[23]),
    .A2(A[11]),
    .ZN(\V3/V2/V3/V4/w3 ));
 OR2_X1 \V3/V2/V3/_0_  (.A1(\V3/V2/V3/c1 ),
    .A2(\V3/V2/V3/c2 ),
    .ZN(\V3/V2/V3/c3 ));
 AND2_X1 \V3/V2/V4/A1/M1/M1/_0_  (.A1(\V3/V2/V4/v2 [0]),
    .A2(\V3/V2/V4/v3 [0]),
    .ZN(\V3/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M1/M1/_1_  (.A(\V3/V2/V4/v2 [0]),
    .B(\V3/V2/V4/v3 [0]),
    .Z(\V3/V2/V4/A1/M1/s1 ));
 AND2_X1 \V3/V2/V4/A1/M1/M2/_0_  (.A1(\V3/V2/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M1/M2/_1_  (.A(\V3/V2/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/V4/s1 [0]));
 OR2_X1 \V3/V2/V4/A1/M1/_0_  (.A1(\V3/V2/V4/A1/M1/c1 ),
    .A2(\V3/V2/V4/A1/M1/c2 ),
    .ZN(\V3/V2/V4/A1/c1 ));
 AND2_X1 \V3/V2/V4/A1/M2/M1/_0_  (.A1(\V3/V2/V4/v2 [1]),
    .A2(\V3/V2/V4/v3 [1]),
    .ZN(\V3/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M2/M1/_1_  (.A(\V3/V2/V4/v2 [1]),
    .B(\V3/V2/V4/v3 [1]),
    .Z(\V3/V2/V4/A1/M2/s1 ));
 AND2_X1 \V3/V2/V4/A1/M2/M2/_0_  (.A1(\V3/V2/V4/A1/M2/s1 ),
    .A2(\V3/V2/V4/A1/c1 ),
    .ZN(\V3/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M2/M2/_1_  (.A(\V3/V2/V4/A1/M2/s1 ),
    .B(\V3/V2/V4/A1/c1 ),
    .Z(\V3/V2/V4/s1 [1]));
 OR2_X1 \V3/V2/V4/A1/M2/_0_  (.A1(\V3/V2/V4/A1/M2/c1 ),
    .A2(\V3/V2/V4/A1/M2/c2 ),
    .ZN(\V3/V2/V4/A1/c2 ));
 AND2_X1 \V3/V2/V4/A1/M3/M1/_0_  (.A1(\V3/V2/V4/v2 [2]),
    .A2(\V3/V2/V4/v3 [2]),
    .ZN(\V3/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M3/M1/_1_  (.A(\V3/V2/V4/v2 [2]),
    .B(\V3/V2/V4/v3 [2]),
    .Z(\V3/V2/V4/A1/M3/s1 ));
 AND2_X1 \V3/V2/V4/A1/M3/M2/_0_  (.A1(\V3/V2/V4/A1/M3/s1 ),
    .A2(\V3/V2/V4/A1/c2 ),
    .ZN(\V3/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M3/M2/_1_  (.A(\V3/V2/V4/A1/M3/s1 ),
    .B(\V3/V2/V4/A1/c2 ),
    .Z(\V3/V2/V4/s1 [2]));
 OR2_X1 \V3/V2/V4/A1/M3/_0_  (.A1(\V3/V2/V4/A1/M3/c1 ),
    .A2(\V3/V2/V4/A1/M3/c2 ),
    .ZN(\V3/V2/V4/A1/c3 ));
 AND2_X1 \V3/V2/V4/A1/M4/M1/_0_  (.A1(\V3/V2/V4/v2 [3]),
    .A2(\V3/V2/V4/v3 [3]),
    .ZN(\V3/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M4/M1/_1_  (.A(\V3/V2/V4/v2 [3]),
    .B(\V3/V2/V4/v3 [3]),
    .Z(\V3/V2/V4/A1/M4/s1 ));
 AND2_X1 \V3/V2/V4/A1/M4/M2/_0_  (.A1(\V3/V2/V4/A1/M4/s1 ),
    .A2(\V3/V2/V4/A1/c3 ),
    .ZN(\V3/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M4/M2/_1_  (.A(\V3/V2/V4/A1/M4/s1 ),
    .B(\V3/V2/V4/A1/c3 ),
    .Z(\V3/V2/V4/s1 [3]));
 OR2_X1 \V3/V2/V4/A1/M4/_0_  (.A1(\V3/V2/V4/A1/M4/c1 ),
    .A2(\V3/V2/V4/A1/M4/c2 ),
    .ZN(\V3/V2/V4/c1 ));
 AND2_X1 \V3/V2/V4/A2/M1/M1/_0_  (.A1(\V3/V2/V4/s1 [0]),
    .A2(\V3/V2/V4/v1 [2]),
    .ZN(\V3/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M1/M1/_1_  (.A(\V3/V2/V4/s1 [0]),
    .B(\V3/V2/V4/v1 [2]),
    .Z(\V3/V2/V4/A2/M1/s1 ));
 AND2_X1 \V3/V2/V4/A2/M1/M2/_0_  (.A1(\V3/V2/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M1/M2/_1_  (.A(\V3/V2/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v4 [2]));
 OR2_X1 \V3/V2/V4/A2/M1/_0_  (.A1(\V3/V2/V4/A2/M1/c1 ),
    .A2(\V3/V2/V4/A2/M1/c2 ),
    .ZN(\V3/V2/V4/A2/c1 ));
 AND2_X1 \V3/V2/V4/A2/M2/M1/_0_  (.A1(\V3/V2/V4/s1 [1]),
    .A2(\V3/V2/V4/v1 [3]),
    .ZN(\V3/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M2/M1/_1_  (.A(\V3/V2/V4/s1 [1]),
    .B(\V3/V2/V4/v1 [3]),
    .Z(\V3/V2/V4/A2/M2/s1 ));
 AND2_X1 \V3/V2/V4/A2/M2/M2/_0_  (.A1(\V3/V2/V4/A2/M2/s1 ),
    .A2(\V3/V2/V4/A2/c1 ),
    .ZN(\V3/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M2/M2/_1_  (.A(\V3/V2/V4/A2/M2/s1 ),
    .B(\V3/V2/V4/A2/c1 ),
    .Z(\V3/V2/v4 [3]));
 OR2_X1 \V3/V2/V4/A2/M2/_0_  (.A1(\V3/V2/V4/A2/M2/c1 ),
    .A2(\V3/V2/V4/A2/M2/c2 ),
    .ZN(\V3/V2/V4/A2/c2 ));
 AND2_X1 \V3/V2/V4/A2/M3/M1/_0_  (.A1(\V3/V2/V4/s1 [2]),
    .A2(ground),
    .ZN(\V3/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M3/M1/_1_  (.A(\V3/V2/V4/s1 [2]),
    .B(ground),
    .Z(\V3/V2/V4/A2/M3/s1 ));
 AND2_X1 \V3/V2/V4/A2/M3/M2/_0_  (.A1(\V3/V2/V4/A2/M3/s1 ),
    .A2(\V3/V2/V4/A2/c2 ),
    .ZN(\V3/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M3/M2/_1_  (.A(\V3/V2/V4/A2/M3/s1 ),
    .B(\V3/V2/V4/A2/c2 ),
    .Z(\V3/V2/V4/s2 [2]));
 OR2_X1 \V3/V2/V4/A2/M3/_0_  (.A1(\V3/V2/V4/A2/M3/c1 ),
    .A2(\V3/V2/V4/A2/M3/c2 ),
    .ZN(\V3/V2/V4/A2/c3 ));
 AND2_X1 \V3/V2/V4/A2/M4/M1/_0_  (.A1(\V3/V2/V4/s1 [3]),
    .A2(ground),
    .ZN(\V3/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M4/M1/_1_  (.A(\V3/V2/V4/s1 [3]),
    .B(ground),
    .Z(\V3/V2/V4/A2/M4/s1 ));
 AND2_X1 \V3/V2/V4/A2/M4/M2/_0_  (.A1(\V3/V2/V4/A2/M4/s1 ),
    .A2(\V3/V2/V4/A2/c3 ),
    .ZN(\V3/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M4/M2/_1_  (.A(\V3/V2/V4/A2/M4/s1 ),
    .B(\V3/V2/V4/A2/c3 ),
    .Z(\V3/V2/V4/s2 [3]));
 OR2_X1 \V3/V2/V4/A2/M4/_0_  (.A1(\V3/V2/V4/A2/M4/c1 ),
    .A2(\V3/V2/V4/A2/M4/c2 ),
    .ZN(\V3/V2/V4/c2 ));
 AND2_X1 \V3/V2/V4/A3/M1/M1/_0_  (.A1(\V3/V2/V4/v4 [0]),
    .A2(\V3/V2/V4/s2 [2]),
    .ZN(\V3/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M1/M1/_1_  (.A(\V3/V2/V4/v4 [0]),
    .B(\V3/V2/V4/s2 [2]),
    .Z(\V3/V2/V4/A3/M1/s1 ));
 AND2_X1 \V3/V2/V4/A3/M1/M2/_0_  (.A1(\V3/V2/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M1/M2/_1_  (.A(\V3/V2/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V2/v4 [4]));
 OR2_X1 \V3/V2/V4/A3/M1/_0_  (.A1(\V3/V2/V4/A3/M1/c1 ),
    .A2(\V3/V2/V4/A3/M1/c2 ),
    .ZN(\V3/V2/V4/A3/c1 ));
 AND2_X1 \V3/V2/V4/A3/M2/M1/_0_  (.A1(\V3/V2/V4/v4 [1]),
    .A2(\V3/V2/V4/s2 [3]),
    .ZN(\V3/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M2/M1/_1_  (.A(\V3/V2/V4/v4 [1]),
    .B(\V3/V2/V4/s2 [3]),
    .Z(\V3/V2/V4/A3/M2/s1 ));
 AND2_X1 \V3/V2/V4/A3/M2/M2/_0_  (.A1(\V3/V2/V4/A3/M2/s1 ),
    .A2(\V3/V2/V4/A3/c1 ),
    .ZN(\V3/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M2/M2/_1_  (.A(\V3/V2/V4/A3/M2/s1 ),
    .B(\V3/V2/V4/A3/c1 ),
    .Z(\V3/V2/v4 [5]));
 OR2_X1 \V3/V2/V4/A3/M2/_0_  (.A1(\V3/V2/V4/A3/M2/c1 ),
    .A2(\V3/V2/V4/A3/M2/c2 ),
    .ZN(\V3/V2/V4/A3/c2 ));
 AND2_X1 \V3/V2/V4/A3/M3/M1/_0_  (.A1(\V3/V2/V4/v4 [2]),
    .A2(\V3/V2/V4/c3 ),
    .ZN(\V3/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M3/M1/_1_  (.A(\V3/V2/V4/v4 [2]),
    .B(\V3/V2/V4/c3 ),
    .Z(\V3/V2/V4/A3/M3/s1 ));
 AND2_X1 \V3/V2/V4/A3/M3/M2/_0_  (.A1(\V3/V2/V4/A3/M3/s1 ),
    .A2(\V3/V2/V4/A3/c2 ),
    .ZN(\V3/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M3/M2/_1_  (.A(\V3/V2/V4/A3/M3/s1 ),
    .B(\V3/V2/V4/A3/c2 ),
    .Z(\V3/V2/v4 [6]));
 OR2_X1 \V3/V2/V4/A3/M3/_0_  (.A1(\V3/V2/V4/A3/M3/c1 ),
    .A2(\V3/V2/V4/A3/M3/c2 ),
    .ZN(\V3/V2/V4/A3/c3 ));
 AND2_X1 \V3/V2/V4/A3/M4/M1/_0_  (.A1(\V3/V2/V4/v4 [3]),
    .A2(ground),
    .ZN(\V3/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M4/M1/_1_  (.A(\V3/V2/V4/v4 [3]),
    .B(ground),
    .Z(\V3/V2/V4/A3/M4/s1 ));
 AND2_X1 \V3/V2/V4/A3/M4/M2/_0_  (.A1(\V3/V2/V4/A3/M4/s1 ),
    .A2(\V3/V2/V4/A3/c3 ),
    .ZN(\V3/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M4/M2/_1_  (.A(\V3/V2/V4/A3/M4/s1 ),
    .B(\V3/V2/V4/A3/c3 ),
    .Z(\V3/V2/v4 [7]));
 OR2_X1 \V3/V2/V4/A3/M4/_0_  (.A1(\V3/V2/V4/A3/M4/c1 ),
    .A2(\V3/V2/V4/A3/M4/c2 ),
    .ZN(\V3/V2/V4/overflow ));
 AND2_X1 \V3/V2/V4/V1/HA1/_0_  (.A1(\V3/V2/V4/V1/w2 ),
    .A2(\V3/V2/V4/V1/w1 ),
    .ZN(\V3/V2/V4/V1/w4 ));
 XOR2_X2 \V3/V2/V4/V1/HA1/_1_  (.A(\V3/V2/V4/V1/w2 ),
    .B(\V3/V2/V4/V1/w1 ),
    .Z(\V3/V2/v4 [1]));
 AND2_X1 \V3/V2/V4/V1/HA2/_0_  (.A1(\V3/V2/V4/V1/w4 ),
    .A2(\V3/V2/V4/V1/w3 ),
    .ZN(\V3/V2/V4/v1 [3]));
 XOR2_X2 \V3/V2/V4/V1/HA2/_1_  (.A(\V3/V2/V4/V1/w4 ),
    .B(\V3/V2/V4/V1/w3 ),
    .Z(\V3/V2/V4/v1 [2]));
 AND2_X1 \V3/V2/V4/V1/_0_  (.A1(A[12]),
    .A2(B[20]),
    .ZN(\V3/V2/v4 [0]));
 AND2_X1 \V3/V2/V4/V1/_1_  (.A1(A[12]),
    .A2(B[21]),
    .ZN(\V3/V2/V4/V1/w1 ));
 AND2_X1 \V3/V2/V4/V1/_2_  (.A1(B[20]),
    .A2(A[13]),
    .ZN(\V3/V2/V4/V1/w2 ));
 AND2_X1 \V3/V2/V4/V1/_3_  (.A1(B[21]),
    .A2(A[13]),
    .ZN(\V3/V2/V4/V1/w3 ));
 AND2_X1 \V3/V2/V4/V2/HA1/_0_  (.A1(\V3/V2/V4/V2/w2 ),
    .A2(\V3/V2/V4/V2/w1 ),
    .ZN(\V3/V2/V4/V2/w4 ));
 XOR2_X2 \V3/V2/V4/V2/HA1/_1_  (.A(\V3/V2/V4/V2/w2 ),
    .B(\V3/V2/V4/V2/w1 ),
    .Z(\V3/V2/V4/v2 [1]));
 AND2_X1 \V3/V2/V4/V2/HA2/_0_  (.A1(\V3/V2/V4/V2/w4 ),
    .A2(\V3/V2/V4/V2/w3 ),
    .ZN(\V3/V2/V4/v2 [3]));
 XOR2_X2 \V3/V2/V4/V2/HA2/_1_  (.A(\V3/V2/V4/V2/w4 ),
    .B(\V3/V2/V4/V2/w3 ),
    .Z(\V3/V2/V4/v2 [2]));
 AND2_X1 \V3/V2/V4/V2/_0_  (.A1(A[14]),
    .A2(B[20]),
    .ZN(\V3/V2/V4/v2 [0]));
 AND2_X1 \V3/V2/V4/V2/_1_  (.A1(A[14]),
    .A2(B[21]),
    .ZN(\V3/V2/V4/V2/w1 ));
 AND2_X1 \V3/V2/V4/V2/_2_  (.A1(B[20]),
    .A2(A[15]),
    .ZN(\V3/V2/V4/V2/w2 ));
 AND2_X1 \V3/V2/V4/V2/_3_  (.A1(B[21]),
    .A2(A[15]),
    .ZN(\V3/V2/V4/V2/w3 ));
 AND2_X1 \V3/V2/V4/V3/HA1/_0_  (.A1(\V3/V2/V4/V3/w2 ),
    .A2(\V3/V2/V4/V3/w1 ),
    .ZN(\V3/V2/V4/V3/w4 ));
 XOR2_X2 \V3/V2/V4/V3/HA1/_1_  (.A(\V3/V2/V4/V3/w2 ),
    .B(\V3/V2/V4/V3/w1 ),
    .Z(\V3/V2/V4/v3 [1]));
 AND2_X1 \V3/V2/V4/V3/HA2/_0_  (.A1(\V3/V2/V4/V3/w4 ),
    .A2(\V3/V2/V4/V3/w3 ),
    .ZN(\V3/V2/V4/v3 [3]));
 XOR2_X2 \V3/V2/V4/V3/HA2/_1_  (.A(\V3/V2/V4/V3/w4 ),
    .B(\V3/V2/V4/V3/w3 ),
    .Z(\V3/V2/V4/v3 [2]));
 AND2_X1 \V3/V2/V4/V3/_0_  (.A1(A[12]),
    .A2(B[22]),
    .ZN(\V3/V2/V4/v3 [0]));
 AND2_X1 \V3/V2/V4/V3/_1_  (.A1(A[12]),
    .A2(B[23]),
    .ZN(\V3/V2/V4/V3/w1 ));
 AND2_X1 \V3/V2/V4/V3/_2_  (.A1(B[22]),
    .A2(A[13]),
    .ZN(\V3/V2/V4/V3/w2 ));
 AND2_X1 \V3/V2/V4/V3/_3_  (.A1(B[23]),
    .A2(A[13]),
    .ZN(\V3/V2/V4/V3/w3 ));
 AND2_X1 \V3/V2/V4/V4/HA1/_0_  (.A1(\V3/V2/V4/V4/w2 ),
    .A2(\V3/V2/V4/V4/w1 ),
    .ZN(\V3/V2/V4/V4/w4 ));
 XOR2_X2 \V3/V2/V4/V4/HA1/_1_  (.A(\V3/V2/V4/V4/w2 ),
    .B(\V3/V2/V4/V4/w1 ),
    .Z(\V3/V2/V4/v4 [1]));
 AND2_X1 \V3/V2/V4/V4/HA2/_0_  (.A1(\V3/V2/V4/V4/w4 ),
    .A2(\V3/V2/V4/V4/w3 ),
    .ZN(\V3/V2/V4/v4 [3]));
 XOR2_X2 \V3/V2/V4/V4/HA2/_1_  (.A(\V3/V2/V4/V4/w4 ),
    .B(\V3/V2/V4/V4/w3 ),
    .Z(\V3/V2/V4/v4 [2]));
 AND2_X1 \V3/V2/V4/V4/_0_  (.A1(A[14]),
    .A2(B[22]),
    .ZN(\V3/V2/V4/v4 [0]));
 AND2_X1 \V3/V2/V4/V4/_1_  (.A1(A[14]),
    .A2(B[23]),
    .ZN(\V3/V2/V4/V4/w1 ));
 AND2_X1 \V3/V2/V4/V4/_2_  (.A1(B[22]),
    .A2(A[15]),
    .ZN(\V3/V2/V4/V4/w2 ));
 AND2_X1 \V3/V2/V4/V4/_3_  (.A1(B[23]),
    .A2(A[15]),
    .ZN(\V3/V2/V4/V4/w3 ));
 OR2_X1 \V3/V2/V4/_0_  (.A1(\V3/V2/V4/c1 ),
    .A2(\V3/V2/V4/c2 ),
    .ZN(\V3/V2/V4/c3 ));
 OR2_X1 \V3/V2/_0_  (.A1(\V3/V2/c1 ),
    .A2(\V3/V2/c2 ),
    .ZN(\V3/V2/c3 ));
 AND2_X1 \V3/V3/A1/A1/M1/M1/_0_  (.A1(\V3/V3/v2 [0]),
    .A2(\V3/V3/v3 [0]),
    .ZN(\V3/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M1/M1/_1_  (.A(\V3/V3/v2 [0]),
    .B(\V3/V3/v3 [0]),
    .Z(\V3/V3/A1/A1/M1/s1 ));
 AND2_X1 \V3/V3/A1/A1/M1/M2/_0_  (.A1(\V3/V3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M1/M2/_1_  (.A(\V3/V3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/s1 [0]));
 OR2_X1 \V3/V3/A1/A1/M1/_0_  (.A1(\V3/V3/A1/A1/M1/c1 ),
    .A2(\V3/V3/A1/A1/M1/c2 ),
    .ZN(\V3/V3/A1/A1/c1 ));
 AND2_X1 \V3/V3/A1/A1/M2/M1/_0_  (.A1(\V3/V3/v2 [1]),
    .A2(\V3/V3/v3 [1]),
    .ZN(\V3/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M2/M1/_1_  (.A(\V3/V3/v2 [1]),
    .B(\V3/V3/v3 [1]),
    .Z(\V3/V3/A1/A1/M2/s1 ));
 AND2_X1 \V3/V3/A1/A1/M2/M2/_0_  (.A1(\V3/V3/A1/A1/M2/s1 ),
    .A2(\V3/V3/A1/A1/c1 ),
    .ZN(\V3/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M2/M2/_1_  (.A(\V3/V3/A1/A1/M2/s1 ),
    .B(\V3/V3/A1/A1/c1 ),
    .Z(\V3/V3/s1 [1]));
 OR2_X1 \V3/V3/A1/A1/M2/_0_  (.A1(\V3/V3/A1/A1/M2/c1 ),
    .A2(\V3/V3/A1/A1/M2/c2 ),
    .ZN(\V3/V3/A1/A1/c2 ));
 AND2_X1 \V3/V3/A1/A1/M3/M1/_0_  (.A1(\V3/V3/v2 [2]),
    .A2(\V3/V3/v3 [2]),
    .ZN(\V3/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M3/M1/_1_  (.A(\V3/V3/v2 [2]),
    .B(\V3/V3/v3 [2]),
    .Z(\V3/V3/A1/A1/M3/s1 ));
 AND2_X1 \V3/V3/A1/A1/M3/M2/_0_  (.A1(\V3/V3/A1/A1/M3/s1 ),
    .A2(\V3/V3/A1/A1/c2 ),
    .ZN(\V3/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M3/M2/_1_  (.A(\V3/V3/A1/A1/M3/s1 ),
    .B(\V3/V3/A1/A1/c2 ),
    .Z(\V3/V3/s1 [2]));
 OR2_X1 \V3/V3/A1/A1/M3/_0_  (.A1(\V3/V3/A1/A1/M3/c1 ),
    .A2(\V3/V3/A1/A1/M3/c2 ),
    .ZN(\V3/V3/A1/A1/c3 ));
 AND2_X1 \V3/V3/A1/A1/M4/M1/_0_  (.A1(\V3/V3/v2 [3]),
    .A2(\V3/V3/v3 [3]),
    .ZN(\V3/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M4/M1/_1_  (.A(\V3/V3/v2 [3]),
    .B(\V3/V3/v3 [3]),
    .Z(\V3/V3/A1/A1/M4/s1 ));
 AND2_X1 \V3/V3/A1/A1/M4/M2/_0_  (.A1(\V3/V3/A1/A1/M4/s1 ),
    .A2(\V3/V3/A1/A1/c3 ),
    .ZN(\V3/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M4/M2/_1_  (.A(\V3/V3/A1/A1/M4/s1 ),
    .B(\V3/V3/A1/A1/c3 ),
    .Z(\V3/V3/s1 [3]));
 OR2_X1 \V3/V3/A1/A1/M4/_0_  (.A1(\V3/V3/A1/A1/M4/c1 ),
    .A2(\V3/V3/A1/A1/M4/c2 ),
    .ZN(\V3/V3/A1/c1 ));
 AND2_X1 \V3/V3/A1/A2/M1/M1/_0_  (.A1(\V3/V3/v2 [4]),
    .A2(\V3/V3/v3 [4]),
    .ZN(\V3/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M1/M1/_1_  (.A(\V3/V3/v2 [4]),
    .B(\V3/V3/v3 [4]),
    .Z(\V3/V3/A1/A2/M1/s1 ));
 AND2_X1 \V3/V3/A1/A2/M1/M2/_0_  (.A1(\V3/V3/A1/A2/M1/s1 ),
    .A2(\V3/V3/A1/c1 ),
    .ZN(\V3/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M1/M2/_1_  (.A(\V3/V3/A1/A2/M1/s1 ),
    .B(\V3/V3/A1/c1 ),
    .Z(\V3/V3/s1 [4]));
 OR2_X1 \V3/V3/A1/A2/M1/_0_  (.A1(\V3/V3/A1/A2/M1/c1 ),
    .A2(\V3/V3/A1/A2/M1/c2 ),
    .ZN(\V3/V3/A1/A2/c1 ));
 AND2_X1 \V3/V3/A1/A2/M2/M1/_0_  (.A1(\V3/V3/v2 [5]),
    .A2(\V3/V3/v3 [5]),
    .ZN(\V3/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M2/M1/_1_  (.A(\V3/V3/v2 [5]),
    .B(\V3/V3/v3 [5]),
    .Z(\V3/V3/A1/A2/M2/s1 ));
 AND2_X1 \V3/V3/A1/A2/M2/M2/_0_  (.A1(\V3/V3/A1/A2/M2/s1 ),
    .A2(\V3/V3/A1/A2/c1 ),
    .ZN(\V3/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M2/M2/_1_  (.A(\V3/V3/A1/A2/M2/s1 ),
    .B(\V3/V3/A1/A2/c1 ),
    .Z(\V3/V3/s1 [5]));
 OR2_X1 \V3/V3/A1/A2/M2/_0_  (.A1(\V3/V3/A1/A2/M2/c1 ),
    .A2(\V3/V3/A1/A2/M2/c2 ),
    .ZN(\V3/V3/A1/A2/c2 ));
 AND2_X1 \V3/V3/A1/A2/M3/M1/_0_  (.A1(\V3/V3/v2 [6]),
    .A2(\V3/V3/v3 [6]),
    .ZN(\V3/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M3/M1/_1_  (.A(\V3/V3/v2 [6]),
    .B(\V3/V3/v3 [6]),
    .Z(\V3/V3/A1/A2/M3/s1 ));
 AND2_X1 \V3/V3/A1/A2/M3/M2/_0_  (.A1(\V3/V3/A1/A2/M3/s1 ),
    .A2(\V3/V3/A1/A2/c2 ),
    .ZN(\V3/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M3/M2/_1_  (.A(\V3/V3/A1/A2/M3/s1 ),
    .B(\V3/V3/A1/A2/c2 ),
    .Z(\V3/V3/s1 [6]));
 OR2_X1 \V3/V3/A1/A2/M3/_0_  (.A1(\V3/V3/A1/A2/M3/c1 ),
    .A2(\V3/V3/A1/A2/M3/c2 ),
    .ZN(\V3/V3/A1/A2/c3 ));
 AND2_X1 \V3/V3/A1/A2/M4/M1/_0_  (.A1(\V3/V3/v2 [7]),
    .A2(\V3/V3/v3 [7]),
    .ZN(\V3/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M4/M1/_1_  (.A(\V3/V3/v2 [7]),
    .B(\V3/V3/v3 [7]),
    .Z(\V3/V3/A1/A2/M4/s1 ));
 AND2_X1 \V3/V3/A1/A2/M4/M2/_0_  (.A1(\V3/V3/A1/A2/M4/s1 ),
    .A2(\V3/V3/A1/A2/c3 ),
    .ZN(\V3/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M4/M2/_1_  (.A(\V3/V3/A1/A2/M4/s1 ),
    .B(\V3/V3/A1/A2/c3 ),
    .Z(\V3/V3/s1 [7]));
 OR2_X1 \V3/V3/A1/A2/M4/_0_  (.A1(\V3/V3/A1/A2/M4/c1 ),
    .A2(\V3/V3/A1/A2/M4/c2 ),
    .ZN(\V3/V3/c1 ));
 AND2_X1 \V3/V3/A2/A1/M1/M1/_0_  (.A1(\V3/V3/s1 [0]),
    .A2(\V3/V3/v1 [4]),
    .ZN(\V3/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M1/M1/_1_  (.A(\V3/V3/s1 [0]),
    .B(\V3/V3/v1 [4]),
    .Z(\V3/V3/A2/A1/M1/s1 ));
 AND2_X1 \V3/V3/A2/A1/M1/M2/_0_  (.A1(\V3/V3/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M1/M2/_1_  (.A(\V3/V3/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v3 [4]));
 OR2_X1 \V3/V3/A2/A1/M1/_0_  (.A1(\V3/V3/A2/A1/M1/c1 ),
    .A2(\V3/V3/A2/A1/M1/c2 ),
    .ZN(\V3/V3/A2/A1/c1 ));
 AND2_X1 \V3/V3/A2/A1/M2/M1/_0_  (.A1(\V3/V3/s1 [1]),
    .A2(\V3/V3/v1 [5]),
    .ZN(\V3/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M2/M1/_1_  (.A(\V3/V3/s1 [1]),
    .B(\V3/V3/v1 [5]),
    .Z(\V3/V3/A2/A1/M2/s1 ));
 AND2_X1 \V3/V3/A2/A1/M2/M2/_0_  (.A1(\V3/V3/A2/A1/M2/s1 ),
    .A2(\V3/V3/A2/A1/c1 ),
    .ZN(\V3/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M2/M2/_1_  (.A(\V3/V3/A2/A1/M2/s1 ),
    .B(\V3/V3/A2/A1/c1 ),
    .Z(\V3/v3 [5]));
 OR2_X1 \V3/V3/A2/A1/M2/_0_  (.A1(\V3/V3/A2/A1/M2/c1 ),
    .A2(\V3/V3/A2/A1/M2/c2 ),
    .ZN(\V3/V3/A2/A1/c2 ));
 AND2_X1 \V3/V3/A2/A1/M3/M1/_0_  (.A1(\V3/V3/s1 [2]),
    .A2(\V3/V3/v1 [6]),
    .ZN(\V3/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M3/M1/_1_  (.A(\V3/V3/s1 [2]),
    .B(\V3/V3/v1 [6]),
    .Z(\V3/V3/A2/A1/M3/s1 ));
 AND2_X1 \V3/V3/A2/A1/M3/M2/_0_  (.A1(\V3/V3/A2/A1/M3/s1 ),
    .A2(\V3/V3/A2/A1/c2 ),
    .ZN(\V3/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M3/M2/_1_  (.A(\V3/V3/A2/A1/M3/s1 ),
    .B(\V3/V3/A2/A1/c2 ),
    .Z(\V3/v3 [6]));
 OR2_X1 \V3/V3/A2/A1/M3/_0_  (.A1(\V3/V3/A2/A1/M3/c1 ),
    .A2(\V3/V3/A2/A1/M3/c2 ),
    .ZN(\V3/V3/A2/A1/c3 ));
 AND2_X1 \V3/V3/A2/A1/M4/M1/_0_  (.A1(\V3/V3/s1 [3]),
    .A2(\V3/V3/v1 [7]),
    .ZN(\V3/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M4/M1/_1_  (.A(\V3/V3/s1 [3]),
    .B(\V3/V3/v1 [7]),
    .Z(\V3/V3/A2/A1/M4/s1 ));
 AND2_X1 \V3/V3/A2/A1/M4/M2/_0_  (.A1(\V3/V3/A2/A1/M4/s1 ),
    .A2(\V3/V3/A2/A1/c3 ),
    .ZN(\V3/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M4/M2/_1_  (.A(\V3/V3/A2/A1/M4/s1 ),
    .B(\V3/V3/A2/A1/c3 ),
    .Z(\V3/v3 [7]));
 OR2_X1 \V3/V3/A2/A1/M4/_0_  (.A1(\V3/V3/A2/A1/M4/c1 ),
    .A2(\V3/V3/A2/A1/M4/c2 ),
    .ZN(\V3/V3/A2/c1 ));
 AND2_X1 \V3/V3/A2/A2/M1/M1/_0_  (.A1(\V3/V3/s1 [4]),
    .A2(ground),
    .ZN(\V3/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M1/M1/_1_  (.A(\V3/V3/s1 [4]),
    .B(ground),
    .Z(\V3/V3/A2/A2/M1/s1 ));
 AND2_X1 \V3/V3/A2/A2/M1/M2/_0_  (.A1(\V3/V3/A2/A2/M1/s1 ),
    .A2(\V3/V3/A2/c1 ),
    .ZN(\V3/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M1/M2/_1_  (.A(\V3/V3/A2/A2/M1/s1 ),
    .B(\V3/V3/A2/c1 ),
    .Z(\V3/V3/s2 [4]));
 OR2_X1 \V3/V3/A2/A2/M1/_0_  (.A1(\V3/V3/A2/A2/M1/c1 ),
    .A2(\V3/V3/A2/A2/M1/c2 ),
    .ZN(\V3/V3/A2/A2/c1 ));
 AND2_X1 \V3/V3/A2/A2/M2/M1/_0_  (.A1(\V3/V3/s1 [5]),
    .A2(ground),
    .ZN(\V3/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M2/M1/_1_  (.A(\V3/V3/s1 [5]),
    .B(ground),
    .Z(\V3/V3/A2/A2/M2/s1 ));
 AND2_X1 \V3/V3/A2/A2/M2/M2/_0_  (.A1(\V3/V3/A2/A2/M2/s1 ),
    .A2(\V3/V3/A2/A2/c1 ),
    .ZN(\V3/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M2/M2/_1_  (.A(\V3/V3/A2/A2/M2/s1 ),
    .B(\V3/V3/A2/A2/c1 ),
    .Z(\V3/V3/s2 [5]));
 OR2_X1 \V3/V3/A2/A2/M2/_0_  (.A1(\V3/V3/A2/A2/M2/c1 ),
    .A2(\V3/V3/A2/A2/M2/c2 ),
    .ZN(\V3/V3/A2/A2/c2 ));
 AND2_X1 \V3/V3/A2/A2/M3/M1/_0_  (.A1(\V3/V3/s1 [6]),
    .A2(ground),
    .ZN(\V3/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M3/M1/_1_  (.A(\V3/V3/s1 [6]),
    .B(ground),
    .Z(\V3/V3/A2/A2/M3/s1 ));
 AND2_X1 \V3/V3/A2/A2/M3/M2/_0_  (.A1(\V3/V3/A2/A2/M3/s1 ),
    .A2(\V3/V3/A2/A2/c2 ),
    .ZN(\V3/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M3/M2/_1_  (.A(\V3/V3/A2/A2/M3/s1 ),
    .B(\V3/V3/A2/A2/c2 ),
    .Z(\V3/V3/s2 [6]));
 OR2_X1 \V3/V3/A2/A2/M3/_0_  (.A1(\V3/V3/A2/A2/M3/c1 ),
    .A2(\V3/V3/A2/A2/M3/c2 ),
    .ZN(\V3/V3/A2/A2/c3 ));
 AND2_X1 \V3/V3/A2/A2/M4/M1/_0_  (.A1(\V3/V3/s1 [7]),
    .A2(ground),
    .ZN(\V3/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M4/M1/_1_  (.A(\V3/V3/s1 [7]),
    .B(ground),
    .Z(\V3/V3/A2/A2/M4/s1 ));
 AND2_X1 \V3/V3/A2/A2/M4/M2/_0_  (.A1(\V3/V3/A2/A2/M4/s1 ),
    .A2(\V3/V3/A2/A2/c3 ),
    .ZN(\V3/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M4/M2/_1_  (.A(\V3/V3/A2/A2/M4/s1 ),
    .B(\V3/V3/A2/A2/c3 ),
    .Z(\V3/V3/s2 [7]));
 OR2_X1 \V3/V3/A2/A2/M4/_0_  (.A1(\V3/V3/A2/A2/M4/c1 ),
    .A2(\V3/V3/A2/A2/M4/c2 ),
    .ZN(\V3/V3/c2 ));
 AND2_X1 \V3/V3/A3/A1/M1/M1/_0_  (.A1(\V3/V3/v4 [0]),
    .A2(\V3/V3/s2 [4]),
    .ZN(\V3/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M1/M1/_1_  (.A(\V3/V3/v4 [0]),
    .B(\V3/V3/s2 [4]),
    .Z(\V3/V3/A3/A1/M1/s1 ));
 AND2_X1 \V3/V3/A3/A1/M1/M2/_0_  (.A1(\V3/V3/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M1/M2/_1_  (.A(\V3/V3/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v3 [8]));
 OR2_X1 \V3/V3/A3/A1/M1/_0_  (.A1(\V3/V3/A3/A1/M1/c1 ),
    .A2(\V3/V3/A3/A1/M1/c2 ),
    .ZN(\V3/V3/A3/A1/c1 ));
 AND2_X1 \V3/V3/A3/A1/M2/M1/_0_  (.A1(\V3/V3/v4 [1]),
    .A2(\V3/V3/s2 [5]),
    .ZN(\V3/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M2/M1/_1_  (.A(\V3/V3/v4 [1]),
    .B(\V3/V3/s2 [5]),
    .Z(\V3/V3/A3/A1/M2/s1 ));
 AND2_X1 \V3/V3/A3/A1/M2/M2/_0_  (.A1(\V3/V3/A3/A1/M2/s1 ),
    .A2(\V3/V3/A3/A1/c1 ),
    .ZN(\V3/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M2/M2/_1_  (.A(\V3/V3/A3/A1/M2/s1 ),
    .B(\V3/V3/A3/A1/c1 ),
    .Z(\V3/v3 [9]));
 OR2_X1 \V3/V3/A3/A1/M2/_0_  (.A1(\V3/V3/A3/A1/M2/c1 ),
    .A2(\V3/V3/A3/A1/M2/c2 ),
    .ZN(\V3/V3/A3/A1/c2 ));
 AND2_X1 \V3/V3/A3/A1/M3/M1/_0_  (.A1(\V3/V3/v4 [2]),
    .A2(\V3/V3/s2 [6]),
    .ZN(\V3/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M3/M1/_1_  (.A(\V3/V3/v4 [2]),
    .B(\V3/V3/s2 [6]),
    .Z(\V3/V3/A3/A1/M3/s1 ));
 AND2_X1 \V3/V3/A3/A1/M3/M2/_0_  (.A1(\V3/V3/A3/A1/M3/s1 ),
    .A2(\V3/V3/A3/A1/c2 ),
    .ZN(\V3/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M3/M2/_1_  (.A(\V3/V3/A3/A1/M3/s1 ),
    .B(\V3/V3/A3/A1/c2 ),
    .Z(\V3/v3 [10]));
 OR2_X1 \V3/V3/A3/A1/M3/_0_  (.A1(\V3/V3/A3/A1/M3/c1 ),
    .A2(\V3/V3/A3/A1/M3/c2 ),
    .ZN(\V3/V3/A3/A1/c3 ));
 AND2_X1 \V3/V3/A3/A1/M4/M1/_0_  (.A1(\V3/V3/v4 [3]),
    .A2(\V3/V3/s2 [7]),
    .ZN(\V3/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M4/M1/_1_  (.A(\V3/V3/v4 [3]),
    .B(\V3/V3/s2 [7]),
    .Z(\V3/V3/A3/A1/M4/s1 ));
 AND2_X1 \V3/V3/A3/A1/M4/M2/_0_  (.A1(\V3/V3/A3/A1/M4/s1 ),
    .A2(\V3/V3/A3/A1/c3 ),
    .ZN(\V3/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M4/M2/_1_  (.A(\V3/V3/A3/A1/M4/s1 ),
    .B(\V3/V3/A3/A1/c3 ),
    .Z(\V3/v3 [11]));
 OR2_X1 \V3/V3/A3/A1/M4/_0_  (.A1(\V3/V3/A3/A1/M4/c1 ),
    .A2(\V3/V3/A3/A1/M4/c2 ),
    .ZN(\V3/V3/A3/c1 ));
 AND2_X1 \V3/V3/A3/A2/M1/M1/_0_  (.A1(\V3/V3/v4 [4]),
    .A2(\V3/V3/c3 ),
    .ZN(\V3/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M1/M1/_1_  (.A(\V3/V3/v4 [4]),
    .B(\V3/V3/c3 ),
    .Z(\V3/V3/A3/A2/M1/s1 ));
 AND2_X1 \V3/V3/A3/A2/M1/M2/_0_  (.A1(\V3/V3/A3/A2/M1/s1 ),
    .A2(\V3/V3/A3/c1 ),
    .ZN(\V3/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M1/M2/_1_  (.A(\V3/V3/A3/A2/M1/s1 ),
    .B(\V3/V3/A3/c1 ),
    .Z(\V3/v3 [12]));
 OR2_X1 \V3/V3/A3/A2/M1/_0_  (.A1(\V3/V3/A3/A2/M1/c1 ),
    .A2(\V3/V3/A3/A2/M1/c2 ),
    .ZN(\V3/V3/A3/A2/c1 ));
 AND2_X1 \V3/V3/A3/A2/M2/M1/_0_  (.A1(\V3/V3/v4 [5]),
    .A2(ground),
    .ZN(\V3/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M2/M1/_1_  (.A(\V3/V3/v4 [5]),
    .B(ground),
    .Z(\V3/V3/A3/A2/M2/s1 ));
 AND2_X1 \V3/V3/A3/A2/M2/M2/_0_  (.A1(\V3/V3/A3/A2/M2/s1 ),
    .A2(\V3/V3/A3/A2/c1 ),
    .ZN(\V3/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M2/M2/_1_  (.A(\V3/V3/A3/A2/M2/s1 ),
    .B(\V3/V3/A3/A2/c1 ),
    .Z(\V3/v3 [13]));
 OR2_X1 \V3/V3/A3/A2/M2/_0_  (.A1(\V3/V3/A3/A2/M2/c1 ),
    .A2(\V3/V3/A3/A2/M2/c2 ),
    .ZN(\V3/V3/A3/A2/c2 ));
 AND2_X1 \V3/V3/A3/A2/M3/M1/_0_  (.A1(\V3/V3/v4 [6]),
    .A2(ground),
    .ZN(\V3/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M3/M1/_1_  (.A(\V3/V3/v4 [6]),
    .B(ground),
    .Z(\V3/V3/A3/A2/M3/s1 ));
 AND2_X1 \V3/V3/A3/A2/M3/M2/_0_  (.A1(\V3/V3/A3/A2/M3/s1 ),
    .A2(\V3/V3/A3/A2/c2 ),
    .ZN(\V3/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M3/M2/_1_  (.A(\V3/V3/A3/A2/M3/s1 ),
    .B(\V3/V3/A3/A2/c2 ),
    .Z(\V3/v3 [14]));
 OR2_X1 \V3/V3/A3/A2/M3/_0_  (.A1(\V3/V3/A3/A2/M3/c1 ),
    .A2(\V3/V3/A3/A2/M3/c2 ),
    .ZN(\V3/V3/A3/A2/c3 ));
 AND2_X1 \V3/V3/A3/A2/M4/M1/_0_  (.A1(\V3/V3/v4 [7]),
    .A2(ground),
    .ZN(\V3/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M4/M1/_1_  (.A(\V3/V3/v4 [7]),
    .B(ground),
    .Z(\V3/V3/A3/A2/M4/s1 ));
 AND2_X1 \V3/V3/A3/A2/M4/M2/_0_  (.A1(\V3/V3/A3/A2/M4/s1 ),
    .A2(\V3/V3/A3/A2/c3 ),
    .ZN(\V3/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M4/M2/_1_  (.A(\V3/V3/A3/A2/M4/s1 ),
    .B(\V3/V3/A3/A2/c3 ),
    .Z(\V3/v3 [15]));
 OR2_X1 \V3/V3/A3/A2/M4/_0_  (.A1(\V3/V3/A3/A2/M4/c1 ),
    .A2(\V3/V3/A3/A2/M4/c2 ),
    .ZN(\V3/V3/overflow ));
 AND2_X1 \V3/V3/V1/A1/M1/M1/_0_  (.A1(\V3/V3/V1/v2 [0]),
    .A2(\V3/V3/V1/v3 [0]),
    .ZN(\V3/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M1/M1/_1_  (.A(\V3/V3/V1/v2 [0]),
    .B(\V3/V3/V1/v3 [0]),
    .Z(\V3/V3/V1/A1/M1/s1 ));
 AND2_X1 \V3/V3/V1/A1/M1/M2/_0_  (.A1(\V3/V3/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M1/M2/_1_  (.A(\V3/V3/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/V1/s1 [0]));
 OR2_X1 \V3/V3/V1/A1/M1/_0_  (.A1(\V3/V3/V1/A1/M1/c1 ),
    .A2(\V3/V3/V1/A1/M1/c2 ),
    .ZN(\V3/V3/V1/A1/c1 ));
 AND2_X1 \V3/V3/V1/A1/M2/M1/_0_  (.A1(\V3/V3/V1/v2 [1]),
    .A2(\V3/V3/V1/v3 [1]),
    .ZN(\V3/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M2/M1/_1_  (.A(\V3/V3/V1/v2 [1]),
    .B(\V3/V3/V1/v3 [1]),
    .Z(\V3/V3/V1/A1/M2/s1 ));
 AND2_X1 \V3/V3/V1/A1/M2/M2/_0_  (.A1(\V3/V3/V1/A1/M2/s1 ),
    .A2(\V3/V3/V1/A1/c1 ),
    .ZN(\V3/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M2/M2/_1_  (.A(\V3/V3/V1/A1/M2/s1 ),
    .B(\V3/V3/V1/A1/c1 ),
    .Z(\V3/V3/V1/s1 [1]));
 OR2_X1 \V3/V3/V1/A1/M2/_0_  (.A1(\V3/V3/V1/A1/M2/c1 ),
    .A2(\V3/V3/V1/A1/M2/c2 ),
    .ZN(\V3/V3/V1/A1/c2 ));
 AND2_X1 \V3/V3/V1/A1/M3/M1/_0_  (.A1(\V3/V3/V1/v2 [2]),
    .A2(\V3/V3/V1/v3 [2]),
    .ZN(\V3/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M3/M1/_1_  (.A(\V3/V3/V1/v2 [2]),
    .B(\V3/V3/V1/v3 [2]),
    .Z(\V3/V3/V1/A1/M3/s1 ));
 AND2_X1 \V3/V3/V1/A1/M3/M2/_0_  (.A1(\V3/V3/V1/A1/M3/s1 ),
    .A2(\V3/V3/V1/A1/c2 ),
    .ZN(\V3/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M3/M2/_1_  (.A(\V3/V3/V1/A1/M3/s1 ),
    .B(\V3/V3/V1/A1/c2 ),
    .Z(\V3/V3/V1/s1 [2]));
 OR2_X1 \V3/V3/V1/A1/M3/_0_  (.A1(\V3/V3/V1/A1/M3/c1 ),
    .A2(\V3/V3/V1/A1/M3/c2 ),
    .ZN(\V3/V3/V1/A1/c3 ));
 AND2_X1 \V3/V3/V1/A1/M4/M1/_0_  (.A1(\V3/V3/V1/v2 [3]),
    .A2(\V3/V3/V1/v3 [3]),
    .ZN(\V3/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M4/M1/_1_  (.A(\V3/V3/V1/v2 [3]),
    .B(\V3/V3/V1/v3 [3]),
    .Z(\V3/V3/V1/A1/M4/s1 ));
 AND2_X1 \V3/V3/V1/A1/M4/M2/_0_  (.A1(\V3/V3/V1/A1/M4/s1 ),
    .A2(\V3/V3/V1/A1/c3 ),
    .ZN(\V3/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M4/M2/_1_  (.A(\V3/V3/V1/A1/M4/s1 ),
    .B(\V3/V3/V1/A1/c3 ),
    .Z(\V3/V3/V1/s1 [3]));
 OR2_X1 \V3/V3/V1/A1/M4/_0_  (.A1(\V3/V3/V1/A1/M4/c1 ),
    .A2(\V3/V3/V1/A1/M4/c2 ),
    .ZN(\V3/V3/V1/c1 ));
 AND2_X1 \V3/V3/V1/A2/M1/M1/_0_  (.A1(\V3/V3/V1/s1 [0]),
    .A2(\V3/V3/V1/v1 [2]),
    .ZN(\V3/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M1/M1/_1_  (.A(\V3/V3/V1/s1 [0]),
    .B(\V3/V3/V1/v1 [2]),
    .Z(\V3/V3/V1/A2/M1/s1 ));
 AND2_X1 \V3/V3/V1/A2/M1/M2/_0_  (.A1(\V3/V3/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M1/M2/_1_  (.A(\V3/V3/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/v3 [2]));
 OR2_X1 \V3/V3/V1/A2/M1/_0_  (.A1(\V3/V3/V1/A2/M1/c1 ),
    .A2(\V3/V3/V1/A2/M1/c2 ),
    .ZN(\V3/V3/V1/A2/c1 ));
 AND2_X1 \V3/V3/V1/A2/M2/M1/_0_  (.A1(\V3/V3/V1/s1 [1]),
    .A2(\V3/V3/V1/v1 [3]),
    .ZN(\V3/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M2/M1/_1_  (.A(\V3/V3/V1/s1 [1]),
    .B(\V3/V3/V1/v1 [3]),
    .Z(\V3/V3/V1/A2/M2/s1 ));
 AND2_X1 \V3/V3/V1/A2/M2/M2/_0_  (.A1(\V3/V3/V1/A2/M2/s1 ),
    .A2(\V3/V3/V1/A2/c1 ),
    .ZN(\V3/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M2/M2/_1_  (.A(\V3/V3/V1/A2/M2/s1 ),
    .B(\V3/V3/V1/A2/c1 ),
    .Z(\V3/v3 [3]));
 OR2_X1 \V3/V3/V1/A2/M2/_0_  (.A1(\V3/V3/V1/A2/M2/c1 ),
    .A2(\V3/V3/V1/A2/M2/c2 ),
    .ZN(\V3/V3/V1/A2/c2 ));
 AND2_X1 \V3/V3/V1/A2/M3/M1/_0_  (.A1(\V3/V3/V1/s1 [2]),
    .A2(ground),
    .ZN(\V3/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M3/M1/_1_  (.A(\V3/V3/V1/s1 [2]),
    .B(ground),
    .Z(\V3/V3/V1/A2/M3/s1 ));
 AND2_X1 \V3/V3/V1/A2/M3/M2/_0_  (.A1(\V3/V3/V1/A2/M3/s1 ),
    .A2(\V3/V3/V1/A2/c2 ),
    .ZN(\V3/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M3/M2/_1_  (.A(\V3/V3/V1/A2/M3/s1 ),
    .B(\V3/V3/V1/A2/c2 ),
    .Z(\V3/V3/V1/s2 [2]));
 OR2_X1 \V3/V3/V1/A2/M3/_0_  (.A1(\V3/V3/V1/A2/M3/c1 ),
    .A2(\V3/V3/V1/A2/M3/c2 ),
    .ZN(\V3/V3/V1/A2/c3 ));
 AND2_X1 \V3/V3/V1/A2/M4/M1/_0_  (.A1(\V3/V3/V1/s1 [3]),
    .A2(ground),
    .ZN(\V3/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M4/M1/_1_  (.A(\V3/V3/V1/s1 [3]),
    .B(ground),
    .Z(\V3/V3/V1/A2/M4/s1 ));
 AND2_X1 \V3/V3/V1/A2/M4/M2/_0_  (.A1(\V3/V3/V1/A2/M4/s1 ),
    .A2(\V3/V3/V1/A2/c3 ),
    .ZN(\V3/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M4/M2/_1_  (.A(\V3/V3/V1/A2/M4/s1 ),
    .B(\V3/V3/V1/A2/c3 ),
    .Z(\V3/V3/V1/s2 [3]));
 OR2_X1 \V3/V3/V1/A2/M4/_0_  (.A1(\V3/V3/V1/A2/M4/c1 ),
    .A2(\V3/V3/V1/A2/M4/c2 ),
    .ZN(\V3/V3/V1/c2 ));
 AND2_X1 \V3/V3/V1/A3/M1/M1/_0_  (.A1(\V3/V3/V1/v4 [0]),
    .A2(\V3/V3/V1/s2 [2]),
    .ZN(\V3/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M1/M1/_1_  (.A(\V3/V3/V1/v4 [0]),
    .B(\V3/V3/V1/s2 [2]),
    .Z(\V3/V3/V1/A3/M1/s1 ));
 AND2_X1 \V3/V3/V1/A3/M1/M2/_0_  (.A1(\V3/V3/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M1/M2/_1_  (.A(\V3/V3/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v1 [4]));
 OR2_X1 \V3/V3/V1/A3/M1/_0_  (.A1(\V3/V3/V1/A3/M1/c1 ),
    .A2(\V3/V3/V1/A3/M1/c2 ),
    .ZN(\V3/V3/V1/A3/c1 ));
 AND2_X1 \V3/V3/V1/A3/M2/M1/_0_  (.A1(\V3/V3/V1/v4 [1]),
    .A2(\V3/V3/V1/s2 [3]),
    .ZN(\V3/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M2/M1/_1_  (.A(\V3/V3/V1/v4 [1]),
    .B(\V3/V3/V1/s2 [3]),
    .Z(\V3/V3/V1/A3/M2/s1 ));
 AND2_X1 \V3/V3/V1/A3/M2/M2/_0_  (.A1(\V3/V3/V1/A3/M2/s1 ),
    .A2(\V3/V3/V1/A3/c1 ),
    .ZN(\V3/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M2/M2/_1_  (.A(\V3/V3/V1/A3/M2/s1 ),
    .B(\V3/V3/V1/A3/c1 ),
    .Z(\V3/V3/v1 [5]));
 OR2_X1 \V3/V3/V1/A3/M2/_0_  (.A1(\V3/V3/V1/A3/M2/c1 ),
    .A2(\V3/V3/V1/A3/M2/c2 ),
    .ZN(\V3/V3/V1/A3/c2 ));
 AND2_X1 \V3/V3/V1/A3/M3/M1/_0_  (.A1(\V3/V3/V1/v4 [2]),
    .A2(\V3/V3/V1/c3 ),
    .ZN(\V3/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M3/M1/_1_  (.A(\V3/V3/V1/v4 [2]),
    .B(\V3/V3/V1/c3 ),
    .Z(\V3/V3/V1/A3/M3/s1 ));
 AND2_X1 \V3/V3/V1/A3/M3/M2/_0_  (.A1(\V3/V3/V1/A3/M3/s1 ),
    .A2(\V3/V3/V1/A3/c2 ),
    .ZN(\V3/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M3/M2/_1_  (.A(\V3/V3/V1/A3/M3/s1 ),
    .B(\V3/V3/V1/A3/c2 ),
    .Z(\V3/V3/v1 [6]));
 OR2_X1 \V3/V3/V1/A3/M3/_0_  (.A1(\V3/V3/V1/A3/M3/c1 ),
    .A2(\V3/V3/V1/A3/M3/c2 ),
    .ZN(\V3/V3/V1/A3/c3 ));
 AND2_X1 \V3/V3/V1/A3/M4/M1/_0_  (.A1(\V3/V3/V1/v4 [3]),
    .A2(ground),
    .ZN(\V3/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M4/M1/_1_  (.A(\V3/V3/V1/v4 [3]),
    .B(ground),
    .Z(\V3/V3/V1/A3/M4/s1 ));
 AND2_X1 \V3/V3/V1/A3/M4/M2/_0_  (.A1(\V3/V3/V1/A3/M4/s1 ),
    .A2(\V3/V3/V1/A3/c3 ),
    .ZN(\V3/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M4/M2/_1_  (.A(\V3/V3/V1/A3/M4/s1 ),
    .B(\V3/V3/V1/A3/c3 ),
    .Z(\V3/V3/v1 [7]));
 OR2_X1 \V3/V3/V1/A3/M4/_0_  (.A1(\V3/V3/V1/A3/M4/c1 ),
    .A2(\V3/V3/V1/A3/M4/c2 ),
    .ZN(\V3/V3/V1/overflow ));
 AND2_X1 \V3/V3/V1/V1/HA1/_0_  (.A1(\V3/V3/V1/V1/w2 ),
    .A2(\V3/V3/V1/V1/w1 ),
    .ZN(\V3/V3/V1/V1/w4 ));
 XOR2_X2 \V3/V3/V1/V1/HA1/_1_  (.A(\V3/V3/V1/V1/w2 ),
    .B(\V3/V3/V1/V1/w1 ),
    .Z(\V3/v3 [1]));
 AND2_X1 \V3/V3/V1/V1/HA2/_0_  (.A1(\V3/V3/V1/V1/w4 ),
    .A2(\V3/V3/V1/V1/w3 ),
    .ZN(\V3/V3/V1/v1 [3]));
 XOR2_X2 \V3/V3/V1/V1/HA2/_1_  (.A(\V3/V3/V1/V1/w4 ),
    .B(\V3/V3/V1/V1/w3 ),
    .Z(\V3/V3/V1/v1 [2]));
 AND2_X1 \V3/V3/V1/V1/_0_  (.A1(A[0]),
    .A2(B[24]),
    .ZN(\V3/v3 [0]));
 AND2_X1 \V3/V3/V1/V1/_1_  (.A1(A[0]),
    .A2(B[25]),
    .ZN(\V3/V3/V1/V1/w1 ));
 AND2_X1 \V3/V3/V1/V1/_2_  (.A1(B[24]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V1/w2 ));
 AND2_X1 \V3/V3/V1/V1/_3_  (.A1(B[25]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V1/w3 ));
 AND2_X1 \V3/V3/V1/V2/HA1/_0_  (.A1(\V3/V3/V1/V2/w2 ),
    .A2(\V3/V3/V1/V2/w1 ),
    .ZN(\V3/V3/V1/V2/w4 ));
 XOR2_X2 \V3/V3/V1/V2/HA1/_1_  (.A(\V3/V3/V1/V2/w2 ),
    .B(\V3/V3/V1/V2/w1 ),
    .Z(\V3/V3/V1/v2 [1]));
 AND2_X1 \V3/V3/V1/V2/HA2/_0_  (.A1(\V3/V3/V1/V2/w4 ),
    .A2(\V3/V3/V1/V2/w3 ),
    .ZN(\V3/V3/V1/v2 [3]));
 XOR2_X2 \V3/V3/V1/V2/HA2/_1_  (.A(\V3/V3/V1/V2/w4 ),
    .B(\V3/V3/V1/V2/w3 ),
    .Z(\V3/V3/V1/v2 [2]));
 AND2_X1 \V3/V3/V1/V2/_0_  (.A1(A[2]),
    .A2(B[24]),
    .ZN(\V3/V3/V1/v2 [0]));
 AND2_X1 \V3/V3/V1/V2/_1_  (.A1(A[2]),
    .A2(B[25]),
    .ZN(\V3/V3/V1/V2/w1 ));
 AND2_X1 \V3/V3/V1/V2/_2_  (.A1(B[24]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V2/w2 ));
 AND2_X1 \V3/V3/V1/V2/_3_  (.A1(B[25]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V2/w3 ));
 AND2_X1 \V3/V3/V1/V3/HA1/_0_  (.A1(\V3/V3/V1/V3/w2 ),
    .A2(\V3/V3/V1/V3/w1 ),
    .ZN(\V3/V3/V1/V3/w4 ));
 XOR2_X2 \V3/V3/V1/V3/HA1/_1_  (.A(\V3/V3/V1/V3/w2 ),
    .B(\V3/V3/V1/V3/w1 ),
    .Z(\V3/V3/V1/v3 [1]));
 AND2_X1 \V3/V3/V1/V3/HA2/_0_  (.A1(\V3/V3/V1/V3/w4 ),
    .A2(\V3/V3/V1/V3/w3 ),
    .ZN(\V3/V3/V1/v3 [3]));
 XOR2_X2 \V3/V3/V1/V3/HA2/_1_  (.A(\V3/V3/V1/V3/w4 ),
    .B(\V3/V3/V1/V3/w3 ),
    .Z(\V3/V3/V1/v3 [2]));
 AND2_X1 \V3/V3/V1/V3/_0_  (.A1(A[0]),
    .A2(B[26]),
    .ZN(\V3/V3/V1/v3 [0]));
 AND2_X1 \V3/V3/V1/V3/_1_  (.A1(A[0]),
    .A2(B[27]),
    .ZN(\V3/V3/V1/V3/w1 ));
 AND2_X1 \V3/V3/V1/V3/_2_  (.A1(B[26]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V3/w2 ));
 AND2_X1 \V3/V3/V1/V3/_3_  (.A1(B[27]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V3/w3 ));
 AND2_X1 \V3/V3/V1/V4/HA1/_0_  (.A1(\V3/V3/V1/V4/w2 ),
    .A2(\V3/V3/V1/V4/w1 ),
    .ZN(\V3/V3/V1/V4/w4 ));
 XOR2_X2 \V3/V3/V1/V4/HA1/_1_  (.A(\V3/V3/V1/V4/w2 ),
    .B(\V3/V3/V1/V4/w1 ),
    .Z(\V3/V3/V1/v4 [1]));
 AND2_X1 \V3/V3/V1/V4/HA2/_0_  (.A1(\V3/V3/V1/V4/w4 ),
    .A2(\V3/V3/V1/V4/w3 ),
    .ZN(\V3/V3/V1/v4 [3]));
 XOR2_X2 \V3/V3/V1/V4/HA2/_1_  (.A(\V3/V3/V1/V4/w4 ),
    .B(\V3/V3/V1/V4/w3 ),
    .Z(\V3/V3/V1/v4 [2]));
 AND2_X1 \V3/V3/V1/V4/_0_  (.A1(A[2]),
    .A2(B[26]),
    .ZN(\V3/V3/V1/v4 [0]));
 AND2_X1 \V3/V3/V1/V4/_1_  (.A1(A[2]),
    .A2(B[27]),
    .ZN(\V3/V3/V1/V4/w1 ));
 AND2_X1 \V3/V3/V1/V4/_2_  (.A1(B[26]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V4/w2 ));
 AND2_X1 \V3/V3/V1/V4/_3_  (.A1(B[27]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V4/w3 ));
 OR2_X1 \V3/V3/V1/_0_  (.A1(\V3/V3/V1/c1 ),
    .A2(\V3/V3/V1/c2 ),
    .ZN(\V3/V3/V1/c3 ));
 AND2_X1 \V3/V3/V2/A1/M1/M1/_0_  (.A1(\V3/V3/V2/v2 [0]),
    .A2(\V3/V3/V2/v3 [0]),
    .ZN(\V3/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M1/M1/_1_  (.A(\V3/V3/V2/v2 [0]),
    .B(\V3/V3/V2/v3 [0]),
    .Z(\V3/V3/V2/A1/M1/s1 ));
 AND2_X1 \V3/V3/V2/A1/M1/M2/_0_  (.A1(\V3/V3/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M1/M2/_1_  (.A(\V3/V3/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/V2/s1 [0]));
 OR2_X1 \V3/V3/V2/A1/M1/_0_  (.A1(\V3/V3/V2/A1/M1/c1 ),
    .A2(\V3/V3/V2/A1/M1/c2 ),
    .ZN(\V3/V3/V2/A1/c1 ));
 AND2_X1 \V3/V3/V2/A1/M2/M1/_0_  (.A1(\V3/V3/V2/v2 [1]),
    .A2(\V3/V3/V2/v3 [1]),
    .ZN(\V3/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M2/M1/_1_  (.A(\V3/V3/V2/v2 [1]),
    .B(\V3/V3/V2/v3 [1]),
    .Z(\V3/V3/V2/A1/M2/s1 ));
 AND2_X1 \V3/V3/V2/A1/M2/M2/_0_  (.A1(\V3/V3/V2/A1/M2/s1 ),
    .A2(\V3/V3/V2/A1/c1 ),
    .ZN(\V3/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M2/M2/_1_  (.A(\V3/V3/V2/A1/M2/s1 ),
    .B(\V3/V3/V2/A1/c1 ),
    .Z(\V3/V3/V2/s1 [1]));
 OR2_X1 \V3/V3/V2/A1/M2/_0_  (.A1(\V3/V3/V2/A1/M2/c1 ),
    .A2(\V3/V3/V2/A1/M2/c2 ),
    .ZN(\V3/V3/V2/A1/c2 ));
 AND2_X1 \V3/V3/V2/A1/M3/M1/_0_  (.A1(\V3/V3/V2/v2 [2]),
    .A2(\V3/V3/V2/v3 [2]),
    .ZN(\V3/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M3/M1/_1_  (.A(\V3/V3/V2/v2 [2]),
    .B(\V3/V3/V2/v3 [2]),
    .Z(\V3/V3/V2/A1/M3/s1 ));
 AND2_X1 \V3/V3/V2/A1/M3/M2/_0_  (.A1(\V3/V3/V2/A1/M3/s1 ),
    .A2(\V3/V3/V2/A1/c2 ),
    .ZN(\V3/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M3/M2/_1_  (.A(\V3/V3/V2/A1/M3/s1 ),
    .B(\V3/V3/V2/A1/c2 ),
    .Z(\V3/V3/V2/s1 [2]));
 OR2_X1 \V3/V3/V2/A1/M3/_0_  (.A1(\V3/V3/V2/A1/M3/c1 ),
    .A2(\V3/V3/V2/A1/M3/c2 ),
    .ZN(\V3/V3/V2/A1/c3 ));
 AND2_X1 \V3/V3/V2/A1/M4/M1/_0_  (.A1(\V3/V3/V2/v2 [3]),
    .A2(\V3/V3/V2/v3 [3]),
    .ZN(\V3/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M4/M1/_1_  (.A(\V3/V3/V2/v2 [3]),
    .B(\V3/V3/V2/v3 [3]),
    .Z(\V3/V3/V2/A1/M4/s1 ));
 AND2_X1 \V3/V3/V2/A1/M4/M2/_0_  (.A1(\V3/V3/V2/A1/M4/s1 ),
    .A2(\V3/V3/V2/A1/c3 ),
    .ZN(\V3/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M4/M2/_1_  (.A(\V3/V3/V2/A1/M4/s1 ),
    .B(\V3/V3/V2/A1/c3 ),
    .Z(\V3/V3/V2/s1 [3]));
 OR2_X1 \V3/V3/V2/A1/M4/_0_  (.A1(\V3/V3/V2/A1/M4/c1 ),
    .A2(\V3/V3/V2/A1/M4/c2 ),
    .ZN(\V3/V3/V2/c1 ));
 AND2_X1 \V3/V3/V2/A2/M1/M1/_0_  (.A1(\V3/V3/V2/s1 [0]),
    .A2(\V3/V3/V2/v1 [2]),
    .ZN(\V3/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M1/M1/_1_  (.A(\V3/V3/V2/s1 [0]),
    .B(\V3/V3/V2/v1 [2]),
    .Z(\V3/V3/V2/A2/M1/s1 ));
 AND2_X1 \V3/V3/V2/A2/M1/M2/_0_  (.A1(\V3/V3/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M1/M2/_1_  (.A(\V3/V3/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v2 [2]));
 OR2_X1 \V3/V3/V2/A2/M1/_0_  (.A1(\V3/V3/V2/A2/M1/c1 ),
    .A2(\V3/V3/V2/A2/M1/c2 ),
    .ZN(\V3/V3/V2/A2/c1 ));
 AND2_X1 \V3/V3/V2/A2/M2/M1/_0_  (.A1(\V3/V3/V2/s1 [1]),
    .A2(\V3/V3/V2/v1 [3]),
    .ZN(\V3/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M2/M1/_1_  (.A(\V3/V3/V2/s1 [1]),
    .B(\V3/V3/V2/v1 [3]),
    .Z(\V3/V3/V2/A2/M2/s1 ));
 AND2_X1 \V3/V3/V2/A2/M2/M2/_0_  (.A1(\V3/V3/V2/A2/M2/s1 ),
    .A2(\V3/V3/V2/A2/c1 ),
    .ZN(\V3/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M2/M2/_1_  (.A(\V3/V3/V2/A2/M2/s1 ),
    .B(\V3/V3/V2/A2/c1 ),
    .Z(\V3/V3/v2 [3]));
 OR2_X1 \V3/V3/V2/A2/M2/_0_  (.A1(\V3/V3/V2/A2/M2/c1 ),
    .A2(\V3/V3/V2/A2/M2/c2 ),
    .ZN(\V3/V3/V2/A2/c2 ));
 AND2_X1 \V3/V3/V2/A2/M3/M1/_0_  (.A1(\V3/V3/V2/s1 [2]),
    .A2(ground),
    .ZN(\V3/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M3/M1/_1_  (.A(\V3/V3/V2/s1 [2]),
    .B(ground),
    .Z(\V3/V3/V2/A2/M3/s1 ));
 AND2_X1 \V3/V3/V2/A2/M3/M2/_0_  (.A1(\V3/V3/V2/A2/M3/s1 ),
    .A2(\V3/V3/V2/A2/c2 ),
    .ZN(\V3/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M3/M2/_1_  (.A(\V3/V3/V2/A2/M3/s1 ),
    .B(\V3/V3/V2/A2/c2 ),
    .Z(\V3/V3/V2/s2 [2]));
 OR2_X1 \V3/V3/V2/A2/M3/_0_  (.A1(\V3/V3/V2/A2/M3/c1 ),
    .A2(\V3/V3/V2/A2/M3/c2 ),
    .ZN(\V3/V3/V2/A2/c3 ));
 AND2_X1 \V3/V3/V2/A2/M4/M1/_0_  (.A1(\V3/V3/V2/s1 [3]),
    .A2(ground),
    .ZN(\V3/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M4/M1/_1_  (.A(\V3/V3/V2/s1 [3]),
    .B(ground),
    .Z(\V3/V3/V2/A2/M4/s1 ));
 AND2_X1 \V3/V3/V2/A2/M4/M2/_0_  (.A1(\V3/V3/V2/A2/M4/s1 ),
    .A2(\V3/V3/V2/A2/c3 ),
    .ZN(\V3/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M4/M2/_1_  (.A(\V3/V3/V2/A2/M4/s1 ),
    .B(\V3/V3/V2/A2/c3 ),
    .Z(\V3/V3/V2/s2 [3]));
 OR2_X1 \V3/V3/V2/A2/M4/_0_  (.A1(\V3/V3/V2/A2/M4/c1 ),
    .A2(\V3/V3/V2/A2/M4/c2 ),
    .ZN(\V3/V3/V2/c2 ));
 AND2_X1 \V3/V3/V2/A3/M1/M1/_0_  (.A1(\V3/V3/V2/v4 [0]),
    .A2(\V3/V3/V2/s2 [2]),
    .ZN(\V3/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M1/M1/_1_  (.A(\V3/V3/V2/v4 [0]),
    .B(\V3/V3/V2/s2 [2]),
    .Z(\V3/V3/V2/A3/M1/s1 ));
 AND2_X1 \V3/V3/V2/A3/M1/M2/_0_  (.A1(\V3/V3/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M1/M2/_1_  (.A(\V3/V3/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v2 [4]));
 OR2_X1 \V3/V3/V2/A3/M1/_0_  (.A1(\V3/V3/V2/A3/M1/c1 ),
    .A2(\V3/V3/V2/A3/M1/c2 ),
    .ZN(\V3/V3/V2/A3/c1 ));
 AND2_X1 \V3/V3/V2/A3/M2/M1/_0_  (.A1(\V3/V3/V2/v4 [1]),
    .A2(\V3/V3/V2/s2 [3]),
    .ZN(\V3/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M2/M1/_1_  (.A(\V3/V3/V2/v4 [1]),
    .B(\V3/V3/V2/s2 [3]),
    .Z(\V3/V3/V2/A3/M2/s1 ));
 AND2_X1 \V3/V3/V2/A3/M2/M2/_0_  (.A1(\V3/V3/V2/A3/M2/s1 ),
    .A2(\V3/V3/V2/A3/c1 ),
    .ZN(\V3/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M2/M2/_1_  (.A(\V3/V3/V2/A3/M2/s1 ),
    .B(\V3/V3/V2/A3/c1 ),
    .Z(\V3/V3/v2 [5]));
 OR2_X1 \V3/V3/V2/A3/M2/_0_  (.A1(\V3/V3/V2/A3/M2/c1 ),
    .A2(\V3/V3/V2/A3/M2/c2 ),
    .ZN(\V3/V3/V2/A3/c2 ));
 AND2_X1 \V3/V3/V2/A3/M3/M1/_0_  (.A1(\V3/V3/V2/v4 [2]),
    .A2(\V3/V3/V2/c3 ),
    .ZN(\V3/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M3/M1/_1_  (.A(\V3/V3/V2/v4 [2]),
    .B(\V3/V3/V2/c3 ),
    .Z(\V3/V3/V2/A3/M3/s1 ));
 AND2_X1 \V3/V3/V2/A3/M3/M2/_0_  (.A1(\V3/V3/V2/A3/M3/s1 ),
    .A2(\V3/V3/V2/A3/c2 ),
    .ZN(\V3/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M3/M2/_1_  (.A(\V3/V3/V2/A3/M3/s1 ),
    .B(\V3/V3/V2/A3/c2 ),
    .Z(\V3/V3/v2 [6]));
 OR2_X1 \V3/V3/V2/A3/M3/_0_  (.A1(\V3/V3/V2/A3/M3/c1 ),
    .A2(\V3/V3/V2/A3/M3/c2 ),
    .ZN(\V3/V3/V2/A3/c3 ));
 AND2_X1 \V3/V3/V2/A3/M4/M1/_0_  (.A1(\V3/V3/V2/v4 [3]),
    .A2(ground),
    .ZN(\V3/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M4/M1/_1_  (.A(\V3/V3/V2/v4 [3]),
    .B(ground),
    .Z(\V3/V3/V2/A3/M4/s1 ));
 AND2_X1 \V3/V3/V2/A3/M4/M2/_0_  (.A1(\V3/V3/V2/A3/M4/s1 ),
    .A2(\V3/V3/V2/A3/c3 ),
    .ZN(\V3/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M4/M2/_1_  (.A(\V3/V3/V2/A3/M4/s1 ),
    .B(\V3/V3/V2/A3/c3 ),
    .Z(\V3/V3/v2 [7]));
 OR2_X1 \V3/V3/V2/A3/M4/_0_  (.A1(\V3/V3/V2/A3/M4/c1 ),
    .A2(\V3/V3/V2/A3/M4/c2 ),
    .ZN(\V3/V3/V2/overflow ));
 AND2_X1 \V3/V3/V2/V1/HA1/_0_  (.A1(\V3/V3/V2/V1/w2 ),
    .A2(\V3/V3/V2/V1/w1 ),
    .ZN(\V3/V3/V2/V1/w4 ));
 XOR2_X2 \V3/V3/V2/V1/HA1/_1_  (.A(\V3/V3/V2/V1/w2 ),
    .B(\V3/V3/V2/V1/w1 ),
    .Z(\V3/V3/v2 [1]));
 AND2_X1 \V3/V3/V2/V1/HA2/_0_  (.A1(\V3/V3/V2/V1/w4 ),
    .A2(\V3/V3/V2/V1/w3 ),
    .ZN(\V3/V3/V2/v1 [3]));
 XOR2_X2 \V3/V3/V2/V1/HA2/_1_  (.A(\V3/V3/V2/V1/w4 ),
    .B(\V3/V3/V2/V1/w3 ),
    .Z(\V3/V3/V2/v1 [2]));
 AND2_X1 \V3/V3/V2/V1/_0_  (.A1(A[4]),
    .A2(B[24]),
    .ZN(\V3/V3/v2 [0]));
 AND2_X1 \V3/V3/V2/V1/_1_  (.A1(A[4]),
    .A2(B[25]),
    .ZN(\V3/V3/V2/V1/w1 ));
 AND2_X1 \V3/V3/V2/V1/_2_  (.A1(B[24]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V1/w2 ));
 AND2_X1 \V3/V3/V2/V1/_3_  (.A1(B[25]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V1/w3 ));
 AND2_X1 \V3/V3/V2/V2/HA1/_0_  (.A1(\V3/V3/V2/V2/w2 ),
    .A2(\V3/V3/V2/V2/w1 ),
    .ZN(\V3/V3/V2/V2/w4 ));
 XOR2_X2 \V3/V3/V2/V2/HA1/_1_  (.A(\V3/V3/V2/V2/w2 ),
    .B(\V3/V3/V2/V2/w1 ),
    .Z(\V3/V3/V2/v2 [1]));
 AND2_X1 \V3/V3/V2/V2/HA2/_0_  (.A1(\V3/V3/V2/V2/w4 ),
    .A2(\V3/V3/V2/V2/w3 ),
    .ZN(\V3/V3/V2/v2 [3]));
 XOR2_X2 \V3/V3/V2/V2/HA2/_1_  (.A(\V3/V3/V2/V2/w4 ),
    .B(\V3/V3/V2/V2/w3 ),
    .Z(\V3/V3/V2/v2 [2]));
 AND2_X1 \V3/V3/V2/V2/_0_  (.A1(A[6]),
    .A2(B[24]),
    .ZN(\V3/V3/V2/v2 [0]));
 AND2_X1 \V3/V3/V2/V2/_1_  (.A1(A[6]),
    .A2(B[25]),
    .ZN(\V3/V3/V2/V2/w1 ));
 AND2_X1 \V3/V3/V2/V2/_2_  (.A1(B[24]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V2/w2 ));
 AND2_X1 \V3/V3/V2/V2/_3_  (.A1(B[25]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V2/w3 ));
 AND2_X1 \V3/V3/V2/V3/HA1/_0_  (.A1(\V3/V3/V2/V3/w2 ),
    .A2(\V3/V3/V2/V3/w1 ),
    .ZN(\V3/V3/V2/V3/w4 ));
 XOR2_X2 \V3/V3/V2/V3/HA1/_1_  (.A(\V3/V3/V2/V3/w2 ),
    .B(\V3/V3/V2/V3/w1 ),
    .Z(\V3/V3/V2/v3 [1]));
 AND2_X1 \V3/V3/V2/V3/HA2/_0_  (.A1(\V3/V3/V2/V3/w4 ),
    .A2(\V3/V3/V2/V3/w3 ),
    .ZN(\V3/V3/V2/v3 [3]));
 XOR2_X2 \V3/V3/V2/V3/HA2/_1_  (.A(\V3/V3/V2/V3/w4 ),
    .B(\V3/V3/V2/V3/w3 ),
    .Z(\V3/V3/V2/v3 [2]));
 AND2_X1 \V3/V3/V2/V3/_0_  (.A1(A[4]),
    .A2(B[26]),
    .ZN(\V3/V3/V2/v3 [0]));
 AND2_X1 \V3/V3/V2/V3/_1_  (.A1(A[4]),
    .A2(B[27]),
    .ZN(\V3/V3/V2/V3/w1 ));
 AND2_X1 \V3/V3/V2/V3/_2_  (.A1(B[26]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V3/w2 ));
 AND2_X1 \V3/V3/V2/V3/_3_  (.A1(B[27]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V3/w3 ));
 AND2_X1 \V3/V3/V2/V4/HA1/_0_  (.A1(\V3/V3/V2/V4/w2 ),
    .A2(\V3/V3/V2/V4/w1 ),
    .ZN(\V3/V3/V2/V4/w4 ));
 XOR2_X2 \V3/V3/V2/V4/HA1/_1_  (.A(\V3/V3/V2/V4/w2 ),
    .B(\V3/V3/V2/V4/w1 ),
    .Z(\V3/V3/V2/v4 [1]));
 AND2_X1 \V3/V3/V2/V4/HA2/_0_  (.A1(\V3/V3/V2/V4/w4 ),
    .A2(\V3/V3/V2/V4/w3 ),
    .ZN(\V3/V3/V2/v4 [3]));
 XOR2_X2 \V3/V3/V2/V4/HA2/_1_  (.A(\V3/V3/V2/V4/w4 ),
    .B(\V3/V3/V2/V4/w3 ),
    .Z(\V3/V3/V2/v4 [2]));
 AND2_X1 \V3/V3/V2/V4/_0_  (.A1(A[6]),
    .A2(B[26]),
    .ZN(\V3/V3/V2/v4 [0]));
 AND2_X1 \V3/V3/V2/V4/_1_  (.A1(A[6]),
    .A2(B[27]),
    .ZN(\V3/V3/V2/V4/w1 ));
 AND2_X1 \V3/V3/V2/V4/_2_  (.A1(B[26]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V4/w2 ));
 AND2_X1 \V3/V3/V2/V4/_3_  (.A1(B[27]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V4/w3 ));
 OR2_X1 \V3/V3/V2/_0_  (.A1(\V3/V3/V2/c1 ),
    .A2(\V3/V3/V2/c2 ),
    .ZN(\V3/V3/V2/c3 ));
 AND2_X1 \V3/V3/V3/A1/M1/M1/_0_  (.A1(\V3/V3/V3/v2 [0]),
    .A2(\V3/V3/V3/v3 [0]),
    .ZN(\V3/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M1/M1/_1_  (.A(\V3/V3/V3/v2 [0]),
    .B(\V3/V3/V3/v3 [0]),
    .Z(\V3/V3/V3/A1/M1/s1 ));
 AND2_X1 \V3/V3/V3/A1/M1/M2/_0_  (.A1(\V3/V3/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M1/M2/_1_  (.A(\V3/V3/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/V3/s1 [0]));
 OR2_X1 \V3/V3/V3/A1/M1/_0_  (.A1(\V3/V3/V3/A1/M1/c1 ),
    .A2(\V3/V3/V3/A1/M1/c2 ),
    .ZN(\V3/V3/V3/A1/c1 ));
 AND2_X1 \V3/V3/V3/A1/M2/M1/_0_  (.A1(\V3/V3/V3/v2 [1]),
    .A2(\V3/V3/V3/v3 [1]),
    .ZN(\V3/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M2/M1/_1_  (.A(\V3/V3/V3/v2 [1]),
    .B(\V3/V3/V3/v3 [1]),
    .Z(\V3/V3/V3/A1/M2/s1 ));
 AND2_X1 \V3/V3/V3/A1/M2/M2/_0_  (.A1(\V3/V3/V3/A1/M2/s1 ),
    .A2(\V3/V3/V3/A1/c1 ),
    .ZN(\V3/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M2/M2/_1_  (.A(\V3/V3/V3/A1/M2/s1 ),
    .B(\V3/V3/V3/A1/c1 ),
    .Z(\V3/V3/V3/s1 [1]));
 OR2_X1 \V3/V3/V3/A1/M2/_0_  (.A1(\V3/V3/V3/A1/M2/c1 ),
    .A2(\V3/V3/V3/A1/M2/c2 ),
    .ZN(\V3/V3/V3/A1/c2 ));
 AND2_X1 \V3/V3/V3/A1/M3/M1/_0_  (.A1(\V3/V3/V3/v2 [2]),
    .A2(\V3/V3/V3/v3 [2]),
    .ZN(\V3/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M3/M1/_1_  (.A(\V3/V3/V3/v2 [2]),
    .B(\V3/V3/V3/v3 [2]),
    .Z(\V3/V3/V3/A1/M3/s1 ));
 AND2_X1 \V3/V3/V3/A1/M3/M2/_0_  (.A1(\V3/V3/V3/A1/M3/s1 ),
    .A2(\V3/V3/V3/A1/c2 ),
    .ZN(\V3/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M3/M2/_1_  (.A(\V3/V3/V3/A1/M3/s1 ),
    .B(\V3/V3/V3/A1/c2 ),
    .Z(\V3/V3/V3/s1 [2]));
 OR2_X1 \V3/V3/V3/A1/M3/_0_  (.A1(\V3/V3/V3/A1/M3/c1 ),
    .A2(\V3/V3/V3/A1/M3/c2 ),
    .ZN(\V3/V3/V3/A1/c3 ));
 AND2_X1 \V3/V3/V3/A1/M4/M1/_0_  (.A1(\V3/V3/V3/v2 [3]),
    .A2(\V3/V3/V3/v3 [3]),
    .ZN(\V3/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M4/M1/_1_  (.A(\V3/V3/V3/v2 [3]),
    .B(\V3/V3/V3/v3 [3]),
    .Z(\V3/V3/V3/A1/M4/s1 ));
 AND2_X1 \V3/V3/V3/A1/M4/M2/_0_  (.A1(\V3/V3/V3/A1/M4/s1 ),
    .A2(\V3/V3/V3/A1/c3 ),
    .ZN(\V3/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M4/M2/_1_  (.A(\V3/V3/V3/A1/M4/s1 ),
    .B(\V3/V3/V3/A1/c3 ),
    .Z(\V3/V3/V3/s1 [3]));
 OR2_X1 \V3/V3/V3/A1/M4/_0_  (.A1(\V3/V3/V3/A1/M4/c1 ),
    .A2(\V3/V3/V3/A1/M4/c2 ),
    .ZN(\V3/V3/V3/c1 ));
 AND2_X1 \V3/V3/V3/A2/M1/M1/_0_  (.A1(\V3/V3/V3/s1 [0]),
    .A2(\V3/V3/V3/v1 [2]),
    .ZN(\V3/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M1/M1/_1_  (.A(\V3/V3/V3/s1 [0]),
    .B(\V3/V3/V3/v1 [2]),
    .Z(\V3/V3/V3/A2/M1/s1 ));
 AND2_X1 \V3/V3/V3/A2/M1/M2/_0_  (.A1(\V3/V3/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M1/M2/_1_  (.A(\V3/V3/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v3 [2]));
 OR2_X1 \V3/V3/V3/A2/M1/_0_  (.A1(\V3/V3/V3/A2/M1/c1 ),
    .A2(\V3/V3/V3/A2/M1/c2 ),
    .ZN(\V3/V3/V3/A2/c1 ));
 AND2_X1 \V3/V3/V3/A2/M2/M1/_0_  (.A1(\V3/V3/V3/s1 [1]),
    .A2(\V3/V3/V3/v1 [3]),
    .ZN(\V3/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M2/M1/_1_  (.A(\V3/V3/V3/s1 [1]),
    .B(\V3/V3/V3/v1 [3]),
    .Z(\V3/V3/V3/A2/M2/s1 ));
 AND2_X1 \V3/V3/V3/A2/M2/M2/_0_  (.A1(\V3/V3/V3/A2/M2/s1 ),
    .A2(\V3/V3/V3/A2/c1 ),
    .ZN(\V3/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M2/M2/_1_  (.A(\V3/V3/V3/A2/M2/s1 ),
    .B(\V3/V3/V3/A2/c1 ),
    .Z(\V3/V3/v3 [3]));
 OR2_X1 \V3/V3/V3/A2/M2/_0_  (.A1(\V3/V3/V3/A2/M2/c1 ),
    .A2(\V3/V3/V3/A2/M2/c2 ),
    .ZN(\V3/V3/V3/A2/c2 ));
 AND2_X1 \V3/V3/V3/A2/M3/M1/_0_  (.A1(\V3/V3/V3/s1 [2]),
    .A2(ground),
    .ZN(\V3/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M3/M1/_1_  (.A(\V3/V3/V3/s1 [2]),
    .B(ground),
    .Z(\V3/V3/V3/A2/M3/s1 ));
 AND2_X1 \V3/V3/V3/A2/M3/M2/_0_  (.A1(\V3/V3/V3/A2/M3/s1 ),
    .A2(\V3/V3/V3/A2/c2 ),
    .ZN(\V3/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M3/M2/_1_  (.A(\V3/V3/V3/A2/M3/s1 ),
    .B(\V3/V3/V3/A2/c2 ),
    .Z(\V3/V3/V3/s2 [2]));
 OR2_X1 \V3/V3/V3/A2/M3/_0_  (.A1(\V3/V3/V3/A2/M3/c1 ),
    .A2(\V3/V3/V3/A2/M3/c2 ),
    .ZN(\V3/V3/V3/A2/c3 ));
 AND2_X1 \V3/V3/V3/A2/M4/M1/_0_  (.A1(\V3/V3/V3/s1 [3]),
    .A2(ground),
    .ZN(\V3/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M4/M1/_1_  (.A(\V3/V3/V3/s1 [3]),
    .B(ground),
    .Z(\V3/V3/V3/A2/M4/s1 ));
 AND2_X1 \V3/V3/V3/A2/M4/M2/_0_  (.A1(\V3/V3/V3/A2/M4/s1 ),
    .A2(\V3/V3/V3/A2/c3 ),
    .ZN(\V3/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M4/M2/_1_  (.A(\V3/V3/V3/A2/M4/s1 ),
    .B(\V3/V3/V3/A2/c3 ),
    .Z(\V3/V3/V3/s2 [3]));
 OR2_X1 \V3/V3/V3/A2/M4/_0_  (.A1(\V3/V3/V3/A2/M4/c1 ),
    .A2(\V3/V3/V3/A2/M4/c2 ),
    .ZN(\V3/V3/V3/c2 ));
 AND2_X1 \V3/V3/V3/A3/M1/M1/_0_  (.A1(\V3/V3/V3/v4 [0]),
    .A2(\V3/V3/V3/s2 [2]),
    .ZN(\V3/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M1/M1/_1_  (.A(\V3/V3/V3/v4 [0]),
    .B(\V3/V3/V3/s2 [2]),
    .Z(\V3/V3/V3/A3/M1/s1 ));
 AND2_X1 \V3/V3/V3/A3/M1/M2/_0_  (.A1(\V3/V3/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M1/M2/_1_  (.A(\V3/V3/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v3 [4]));
 OR2_X1 \V3/V3/V3/A3/M1/_0_  (.A1(\V3/V3/V3/A3/M1/c1 ),
    .A2(\V3/V3/V3/A3/M1/c2 ),
    .ZN(\V3/V3/V3/A3/c1 ));
 AND2_X1 \V3/V3/V3/A3/M2/M1/_0_  (.A1(\V3/V3/V3/v4 [1]),
    .A2(\V3/V3/V3/s2 [3]),
    .ZN(\V3/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M2/M1/_1_  (.A(\V3/V3/V3/v4 [1]),
    .B(\V3/V3/V3/s2 [3]),
    .Z(\V3/V3/V3/A3/M2/s1 ));
 AND2_X1 \V3/V3/V3/A3/M2/M2/_0_  (.A1(\V3/V3/V3/A3/M2/s1 ),
    .A2(\V3/V3/V3/A3/c1 ),
    .ZN(\V3/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M2/M2/_1_  (.A(\V3/V3/V3/A3/M2/s1 ),
    .B(\V3/V3/V3/A3/c1 ),
    .Z(\V3/V3/v3 [5]));
 OR2_X1 \V3/V3/V3/A3/M2/_0_  (.A1(\V3/V3/V3/A3/M2/c1 ),
    .A2(\V3/V3/V3/A3/M2/c2 ),
    .ZN(\V3/V3/V3/A3/c2 ));
 AND2_X1 \V3/V3/V3/A3/M3/M1/_0_  (.A1(\V3/V3/V3/v4 [2]),
    .A2(\V3/V3/V3/c3 ),
    .ZN(\V3/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M3/M1/_1_  (.A(\V3/V3/V3/v4 [2]),
    .B(\V3/V3/V3/c3 ),
    .Z(\V3/V3/V3/A3/M3/s1 ));
 AND2_X1 \V3/V3/V3/A3/M3/M2/_0_  (.A1(\V3/V3/V3/A3/M3/s1 ),
    .A2(\V3/V3/V3/A3/c2 ),
    .ZN(\V3/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M3/M2/_1_  (.A(\V3/V3/V3/A3/M3/s1 ),
    .B(\V3/V3/V3/A3/c2 ),
    .Z(\V3/V3/v3 [6]));
 OR2_X1 \V3/V3/V3/A3/M3/_0_  (.A1(\V3/V3/V3/A3/M3/c1 ),
    .A2(\V3/V3/V3/A3/M3/c2 ),
    .ZN(\V3/V3/V3/A3/c3 ));
 AND2_X1 \V3/V3/V3/A3/M4/M1/_0_  (.A1(\V3/V3/V3/v4 [3]),
    .A2(ground),
    .ZN(\V3/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M4/M1/_1_  (.A(\V3/V3/V3/v4 [3]),
    .B(ground),
    .Z(\V3/V3/V3/A3/M4/s1 ));
 AND2_X1 \V3/V3/V3/A3/M4/M2/_0_  (.A1(\V3/V3/V3/A3/M4/s1 ),
    .A2(\V3/V3/V3/A3/c3 ),
    .ZN(\V3/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M4/M2/_1_  (.A(\V3/V3/V3/A3/M4/s1 ),
    .B(\V3/V3/V3/A3/c3 ),
    .Z(\V3/V3/v3 [7]));
 OR2_X1 \V3/V3/V3/A3/M4/_0_  (.A1(\V3/V3/V3/A3/M4/c1 ),
    .A2(\V3/V3/V3/A3/M4/c2 ),
    .ZN(\V3/V3/V3/overflow ));
 AND2_X1 \V3/V3/V3/V1/HA1/_0_  (.A1(\V3/V3/V3/V1/w2 ),
    .A2(\V3/V3/V3/V1/w1 ),
    .ZN(\V3/V3/V3/V1/w4 ));
 XOR2_X2 \V3/V3/V3/V1/HA1/_1_  (.A(\V3/V3/V3/V1/w2 ),
    .B(\V3/V3/V3/V1/w1 ),
    .Z(\V3/V3/v3 [1]));
 AND2_X1 \V3/V3/V3/V1/HA2/_0_  (.A1(\V3/V3/V3/V1/w4 ),
    .A2(\V3/V3/V3/V1/w3 ),
    .ZN(\V3/V3/V3/v1 [3]));
 XOR2_X2 \V3/V3/V3/V1/HA2/_1_  (.A(\V3/V3/V3/V1/w4 ),
    .B(\V3/V3/V3/V1/w3 ),
    .Z(\V3/V3/V3/v1 [2]));
 AND2_X1 \V3/V3/V3/V1/_0_  (.A1(A[0]),
    .A2(B[28]),
    .ZN(\V3/V3/v3 [0]));
 AND2_X1 \V3/V3/V3/V1/_1_  (.A1(A[0]),
    .A2(B[29]),
    .ZN(\V3/V3/V3/V1/w1 ));
 AND2_X1 \V3/V3/V3/V1/_2_  (.A1(B[28]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V1/w2 ));
 AND2_X1 \V3/V3/V3/V1/_3_  (.A1(B[29]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V1/w3 ));
 AND2_X1 \V3/V3/V3/V2/HA1/_0_  (.A1(\V3/V3/V3/V2/w2 ),
    .A2(\V3/V3/V3/V2/w1 ),
    .ZN(\V3/V3/V3/V2/w4 ));
 XOR2_X2 \V3/V3/V3/V2/HA1/_1_  (.A(\V3/V3/V3/V2/w2 ),
    .B(\V3/V3/V3/V2/w1 ),
    .Z(\V3/V3/V3/v2 [1]));
 AND2_X1 \V3/V3/V3/V2/HA2/_0_  (.A1(\V3/V3/V3/V2/w4 ),
    .A2(\V3/V3/V3/V2/w3 ),
    .ZN(\V3/V3/V3/v2 [3]));
 XOR2_X2 \V3/V3/V3/V2/HA2/_1_  (.A(\V3/V3/V3/V2/w4 ),
    .B(\V3/V3/V3/V2/w3 ),
    .Z(\V3/V3/V3/v2 [2]));
 AND2_X1 \V3/V3/V3/V2/_0_  (.A1(A[2]),
    .A2(B[28]),
    .ZN(\V3/V3/V3/v2 [0]));
 AND2_X1 \V3/V3/V3/V2/_1_  (.A1(A[2]),
    .A2(B[29]),
    .ZN(\V3/V3/V3/V2/w1 ));
 AND2_X1 \V3/V3/V3/V2/_2_  (.A1(B[28]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V2/w2 ));
 AND2_X1 \V3/V3/V3/V2/_3_  (.A1(B[29]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V2/w3 ));
 AND2_X1 \V3/V3/V3/V3/HA1/_0_  (.A1(\V3/V3/V3/V3/w2 ),
    .A2(\V3/V3/V3/V3/w1 ),
    .ZN(\V3/V3/V3/V3/w4 ));
 XOR2_X2 \V3/V3/V3/V3/HA1/_1_  (.A(\V3/V3/V3/V3/w2 ),
    .B(\V3/V3/V3/V3/w1 ),
    .Z(\V3/V3/V3/v3 [1]));
 AND2_X1 \V3/V3/V3/V3/HA2/_0_  (.A1(\V3/V3/V3/V3/w4 ),
    .A2(\V3/V3/V3/V3/w3 ),
    .ZN(\V3/V3/V3/v3 [3]));
 XOR2_X2 \V3/V3/V3/V3/HA2/_1_  (.A(\V3/V3/V3/V3/w4 ),
    .B(\V3/V3/V3/V3/w3 ),
    .Z(\V3/V3/V3/v3 [2]));
 AND2_X1 \V3/V3/V3/V3/_0_  (.A1(A[0]),
    .A2(B[30]),
    .ZN(\V3/V3/V3/v3 [0]));
 AND2_X1 \V3/V3/V3/V3/_1_  (.A1(A[0]),
    .A2(B[31]),
    .ZN(\V3/V3/V3/V3/w1 ));
 AND2_X1 \V3/V3/V3/V3/_2_  (.A1(B[30]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V3/w2 ));
 AND2_X1 \V3/V3/V3/V3/_3_  (.A1(B[31]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V3/w3 ));
 AND2_X1 \V3/V3/V3/V4/HA1/_0_  (.A1(\V3/V3/V3/V4/w2 ),
    .A2(\V3/V3/V3/V4/w1 ),
    .ZN(\V3/V3/V3/V4/w4 ));
 XOR2_X2 \V3/V3/V3/V4/HA1/_1_  (.A(\V3/V3/V3/V4/w2 ),
    .B(\V3/V3/V3/V4/w1 ),
    .Z(\V3/V3/V3/v4 [1]));
 AND2_X1 \V3/V3/V3/V4/HA2/_0_  (.A1(\V3/V3/V3/V4/w4 ),
    .A2(\V3/V3/V3/V4/w3 ),
    .ZN(\V3/V3/V3/v4 [3]));
 XOR2_X2 \V3/V3/V3/V4/HA2/_1_  (.A(\V3/V3/V3/V4/w4 ),
    .B(\V3/V3/V3/V4/w3 ),
    .Z(\V3/V3/V3/v4 [2]));
 AND2_X1 \V3/V3/V3/V4/_0_  (.A1(A[2]),
    .A2(B[30]),
    .ZN(\V3/V3/V3/v4 [0]));
 AND2_X1 \V3/V3/V3/V4/_1_  (.A1(A[2]),
    .A2(B[31]),
    .ZN(\V3/V3/V3/V4/w1 ));
 AND2_X1 \V3/V3/V3/V4/_2_  (.A1(B[30]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V4/w2 ));
 AND2_X1 \V3/V3/V3/V4/_3_  (.A1(B[31]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V4/w3 ));
 OR2_X1 \V3/V3/V3/_0_  (.A1(\V3/V3/V3/c1 ),
    .A2(\V3/V3/V3/c2 ),
    .ZN(\V3/V3/V3/c3 ));
 AND2_X1 \V3/V3/V4/A1/M1/M1/_0_  (.A1(\V3/V3/V4/v2 [0]),
    .A2(\V3/V3/V4/v3 [0]),
    .ZN(\V3/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M1/M1/_1_  (.A(\V3/V3/V4/v2 [0]),
    .B(\V3/V3/V4/v3 [0]),
    .Z(\V3/V3/V4/A1/M1/s1 ));
 AND2_X1 \V3/V3/V4/A1/M1/M2/_0_  (.A1(\V3/V3/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M1/M2/_1_  (.A(\V3/V3/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/V4/s1 [0]));
 OR2_X1 \V3/V3/V4/A1/M1/_0_  (.A1(\V3/V3/V4/A1/M1/c1 ),
    .A2(\V3/V3/V4/A1/M1/c2 ),
    .ZN(\V3/V3/V4/A1/c1 ));
 AND2_X1 \V3/V3/V4/A1/M2/M1/_0_  (.A1(\V3/V3/V4/v2 [1]),
    .A2(\V3/V3/V4/v3 [1]),
    .ZN(\V3/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M2/M1/_1_  (.A(\V3/V3/V4/v2 [1]),
    .B(\V3/V3/V4/v3 [1]),
    .Z(\V3/V3/V4/A1/M2/s1 ));
 AND2_X1 \V3/V3/V4/A1/M2/M2/_0_  (.A1(\V3/V3/V4/A1/M2/s1 ),
    .A2(\V3/V3/V4/A1/c1 ),
    .ZN(\V3/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M2/M2/_1_  (.A(\V3/V3/V4/A1/M2/s1 ),
    .B(\V3/V3/V4/A1/c1 ),
    .Z(\V3/V3/V4/s1 [1]));
 OR2_X1 \V3/V3/V4/A1/M2/_0_  (.A1(\V3/V3/V4/A1/M2/c1 ),
    .A2(\V3/V3/V4/A1/M2/c2 ),
    .ZN(\V3/V3/V4/A1/c2 ));
 AND2_X1 \V3/V3/V4/A1/M3/M1/_0_  (.A1(\V3/V3/V4/v2 [2]),
    .A2(\V3/V3/V4/v3 [2]),
    .ZN(\V3/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M3/M1/_1_  (.A(\V3/V3/V4/v2 [2]),
    .B(\V3/V3/V4/v3 [2]),
    .Z(\V3/V3/V4/A1/M3/s1 ));
 AND2_X1 \V3/V3/V4/A1/M3/M2/_0_  (.A1(\V3/V3/V4/A1/M3/s1 ),
    .A2(\V3/V3/V4/A1/c2 ),
    .ZN(\V3/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M3/M2/_1_  (.A(\V3/V3/V4/A1/M3/s1 ),
    .B(\V3/V3/V4/A1/c2 ),
    .Z(\V3/V3/V4/s1 [2]));
 OR2_X1 \V3/V3/V4/A1/M3/_0_  (.A1(\V3/V3/V4/A1/M3/c1 ),
    .A2(\V3/V3/V4/A1/M3/c2 ),
    .ZN(\V3/V3/V4/A1/c3 ));
 AND2_X1 \V3/V3/V4/A1/M4/M1/_0_  (.A1(\V3/V3/V4/v2 [3]),
    .A2(\V3/V3/V4/v3 [3]),
    .ZN(\V3/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M4/M1/_1_  (.A(\V3/V3/V4/v2 [3]),
    .B(\V3/V3/V4/v3 [3]),
    .Z(\V3/V3/V4/A1/M4/s1 ));
 AND2_X1 \V3/V3/V4/A1/M4/M2/_0_  (.A1(\V3/V3/V4/A1/M4/s1 ),
    .A2(\V3/V3/V4/A1/c3 ),
    .ZN(\V3/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M4/M2/_1_  (.A(\V3/V3/V4/A1/M4/s1 ),
    .B(\V3/V3/V4/A1/c3 ),
    .Z(\V3/V3/V4/s1 [3]));
 OR2_X1 \V3/V3/V4/A1/M4/_0_  (.A1(\V3/V3/V4/A1/M4/c1 ),
    .A2(\V3/V3/V4/A1/M4/c2 ),
    .ZN(\V3/V3/V4/c1 ));
 AND2_X1 \V3/V3/V4/A2/M1/M1/_0_  (.A1(\V3/V3/V4/s1 [0]),
    .A2(\V3/V3/V4/v1 [2]),
    .ZN(\V3/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M1/M1/_1_  (.A(\V3/V3/V4/s1 [0]),
    .B(\V3/V3/V4/v1 [2]),
    .Z(\V3/V3/V4/A2/M1/s1 ));
 AND2_X1 \V3/V3/V4/A2/M1/M2/_0_  (.A1(\V3/V3/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M1/M2/_1_  (.A(\V3/V3/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v4 [2]));
 OR2_X1 \V3/V3/V4/A2/M1/_0_  (.A1(\V3/V3/V4/A2/M1/c1 ),
    .A2(\V3/V3/V4/A2/M1/c2 ),
    .ZN(\V3/V3/V4/A2/c1 ));
 AND2_X1 \V3/V3/V4/A2/M2/M1/_0_  (.A1(\V3/V3/V4/s1 [1]),
    .A2(\V3/V3/V4/v1 [3]),
    .ZN(\V3/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M2/M1/_1_  (.A(\V3/V3/V4/s1 [1]),
    .B(\V3/V3/V4/v1 [3]),
    .Z(\V3/V3/V4/A2/M2/s1 ));
 AND2_X1 \V3/V3/V4/A2/M2/M2/_0_  (.A1(\V3/V3/V4/A2/M2/s1 ),
    .A2(\V3/V3/V4/A2/c1 ),
    .ZN(\V3/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M2/M2/_1_  (.A(\V3/V3/V4/A2/M2/s1 ),
    .B(\V3/V3/V4/A2/c1 ),
    .Z(\V3/V3/v4 [3]));
 OR2_X1 \V3/V3/V4/A2/M2/_0_  (.A1(\V3/V3/V4/A2/M2/c1 ),
    .A2(\V3/V3/V4/A2/M2/c2 ),
    .ZN(\V3/V3/V4/A2/c2 ));
 AND2_X1 \V3/V3/V4/A2/M3/M1/_0_  (.A1(\V3/V3/V4/s1 [2]),
    .A2(ground),
    .ZN(\V3/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M3/M1/_1_  (.A(\V3/V3/V4/s1 [2]),
    .B(ground),
    .Z(\V3/V3/V4/A2/M3/s1 ));
 AND2_X1 \V3/V3/V4/A2/M3/M2/_0_  (.A1(\V3/V3/V4/A2/M3/s1 ),
    .A2(\V3/V3/V4/A2/c2 ),
    .ZN(\V3/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M3/M2/_1_  (.A(\V3/V3/V4/A2/M3/s1 ),
    .B(\V3/V3/V4/A2/c2 ),
    .Z(\V3/V3/V4/s2 [2]));
 OR2_X1 \V3/V3/V4/A2/M3/_0_  (.A1(\V3/V3/V4/A2/M3/c1 ),
    .A2(\V3/V3/V4/A2/M3/c2 ),
    .ZN(\V3/V3/V4/A2/c3 ));
 AND2_X1 \V3/V3/V4/A2/M4/M1/_0_  (.A1(\V3/V3/V4/s1 [3]),
    .A2(ground),
    .ZN(\V3/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M4/M1/_1_  (.A(\V3/V3/V4/s1 [3]),
    .B(ground),
    .Z(\V3/V3/V4/A2/M4/s1 ));
 AND2_X1 \V3/V3/V4/A2/M4/M2/_0_  (.A1(\V3/V3/V4/A2/M4/s1 ),
    .A2(\V3/V3/V4/A2/c3 ),
    .ZN(\V3/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M4/M2/_1_  (.A(\V3/V3/V4/A2/M4/s1 ),
    .B(\V3/V3/V4/A2/c3 ),
    .Z(\V3/V3/V4/s2 [3]));
 OR2_X1 \V3/V3/V4/A2/M4/_0_  (.A1(\V3/V3/V4/A2/M4/c1 ),
    .A2(\V3/V3/V4/A2/M4/c2 ),
    .ZN(\V3/V3/V4/c2 ));
 AND2_X1 \V3/V3/V4/A3/M1/M1/_0_  (.A1(\V3/V3/V4/v4 [0]),
    .A2(\V3/V3/V4/s2 [2]),
    .ZN(\V3/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M1/M1/_1_  (.A(\V3/V3/V4/v4 [0]),
    .B(\V3/V3/V4/s2 [2]),
    .Z(\V3/V3/V4/A3/M1/s1 ));
 AND2_X1 \V3/V3/V4/A3/M1/M2/_0_  (.A1(\V3/V3/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M1/M2/_1_  (.A(\V3/V3/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V3/v4 [4]));
 OR2_X1 \V3/V3/V4/A3/M1/_0_  (.A1(\V3/V3/V4/A3/M1/c1 ),
    .A2(\V3/V3/V4/A3/M1/c2 ),
    .ZN(\V3/V3/V4/A3/c1 ));
 AND2_X1 \V3/V3/V4/A3/M2/M1/_0_  (.A1(\V3/V3/V4/v4 [1]),
    .A2(\V3/V3/V4/s2 [3]),
    .ZN(\V3/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M2/M1/_1_  (.A(\V3/V3/V4/v4 [1]),
    .B(\V3/V3/V4/s2 [3]),
    .Z(\V3/V3/V4/A3/M2/s1 ));
 AND2_X1 \V3/V3/V4/A3/M2/M2/_0_  (.A1(\V3/V3/V4/A3/M2/s1 ),
    .A2(\V3/V3/V4/A3/c1 ),
    .ZN(\V3/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M2/M2/_1_  (.A(\V3/V3/V4/A3/M2/s1 ),
    .B(\V3/V3/V4/A3/c1 ),
    .Z(\V3/V3/v4 [5]));
 OR2_X1 \V3/V3/V4/A3/M2/_0_  (.A1(\V3/V3/V4/A3/M2/c1 ),
    .A2(\V3/V3/V4/A3/M2/c2 ),
    .ZN(\V3/V3/V4/A3/c2 ));
 AND2_X1 \V3/V3/V4/A3/M3/M1/_0_  (.A1(\V3/V3/V4/v4 [2]),
    .A2(\V3/V3/V4/c3 ),
    .ZN(\V3/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M3/M1/_1_  (.A(\V3/V3/V4/v4 [2]),
    .B(\V3/V3/V4/c3 ),
    .Z(\V3/V3/V4/A3/M3/s1 ));
 AND2_X1 \V3/V3/V4/A3/M3/M2/_0_  (.A1(\V3/V3/V4/A3/M3/s1 ),
    .A2(\V3/V3/V4/A3/c2 ),
    .ZN(\V3/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M3/M2/_1_  (.A(\V3/V3/V4/A3/M3/s1 ),
    .B(\V3/V3/V4/A3/c2 ),
    .Z(\V3/V3/v4 [6]));
 OR2_X1 \V3/V3/V4/A3/M3/_0_  (.A1(\V3/V3/V4/A3/M3/c1 ),
    .A2(\V3/V3/V4/A3/M3/c2 ),
    .ZN(\V3/V3/V4/A3/c3 ));
 AND2_X1 \V3/V3/V4/A3/M4/M1/_0_  (.A1(\V3/V3/V4/v4 [3]),
    .A2(ground),
    .ZN(\V3/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M4/M1/_1_  (.A(\V3/V3/V4/v4 [3]),
    .B(ground),
    .Z(\V3/V3/V4/A3/M4/s1 ));
 AND2_X1 \V3/V3/V4/A3/M4/M2/_0_  (.A1(\V3/V3/V4/A3/M4/s1 ),
    .A2(\V3/V3/V4/A3/c3 ),
    .ZN(\V3/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M4/M2/_1_  (.A(\V3/V3/V4/A3/M4/s1 ),
    .B(\V3/V3/V4/A3/c3 ),
    .Z(\V3/V3/v4 [7]));
 OR2_X1 \V3/V3/V4/A3/M4/_0_  (.A1(\V3/V3/V4/A3/M4/c1 ),
    .A2(\V3/V3/V4/A3/M4/c2 ),
    .ZN(\V3/V3/V4/overflow ));
 AND2_X1 \V3/V3/V4/V1/HA1/_0_  (.A1(\V3/V3/V4/V1/w2 ),
    .A2(\V3/V3/V4/V1/w1 ),
    .ZN(\V3/V3/V4/V1/w4 ));
 XOR2_X2 \V3/V3/V4/V1/HA1/_1_  (.A(\V3/V3/V4/V1/w2 ),
    .B(\V3/V3/V4/V1/w1 ),
    .Z(\V3/V3/v4 [1]));
 AND2_X1 \V3/V3/V4/V1/HA2/_0_  (.A1(\V3/V3/V4/V1/w4 ),
    .A2(\V3/V3/V4/V1/w3 ),
    .ZN(\V3/V3/V4/v1 [3]));
 XOR2_X2 \V3/V3/V4/V1/HA2/_1_  (.A(\V3/V3/V4/V1/w4 ),
    .B(\V3/V3/V4/V1/w3 ),
    .Z(\V3/V3/V4/v1 [2]));
 AND2_X1 \V3/V3/V4/V1/_0_  (.A1(A[4]),
    .A2(B[28]),
    .ZN(\V3/V3/v4 [0]));
 AND2_X1 \V3/V3/V4/V1/_1_  (.A1(A[4]),
    .A2(B[29]),
    .ZN(\V3/V3/V4/V1/w1 ));
 AND2_X1 \V3/V3/V4/V1/_2_  (.A1(B[28]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V1/w2 ));
 AND2_X1 \V3/V3/V4/V1/_3_  (.A1(B[29]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V1/w3 ));
 AND2_X1 \V3/V3/V4/V2/HA1/_0_  (.A1(\V3/V3/V4/V2/w2 ),
    .A2(\V3/V3/V4/V2/w1 ),
    .ZN(\V3/V3/V4/V2/w4 ));
 XOR2_X2 \V3/V3/V4/V2/HA1/_1_  (.A(\V3/V3/V4/V2/w2 ),
    .B(\V3/V3/V4/V2/w1 ),
    .Z(\V3/V3/V4/v2 [1]));
 AND2_X1 \V3/V3/V4/V2/HA2/_0_  (.A1(\V3/V3/V4/V2/w4 ),
    .A2(\V3/V3/V4/V2/w3 ),
    .ZN(\V3/V3/V4/v2 [3]));
 XOR2_X2 \V3/V3/V4/V2/HA2/_1_  (.A(\V3/V3/V4/V2/w4 ),
    .B(\V3/V3/V4/V2/w3 ),
    .Z(\V3/V3/V4/v2 [2]));
 AND2_X1 \V3/V3/V4/V2/_0_  (.A1(A[6]),
    .A2(B[28]),
    .ZN(\V3/V3/V4/v2 [0]));
 AND2_X1 \V3/V3/V4/V2/_1_  (.A1(A[6]),
    .A2(B[29]),
    .ZN(\V3/V3/V4/V2/w1 ));
 AND2_X1 \V3/V3/V4/V2/_2_  (.A1(B[28]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V2/w2 ));
 AND2_X1 \V3/V3/V4/V2/_3_  (.A1(B[29]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V2/w3 ));
 AND2_X1 \V3/V3/V4/V3/HA1/_0_  (.A1(\V3/V3/V4/V3/w2 ),
    .A2(\V3/V3/V4/V3/w1 ),
    .ZN(\V3/V3/V4/V3/w4 ));
 XOR2_X2 \V3/V3/V4/V3/HA1/_1_  (.A(\V3/V3/V4/V3/w2 ),
    .B(\V3/V3/V4/V3/w1 ),
    .Z(\V3/V3/V4/v3 [1]));
 AND2_X1 \V3/V3/V4/V3/HA2/_0_  (.A1(\V3/V3/V4/V3/w4 ),
    .A2(\V3/V3/V4/V3/w3 ),
    .ZN(\V3/V3/V4/v3 [3]));
 XOR2_X2 \V3/V3/V4/V3/HA2/_1_  (.A(\V3/V3/V4/V3/w4 ),
    .B(\V3/V3/V4/V3/w3 ),
    .Z(\V3/V3/V4/v3 [2]));
 AND2_X1 \V3/V3/V4/V3/_0_  (.A1(A[4]),
    .A2(B[30]),
    .ZN(\V3/V3/V4/v3 [0]));
 AND2_X1 \V3/V3/V4/V3/_1_  (.A1(A[4]),
    .A2(B[31]),
    .ZN(\V3/V3/V4/V3/w1 ));
 AND2_X1 \V3/V3/V4/V3/_2_  (.A1(B[30]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V3/w2 ));
 AND2_X1 \V3/V3/V4/V3/_3_  (.A1(B[31]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V3/w3 ));
 AND2_X1 \V3/V3/V4/V4/HA1/_0_  (.A1(\V3/V3/V4/V4/w2 ),
    .A2(\V3/V3/V4/V4/w1 ),
    .ZN(\V3/V3/V4/V4/w4 ));
 XOR2_X2 \V3/V3/V4/V4/HA1/_1_  (.A(\V3/V3/V4/V4/w2 ),
    .B(\V3/V3/V4/V4/w1 ),
    .Z(\V3/V3/V4/v4 [1]));
 AND2_X1 \V3/V3/V4/V4/HA2/_0_  (.A1(\V3/V3/V4/V4/w4 ),
    .A2(\V3/V3/V4/V4/w3 ),
    .ZN(\V3/V3/V4/v4 [3]));
 XOR2_X2 \V3/V3/V4/V4/HA2/_1_  (.A(\V3/V3/V4/V4/w4 ),
    .B(\V3/V3/V4/V4/w3 ),
    .Z(\V3/V3/V4/v4 [2]));
 AND2_X1 \V3/V3/V4/V4/_0_  (.A1(A[6]),
    .A2(B[30]),
    .ZN(\V3/V3/V4/v4 [0]));
 AND2_X1 \V3/V3/V4/V4/_1_  (.A1(A[6]),
    .A2(B[31]),
    .ZN(\V3/V3/V4/V4/w1 ));
 AND2_X1 \V3/V3/V4/V4/_2_  (.A1(B[30]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V4/w2 ));
 AND2_X1 \V3/V3/V4/V4/_3_  (.A1(B[31]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V4/w3 ));
 OR2_X1 \V3/V3/V4/_0_  (.A1(\V3/V3/V4/c1 ),
    .A2(\V3/V3/V4/c2 ),
    .ZN(\V3/V3/V4/c3 ));
 OR2_X1 \V3/V3/_0_  (.A1(\V3/V3/c1 ),
    .A2(\V3/V3/c2 ),
    .ZN(\V3/V3/c3 ));
 AND2_X1 \V3/V4/A1/A1/M1/M1/_0_  (.A1(\V3/V4/v2 [0]),
    .A2(\V3/V4/v3 [0]),
    .ZN(\V3/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M1/M1/_1_  (.A(\V3/V4/v2 [0]),
    .B(\V3/V4/v3 [0]),
    .Z(\V3/V4/A1/A1/M1/s1 ));
 AND2_X1 \V3/V4/A1/A1/M1/M2/_0_  (.A1(\V3/V4/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M1/M2/_1_  (.A(\V3/V4/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/s1 [0]));
 OR2_X1 \V3/V4/A1/A1/M1/_0_  (.A1(\V3/V4/A1/A1/M1/c1 ),
    .A2(\V3/V4/A1/A1/M1/c2 ),
    .ZN(\V3/V4/A1/A1/c1 ));
 AND2_X1 \V3/V4/A1/A1/M2/M1/_0_  (.A1(\V3/V4/v2 [1]),
    .A2(\V3/V4/v3 [1]),
    .ZN(\V3/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M2/M1/_1_  (.A(\V3/V4/v2 [1]),
    .B(\V3/V4/v3 [1]),
    .Z(\V3/V4/A1/A1/M2/s1 ));
 AND2_X1 \V3/V4/A1/A1/M2/M2/_0_  (.A1(\V3/V4/A1/A1/M2/s1 ),
    .A2(\V3/V4/A1/A1/c1 ),
    .ZN(\V3/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M2/M2/_1_  (.A(\V3/V4/A1/A1/M2/s1 ),
    .B(\V3/V4/A1/A1/c1 ),
    .Z(\V3/V4/s1 [1]));
 OR2_X1 \V3/V4/A1/A1/M2/_0_  (.A1(\V3/V4/A1/A1/M2/c1 ),
    .A2(\V3/V4/A1/A1/M2/c2 ),
    .ZN(\V3/V4/A1/A1/c2 ));
 AND2_X1 \V3/V4/A1/A1/M3/M1/_0_  (.A1(\V3/V4/v2 [2]),
    .A2(\V3/V4/v3 [2]),
    .ZN(\V3/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M3/M1/_1_  (.A(\V3/V4/v2 [2]),
    .B(\V3/V4/v3 [2]),
    .Z(\V3/V4/A1/A1/M3/s1 ));
 AND2_X1 \V3/V4/A1/A1/M3/M2/_0_  (.A1(\V3/V4/A1/A1/M3/s1 ),
    .A2(\V3/V4/A1/A1/c2 ),
    .ZN(\V3/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M3/M2/_1_  (.A(\V3/V4/A1/A1/M3/s1 ),
    .B(\V3/V4/A1/A1/c2 ),
    .Z(\V3/V4/s1 [2]));
 OR2_X1 \V3/V4/A1/A1/M3/_0_  (.A1(\V3/V4/A1/A1/M3/c1 ),
    .A2(\V3/V4/A1/A1/M3/c2 ),
    .ZN(\V3/V4/A1/A1/c3 ));
 AND2_X1 \V3/V4/A1/A1/M4/M1/_0_  (.A1(\V3/V4/v2 [3]),
    .A2(\V3/V4/v3 [3]),
    .ZN(\V3/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M4/M1/_1_  (.A(\V3/V4/v2 [3]),
    .B(\V3/V4/v3 [3]),
    .Z(\V3/V4/A1/A1/M4/s1 ));
 AND2_X1 \V3/V4/A1/A1/M4/M2/_0_  (.A1(\V3/V4/A1/A1/M4/s1 ),
    .A2(\V3/V4/A1/A1/c3 ),
    .ZN(\V3/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M4/M2/_1_  (.A(\V3/V4/A1/A1/M4/s1 ),
    .B(\V3/V4/A1/A1/c3 ),
    .Z(\V3/V4/s1 [3]));
 OR2_X1 \V3/V4/A1/A1/M4/_0_  (.A1(\V3/V4/A1/A1/M4/c1 ),
    .A2(\V3/V4/A1/A1/M4/c2 ),
    .ZN(\V3/V4/A1/c1 ));
 AND2_X1 \V3/V4/A1/A2/M1/M1/_0_  (.A1(\V3/V4/v2 [4]),
    .A2(\V3/V4/v3 [4]),
    .ZN(\V3/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M1/M1/_1_  (.A(\V3/V4/v2 [4]),
    .B(\V3/V4/v3 [4]),
    .Z(\V3/V4/A1/A2/M1/s1 ));
 AND2_X1 \V3/V4/A1/A2/M1/M2/_0_  (.A1(\V3/V4/A1/A2/M1/s1 ),
    .A2(\V3/V4/A1/c1 ),
    .ZN(\V3/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M1/M2/_1_  (.A(\V3/V4/A1/A2/M1/s1 ),
    .B(\V3/V4/A1/c1 ),
    .Z(\V3/V4/s1 [4]));
 OR2_X1 \V3/V4/A1/A2/M1/_0_  (.A1(\V3/V4/A1/A2/M1/c1 ),
    .A2(\V3/V4/A1/A2/M1/c2 ),
    .ZN(\V3/V4/A1/A2/c1 ));
 AND2_X1 \V3/V4/A1/A2/M2/M1/_0_  (.A1(\V3/V4/v2 [5]),
    .A2(\V3/V4/v3 [5]),
    .ZN(\V3/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M2/M1/_1_  (.A(\V3/V4/v2 [5]),
    .B(\V3/V4/v3 [5]),
    .Z(\V3/V4/A1/A2/M2/s1 ));
 AND2_X1 \V3/V4/A1/A2/M2/M2/_0_  (.A1(\V3/V4/A1/A2/M2/s1 ),
    .A2(\V3/V4/A1/A2/c1 ),
    .ZN(\V3/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M2/M2/_1_  (.A(\V3/V4/A1/A2/M2/s1 ),
    .B(\V3/V4/A1/A2/c1 ),
    .Z(\V3/V4/s1 [5]));
 OR2_X1 \V3/V4/A1/A2/M2/_0_  (.A1(\V3/V4/A1/A2/M2/c1 ),
    .A2(\V3/V4/A1/A2/M2/c2 ),
    .ZN(\V3/V4/A1/A2/c2 ));
 AND2_X1 \V3/V4/A1/A2/M3/M1/_0_  (.A1(\V3/V4/v2 [6]),
    .A2(\V3/V4/v3 [6]),
    .ZN(\V3/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M3/M1/_1_  (.A(\V3/V4/v2 [6]),
    .B(\V3/V4/v3 [6]),
    .Z(\V3/V4/A1/A2/M3/s1 ));
 AND2_X1 \V3/V4/A1/A2/M3/M2/_0_  (.A1(\V3/V4/A1/A2/M3/s1 ),
    .A2(\V3/V4/A1/A2/c2 ),
    .ZN(\V3/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M3/M2/_1_  (.A(\V3/V4/A1/A2/M3/s1 ),
    .B(\V3/V4/A1/A2/c2 ),
    .Z(\V3/V4/s1 [6]));
 OR2_X1 \V3/V4/A1/A2/M3/_0_  (.A1(\V3/V4/A1/A2/M3/c1 ),
    .A2(\V3/V4/A1/A2/M3/c2 ),
    .ZN(\V3/V4/A1/A2/c3 ));
 AND2_X1 \V3/V4/A1/A2/M4/M1/_0_  (.A1(\V3/V4/v2 [7]),
    .A2(\V3/V4/v3 [7]),
    .ZN(\V3/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M4/M1/_1_  (.A(\V3/V4/v2 [7]),
    .B(\V3/V4/v3 [7]),
    .Z(\V3/V4/A1/A2/M4/s1 ));
 AND2_X1 \V3/V4/A1/A2/M4/M2/_0_  (.A1(\V3/V4/A1/A2/M4/s1 ),
    .A2(\V3/V4/A1/A2/c3 ),
    .ZN(\V3/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M4/M2/_1_  (.A(\V3/V4/A1/A2/M4/s1 ),
    .B(\V3/V4/A1/A2/c3 ),
    .Z(\V3/V4/s1 [7]));
 OR2_X1 \V3/V4/A1/A2/M4/_0_  (.A1(\V3/V4/A1/A2/M4/c1 ),
    .A2(\V3/V4/A1/A2/M4/c2 ),
    .ZN(\V3/V4/c1 ));
 AND2_X1 \V3/V4/A2/A1/M1/M1/_0_  (.A1(\V3/V4/s1 [0]),
    .A2(\V3/V4/v1 [4]),
    .ZN(\V3/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M1/M1/_1_  (.A(\V3/V4/s1 [0]),
    .B(\V3/V4/v1 [4]),
    .Z(\V3/V4/A2/A1/M1/s1 ));
 AND2_X1 \V3/V4/A2/A1/M1/M2/_0_  (.A1(\V3/V4/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M1/M2/_1_  (.A(\V3/V4/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v4 [4]));
 OR2_X1 \V3/V4/A2/A1/M1/_0_  (.A1(\V3/V4/A2/A1/M1/c1 ),
    .A2(\V3/V4/A2/A1/M1/c2 ),
    .ZN(\V3/V4/A2/A1/c1 ));
 AND2_X1 \V3/V4/A2/A1/M2/M1/_0_  (.A1(\V3/V4/s1 [1]),
    .A2(\V3/V4/v1 [5]),
    .ZN(\V3/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M2/M1/_1_  (.A(\V3/V4/s1 [1]),
    .B(\V3/V4/v1 [5]),
    .Z(\V3/V4/A2/A1/M2/s1 ));
 AND2_X1 \V3/V4/A2/A1/M2/M2/_0_  (.A1(\V3/V4/A2/A1/M2/s1 ),
    .A2(\V3/V4/A2/A1/c1 ),
    .ZN(\V3/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M2/M2/_1_  (.A(\V3/V4/A2/A1/M2/s1 ),
    .B(\V3/V4/A2/A1/c1 ),
    .Z(\V3/v4 [5]));
 OR2_X1 \V3/V4/A2/A1/M2/_0_  (.A1(\V3/V4/A2/A1/M2/c1 ),
    .A2(\V3/V4/A2/A1/M2/c2 ),
    .ZN(\V3/V4/A2/A1/c2 ));
 AND2_X1 \V3/V4/A2/A1/M3/M1/_0_  (.A1(\V3/V4/s1 [2]),
    .A2(\V3/V4/v1 [6]),
    .ZN(\V3/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M3/M1/_1_  (.A(\V3/V4/s1 [2]),
    .B(\V3/V4/v1 [6]),
    .Z(\V3/V4/A2/A1/M3/s1 ));
 AND2_X1 \V3/V4/A2/A1/M3/M2/_0_  (.A1(\V3/V4/A2/A1/M3/s1 ),
    .A2(\V3/V4/A2/A1/c2 ),
    .ZN(\V3/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M3/M2/_1_  (.A(\V3/V4/A2/A1/M3/s1 ),
    .B(\V3/V4/A2/A1/c2 ),
    .Z(\V3/v4 [6]));
 OR2_X1 \V3/V4/A2/A1/M3/_0_  (.A1(\V3/V4/A2/A1/M3/c1 ),
    .A2(\V3/V4/A2/A1/M3/c2 ),
    .ZN(\V3/V4/A2/A1/c3 ));
 AND2_X1 \V3/V4/A2/A1/M4/M1/_0_  (.A1(\V3/V4/s1 [3]),
    .A2(\V3/V4/v1 [7]),
    .ZN(\V3/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M4/M1/_1_  (.A(\V3/V4/s1 [3]),
    .B(\V3/V4/v1 [7]),
    .Z(\V3/V4/A2/A1/M4/s1 ));
 AND2_X1 \V3/V4/A2/A1/M4/M2/_0_  (.A1(\V3/V4/A2/A1/M4/s1 ),
    .A2(\V3/V4/A2/A1/c3 ),
    .ZN(\V3/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M4/M2/_1_  (.A(\V3/V4/A2/A1/M4/s1 ),
    .B(\V3/V4/A2/A1/c3 ),
    .Z(\V3/v4 [7]));
 OR2_X1 \V3/V4/A2/A1/M4/_0_  (.A1(\V3/V4/A2/A1/M4/c1 ),
    .A2(\V3/V4/A2/A1/M4/c2 ),
    .ZN(\V3/V4/A2/c1 ));
 AND2_X1 \V3/V4/A2/A2/M1/M1/_0_  (.A1(\V3/V4/s1 [4]),
    .A2(ground),
    .ZN(\V3/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M1/M1/_1_  (.A(\V3/V4/s1 [4]),
    .B(ground),
    .Z(\V3/V4/A2/A2/M1/s1 ));
 AND2_X1 \V3/V4/A2/A2/M1/M2/_0_  (.A1(\V3/V4/A2/A2/M1/s1 ),
    .A2(\V3/V4/A2/c1 ),
    .ZN(\V3/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M1/M2/_1_  (.A(\V3/V4/A2/A2/M1/s1 ),
    .B(\V3/V4/A2/c1 ),
    .Z(\V3/V4/s2 [4]));
 OR2_X1 \V3/V4/A2/A2/M1/_0_  (.A1(\V3/V4/A2/A2/M1/c1 ),
    .A2(\V3/V4/A2/A2/M1/c2 ),
    .ZN(\V3/V4/A2/A2/c1 ));
 AND2_X1 \V3/V4/A2/A2/M2/M1/_0_  (.A1(\V3/V4/s1 [5]),
    .A2(ground),
    .ZN(\V3/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M2/M1/_1_  (.A(\V3/V4/s1 [5]),
    .B(ground),
    .Z(\V3/V4/A2/A2/M2/s1 ));
 AND2_X1 \V3/V4/A2/A2/M2/M2/_0_  (.A1(\V3/V4/A2/A2/M2/s1 ),
    .A2(\V3/V4/A2/A2/c1 ),
    .ZN(\V3/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M2/M2/_1_  (.A(\V3/V4/A2/A2/M2/s1 ),
    .B(\V3/V4/A2/A2/c1 ),
    .Z(\V3/V4/s2 [5]));
 OR2_X1 \V3/V4/A2/A2/M2/_0_  (.A1(\V3/V4/A2/A2/M2/c1 ),
    .A2(\V3/V4/A2/A2/M2/c2 ),
    .ZN(\V3/V4/A2/A2/c2 ));
 AND2_X1 \V3/V4/A2/A2/M3/M1/_0_  (.A1(\V3/V4/s1 [6]),
    .A2(ground),
    .ZN(\V3/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M3/M1/_1_  (.A(\V3/V4/s1 [6]),
    .B(ground),
    .Z(\V3/V4/A2/A2/M3/s1 ));
 AND2_X1 \V3/V4/A2/A2/M3/M2/_0_  (.A1(\V3/V4/A2/A2/M3/s1 ),
    .A2(\V3/V4/A2/A2/c2 ),
    .ZN(\V3/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M3/M2/_1_  (.A(\V3/V4/A2/A2/M3/s1 ),
    .B(\V3/V4/A2/A2/c2 ),
    .Z(\V3/V4/s2 [6]));
 OR2_X1 \V3/V4/A2/A2/M3/_0_  (.A1(\V3/V4/A2/A2/M3/c1 ),
    .A2(\V3/V4/A2/A2/M3/c2 ),
    .ZN(\V3/V4/A2/A2/c3 ));
 AND2_X1 \V3/V4/A2/A2/M4/M1/_0_  (.A1(\V3/V4/s1 [7]),
    .A2(ground),
    .ZN(\V3/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M4/M1/_1_  (.A(\V3/V4/s1 [7]),
    .B(ground),
    .Z(\V3/V4/A2/A2/M4/s1 ));
 AND2_X1 \V3/V4/A2/A2/M4/M2/_0_  (.A1(\V3/V4/A2/A2/M4/s1 ),
    .A2(\V3/V4/A2/A2/c3 ),
    .ZN(\V3/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M4/M2/_1_  (.A(\V3/V4/A2/A2/M4/s1 ),
    .B(\V3/V4/A2/A2/c3 ),
    .Z(\V3/V4/s2 [7]));
 OR2_X1 \V3/V4/A2/A2/M4/_0_  (.A1(\V3/V4/A2/A2/M4/c1 ),
    .A2(\V3/V4/A2/A2/M4/c2 ),
    .ZN(\V3/V4/c2 ));
 AND2_X1 \V3/V4/A3/A1/M1/M1/_0_  (.A1(\V3/V4/v4 [0]),
    .A2(\V3/V4/s2 [4]),
    .ZN(\V3/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M1/M1/_1_  (.A(\V3/V4/v4 [0]),
    .B(\V3/V4/s2 [4]),
    .Z(\V3/V4/A3/A1/M1/s1 ));
 AND2_X1 \V3/V4/A3/A1/M1/M2/_0_  (.A1(\V3/V4/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M1/M2/_1_  (.A(\V3/V4/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/v4 [8]));
 OR2_X1 \V3/V4/A3/A1/M1/_0_  (.A1(\V3/V4/A3/A1/M1/c1 ),
    .A2(\V3/V4/A3/A1/M1/c2 ),
    .ZN(\V3/V4/A3/A1/c1 ));
 AND2_X1 \V3/V4/A3/A1/M2/M1/_0_  (.A1(\V3/V4/v4 [1]),
    .A2(\V3/V4/s2 [5]),
    .ZN(\V3/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M2/M1/_1_  (.A(\V3/V4/v4 [1]),
    .B(\V3/V4/s2 [5]),
    .Z(\V3/V4/A3/A1/M2/s1 ));
 AND2_X1 \V3/V4/A3/A1/M2/M2/_0_  (.A1(\V3/V4/A3/A1/M2/s1 ),
    .A2(\V3/V4/A3/A1/c1 ),
    .ZN(\V3/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M2/M2/_1_  (.A(\V3/V4/A3/A1/M2/s1 ),
    .B(\V3/V4/A3/A1/c1 ),
    .Z(\V3/v4 [9]));
 OR2_X1 \V3/V4/A3/A1/M2/_0_  (.A1(\V3/V4/A3/A1/M2/c1 ),
    .A2(\V3/V4/A3/A1/M2/c2 ),
    .ZN(\V3/V4/A3/A1/c2 ));
 AND2_X1 \V3/V4/A3/A1/M3/M1/_0_  (.A1(\V3/V4/v4 [2]),
    .A2(\V3/V4/s2 [6]),
    .ZN(\V3/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M3/M1/_1_  (.A(\V3/V4/v4 [2]),
    .B(\V3/V4/s2 [6]),
    .Z(\V3/V4/A3/A1/M3/s1 ));
 AND2_X1 \V3/V4/A3/A1/M3/M2/_0_  (.A1(\V3/V4/A3/A1/M3/s1 ),
    .A2(\V3/V4/A3/A1/c2 ),
    .ZN(\V3/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M3/M2/_1_  (.A(\V3/V4/A3/A1/M3/s1 ),
    .B(\V3/V4/A3/A1/c2 ),
    .Z(\V3/v4 [10]));
 OR2_X1 \V3/V4/A3/A1/M3/_0_  (.A1(\V3/V4/A3/A1/M3/c1 ),
    .A2(\V3/V4/A3/A1/M3/c2 ),
    .ZN(\V3/V4/A3/A1/c3 ));
 AND2_X1 \V3/V4/A3/A1/M4/M1/_0_  (.A1(\V3/V4/v4 [3]),
    .A2(\V3/V4/s2 [7]),
    .ZN(\V3/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M4/M1/_1_  (.A(\V3/V4/v4 [3]),
    .B(\V3/V4/s2 [7]),
    .Z(\V3/V4/A3/A1/M4/s1 ));
 AND2_X1 \V3/V4/A3/A1/M4/M2/_0_  (.A1(\V3/V4/A3/A1/M4/s1 ),
    .A2(\V3/V4/A3/A1/c3 ),
    .ZN(\V3/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M4/M2/_1_  (.A(\V3/V4/A3/A1/M4/s1 ),
    .B(\V3/V4/A3/A1/c3 ),
    .Z(\V3/v4 [11]));
 OR2_X1 \V3/V4/A3/A1/M4/_0_  (.A1(\V3/V4/A3/A1/M4/c1 ),
    .A2(\V3/V4/A3/A1/M4/c2 ),
    .ZN(\V3/V4/A3/c1 ));
 AND2_X1 \V3/V4/A3/A2/M1/M1/_0_  (.A1(\V3/V4/v4 [4]),
    .A2(\V3/V4/c3 ),
    .ZN(\V3/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M1/M1/_1_  (.A(\V3/V4/v4 [4]),
    .B(\V3/V4/c3 ),
    .Z(\V3/V4/A3/A2/M1/s1 ));
 AND2_X1 \V3/V4/A3/A2/M1/M2/_0_  (.A1(\V3/V4/A3/A2/M1/s1 ),
    .A2(\V3/V4/A3/c1 ),
    .ZN(\V3/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M1/M2/_1_  (.A(\V3/V4/A3/A2/M1/s1 ),
    .B(\V3/V4/A3/c1 ),
    .Z(\V3/v4 [12]));
 OR2_X1 \V3/V4/A3/A2/M1/_0_  (.A1(\V3/V4/A3/A2/M1/c1 ),
    .A2(\V3/V4/A3/A2/M1/c2 ),
    .ZN(\V3/V4/A3/A2/c1 ));
 AND2_X1 \V3/V4/A3/A2/M2/M1/_0_  (.A1(\V3/V4/v4 [5]),
    .A2(ground),
    .ZN(\V3/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M2/M1/_1_  (.A(\V3/V4/v4 [5]),
    .B(ground),
    .Z(\V3/V4/A3/A2/M2/s1 ));
 AND2_X1 \V3/V4/A3/A2/M2/M2/_0_  (.A1(\V3/V4/A3/A2/M2/s1 ),
    .A2(\V3/V4/A3/A2/c1 ),
    .ZN(\V3/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M2/M2/_1_  (.A(\V3/V4/A3/A2/M2/s1 ),
    .B(\V3/V4/A3/A2/c1 ),
    .Z(\V3/v4 [13]));
 OR2_X1 \V3/V4/A3/A2/M2/_0_  (.A1(\V3/V4/A3/A2/M2/c1 ),
    .A2(\V3/V4/A3/A2/M2/c2 ),
    .ZN(\V3/V4/A3/A2/c2 ));
 AND2_X1 \V3/V4/A3/A2/M3/M1/_0_  (.A1(\V3/V4/v4 [6]),
    .A2(ground),
    .ZN(\V3/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M3/M1/_1_  (.A(\V3/V4/v4 [6]),
    .B(ground),
    .Z(\V3/V4/A3/A2/M3/s1 ));
 AND2_X1 \V3/V4/A3/A2/M3/M2/_0_  (.A1(\V3/V4/A3/A2/M3/s1 ),
    .A2(\V3/V4/A3/A2/c2 ),
    .ZN(\V3/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M3/M2/_1_  (.A(\V3/V4/A3/A2/M3/s1 ),
    .B(\V3/V4/A3/A2/c2 ),
    .Z(\V3/v4 [14]));
 OR2_X1 \V3/V4/A3/A2/M3/_0_  (.A1(\V3/V4/A3/A2/M3/c1 ),
    .A2(\V3/V4/A3/A2/M3/c2 ),
    .ZN(\V3/V4/A3/A2/c3 ));
 AND2_X1 \V3/V4/A3/A2/M4/M1/_0_  (.A1(\V3/V4/v4 [7]),
    .A2(ground),
    .ZN(\V3/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M4/M1/_1_  (.A(\V3/V4/v4 [7]),
    .B(ground),
    .Z(\V3/V4/A3/A2/M4/s1 ));
 AND2_X1 \V3/V4/A3/A2/M4/M2/_0_  (.A1(\V3/V4/A3/A2/M4/s1 ),
    .A2(\V3/V4/A3/A2/c3 ),
    .ZN(\V3/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M4/M2/_1_  (.A(\V3/V4/A3/A2/M4/s1 ),
    .B(\V3/V4/A3/A2/c3 ),
    .Z(\V3/v4 [15]));
 OR2_X1 \V3/V4/A3/A2/M4/_0_  (.A1(\V3/V4/A3/A2/M4/c1 ),
    .A2(\V3/V4/A3/A2/M4/c2 ),
    .ZN(\V3/V4/overflow ));
 AND2_X1 \V3/V4/V1/A1/M1/M1/_0_  (.A1(\V3/V4/V1/v2 [0]),
    .A2(\V3/V4/V1/v3 [0]),
    .ZN(\V3/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M1/M1/_1_  (.A(\V3/V4/V1/v2 [0]),
    .B(\V3/V4/V1/v3 [0]),
    .Z(\V3/V4/V1/A1/M1/s1 ));
 AND2_X1 \V3/V4/V1/A1/M1/M2/_0_  (.A1(\V3/V4/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M1/M2/_1_  (.A(\V3/V4/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/V1/s1 [0]));
 OR2_X1 \V3/V4/V1/A1/M1/_0_  (.A1(\V3/V4/V1/A1/M1/c1 ),
    .A2(\V3/V4/V1/A1/M1/c2 ),
    .ZN(\V3/V4/V1/A1/c1 ));
 AND2_X1 \V3/V4/V1/A1/M2/M1/_0_  (.A1(\V3/V4/V1/v2 [1]),
    .A2(\V3/V4/V1/v3 [1]),
    .ZN(\V3/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M2/M1/_1_  (.A(\V3/V4/V1/v2 [1]),
    .B(\V3/V4/V1/v3 [1]),
    .Z(\V3/V4/V1/A1/M2/s1 ));
 AND2_X1 \V3/V4/V1/A1/M2/M2/_0_  (.A1(\V3/V4/V1/A1/M2/s1 ),
    .A2(\V3/V4/V1/A1/c1 ),
    .ZN(\V3/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M2/M2/_1_  (.A(\V3/V4/V1/A1/M2/s1 ),
    .B(\V3/V4/V1/A1/c1 ),
    .Z(\V3/V4/V1/s1 [1]));
 OR2_X1 \V3/V4/V1/A1/M2/_0_  (.A1(\V3/V4/V1/A1/M2/c1 ),
    .A2(\V3/V4/V1/A1/M2/c2 ),
    .ZN(\V3/V4/V1/A1/c2 ));
 AND2_X1 \V3/V4/V1/A1/M3/M1/_0_  (.A1(\V3/V4/V1/v2 [2]),
    .A2(\V3/V4/V1/v3 [2]),
    .ZN(\V3/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M3/M1/_1_  (.A(\V3/V4/V1/v2 [2]),
    .B(\V3/V4/V1/v3 [2]),
    .Z(\V3/V4/V1/A1/M3/s1 ));
 AND2_X1 \V3/V4/V1/A1/M3/M2/_0_  (.A1(\V3/V4/V1/A1/M3/s1 ),
    .A2(\V3/V4/V1/A1/c2 ),
    .ZN(\V3/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M3/M2/_1_  (.A(\V3/V4/V1/A1/M3/s1 ),
    .B(\V3/V4/V1/A1/c2 ),
    .Z(\V3/V4/V1/s1 [2]));
 OR2_X1 \V3/V4/V1/A1/M3/_0_  (.A1(\V3/V4/V1/A1/M3/c1 ),
    .A2(\V3/V4/V1/A1/M3/c2 ),
    .ZN(\V3/V4/V1/A1/c3 ));
 AND2_X1 \V3/V4/V1/A1/M4/M1/_0_  (.A1(\V3/V4/V1/v2 [3]),
    .A2(\V3/V4/V1/v3 [3]),
    .ZN(\V3/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M4/M1/_1_  (.A(\V3/V4/V1/v2 [3]),
    .B(\V3/V4/V1/v3 [3]),
    .Z(\V3/V4/V1/A1/M4/s1 ));
 AND2_X1 \V3/V4/V1/A1/M4/M2/_0_  (.A1(\V3/V4/V1/A1/M4/s1 ),
    .A2(\V3/V4/V1/A1/c3 ),
    .ZN(\V3/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M4/M2/_1_  (.A(\V3/V4/V1/A1/M4/s1 ),
    .B(\V3/V4/V1/A1/c3 ),
    .Z(\V3/V4/V1/s1 [3]));
 OR2_X1 \V3/V4/V1/A1/M4/_0_  (.A1(\V3/V4/V1/A1/M4/c1 ),
    .A2(\V3/V4/V1/A1/M4/c2 ),
    .ZN(\V3/V4/V1/c1 ));
 AND2_X1 \V3/V4/V1/A2/M1/M1/_0_  (.A1(\V3/V4/V1/s1 [0]),
    .A2(\V3/V4/V1/v1 [2]),
    .ZN(\V3/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M1/M1/_1_  (.A(\V3/V4/V1/s1 [0]),
    .B(\V3/V4/V1/v1 [2]),
    .Z(\V3/V4/V1/A2/M1/s1 ));
 AND2_X1 \V3/V4/V1/A2/M1/M2/_0_  (.A1(\V3/V4/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M1/M2/_1_  (.A(\V3/V4/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/v4 [2]));
 OR2_X1 \V3/V4/V1/A2/M1/_0_  (.A1(\V3/V4/V1/A2/M1/c1 ),
    .A2(\V3/V4/V1/A2/M1/c2 ),
    .ZN(\V3/V4/V1/A2/c1 ));
 AND2_X1 \V3/V4/V1/A2/M2/M1/_0_  (.A1(\V3/V4/V1/s1 [1]),
    .A2(\V3/V4/V1/v1 [3]),
    .ZN(\V3/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M2/M1/_1_  (.A(\V3/V4/V1/s1 [1]),
    .B(\V3/V4/V1/v1 [3]),
    .Z(\V3/V4/V1/A2/M2/s1 ));
 AND2_X1 \V3/V4/V1/A2/M2/M2/_0_  (.A1(\V3/V4/V1/A2/M2/s1 ),
    .A2(\V3/V4/V1/A2/c1 ),
    .ZN(\V3/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M2/M2/_1_  (.A(\V3/V4/V1/A2/M2/s1 ),
    .B(\V3/V4/V1/A2/c1 ),
    .Z(\V3/v4 [3]));
 OR2_X1 \V3/V4/V1/A2/M2/_0_  (.A1(\V3/V4/V1/A2/M2/c1 ),
    .A2(\V3/V4/V1/A2/M2/c2 ),
    .ZN(\V3/V4/V1/A2/c2 ));
 AND2_X1 \V3/V4/V1/A2/M3/M1/_0_  (.A1(\V3/V4/V1/s1 [2]),
    .A2(ground),
    .ZN(\V3/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M3/M1/_1_  (.A(\V3/V4/V1/s1 [2]),
    .B(ground),
    .Z(\V3/V4/V1/A2/M3/s1 ));
 AND2_X1 \V3/V4/V1/A2/M3/M2/_0_  (.A1(\V3/V4/V1/A2/M3/s1 ),
    .A2(\V3/V4/V1/A2/c2 ),
    .ZN(\V3/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M3/M2/_1_  (.A(\V3/V4/V1/A2/M3/s1 ),
    .B(\V3/V4/V1/A2/c2 ),
    .Z(\V3/V4/V1/s2 [2]));
 OR2_X1 \V3/V4/V1/A2/M3/_0_  (.A1(\V3/V4/V1/A2/M3/c1 ),
    .A2(\V3/V4/V1/A2/M3/c2 ),
    .ZN(\V3/V4/V1/A2/c3 ));
 AND2_X1 \V3/V4/V1/A2/M4/M1/_0_  (.A1(\V3/V4/V1/s1 [3]),
    .A2(ground),
    .ZN(\V3/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M4/M1/_1_  (.A(\V3/V4/V1/s1 [3]),
    .B(ground),
    .Z(\V3/V4/V1/A2/M4/s1 ));
 AND2_X1 \V3/V4/V1/A2/M4/M2/_0_  (.A1(\V3/V4/V1/A2/M4/s1 ),
    .A2(\V3/V4/V1/A2/c3 ),
    .ZN(\V3/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M4/M2/_1_  (.A(\V3/V4/V1/A2/M4/s1 ),
    .B(\V3/V4/V1/A2/c3 ),
    .Z(\V3/V4/V1/s2 [3]));
 OR2_X1 \V3/V4/V1/A2/M4/_0_  (.A1(\V3/V4/V1/A2/M4/c1 ),
    .A2(\V3/V4/V1/A2/M4/c2 ),
    .ZN(\V3/V4/V1/c2 ));
 AND2_X1 \V3/V4/V1/A3/M1/M1/_0_  (.A1(\V3/V4/V1/v4 [0]),
    .A2(\V3/V4/V1/s2 [2]),
    .ZN(\V3/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M1/M1/_1_  (.A(\V3/V4/V1/v4 [0]),
    .B(\V3/V4/V1/s2 [2]),
    .Z(\V3/V4/V1/A3/M1/s1 ));
 AND2_X1 \V3/V4/V1/A3/M1/M2/_0_  (.A1(\V3/V4/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M1/M2/_1_  (.A(\V3/V4/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v1 [4]));
 OR2_X1 \V3/V4/V1/A3/M1/_0_  (.A1(\V3/V4/V1/A3/M1/c1 ),
    .A2(\V3/V4/V1/A3/M1/c2 ),
    .ZN(\V3/V4/V1/A3/c1 ));
 AND2_X1 \V3/V4/V1/A3/M2/M1/_0_  (.A1(\V3/V4/V1/v4 [1]),
    .A2(\V3/V4/V1/s2 [3]),
    .ZN(\V3/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M2/M1/_1_  (.A(\V3/V4/V1/v4 [1]),
    .B(\V3/V4/V1/s2 [3]),
    .Z(\V3/V4/V1/A3/M2/s1 ));
 AND2_X1 \V3/V4/V1/A3/M2/M2/_0_  (.A1(\V3/V4/V1/A3/M2/s1 ),
    .A2(\V3/V4/V1/A3/c1 ),
    .ZN(\V3/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M2/M2/_1_  (.A(\V3/V4/V1/A3/M2/s1 ),
    .B(\V3/V4/V1/A3/c1 ),
    .Z(\V3/V4/v1 [5]));
 OR2_X1 \V3/V4/V1/A3/M2/_0_  (.A1(\V3/V4/V1/A3/M2/c1 ),
    .A2(\V3/V4/V1/A3/M2/c2 ),
    .ZN(\V3/V4/V1/A3/c2 ));
 AND2_X1 \V3/V4/V1/A3/M3/M1/_0_  (.A1(\V3/V4/V1/v4 [2]),
    .A2(\V3/V4/V1/c3 ),
    .ZN(\V3/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M3/M1/_1_  (.A(\V3/V4/V1/v4 [2]),
    .B(\V3/V4/V1/c3 ),
    .Z(\V3/V4/V1/A3/M3/s1 ));
 AND2_X1 \V3/V4/V1/A3/M3/M2/_0_  (.A1(\V3/V4/V1/A3/M3/s1 ),
    .A2(\V3/V4/V1/A3/c2 ),
    .ZN(\V3/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M3/M2/_1_  (.A(\V3/V4/V1/A3/M3/s1 ),
    .B(\V3/V4/V1/A3/c2 ),
    .Z(\V3/V4/v1 [6]));
 OR2_X1 \V3/V4/V1/A3/M3/_0_  (.A1(\V3/V4/V1/A3/M3/c1 ),
    .A2(\V3/V4/V1/A3/M3/c2 ),
    .ZN(\V3/V4/V1/A3/c3 ));
 AND2_X1 \V3/V4/V1/A3/M4/M1/_0_  (.A1(\V3/V4/V1/v4 [3]),
    .A2(ground),
    .ZN(\V3/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M4/M1/_1_  (.A(\V3/V4/V1/v4 [3]),
    .B(ground),
    .Z(\V3/V4/V1/A3/M4/s1 ));
 AND2_X1 \V3/V4/V1/A3/M4/M2/_0_  (.A1(\V3/V4/V1/A3/M4/s1 ),
    .A2(\V3/V4/V1/A3/c3 ),
    .ZN(\V3/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M4/M2/_1_  (.A(\V3/V4/V1/A3/M4/s1 ),
    .B(\V3/V4/V1/A3/c3 ),
    .Z(\V3/V4/v1 [7]));
 OR2_X1 \V3/V4/V1/A3/M4/_0_  (.A1(\V3/V4/V1/A3/M4/c1 ),
    .A2(\V3/V4/V1/A3/M4/c2 ),
    .ZN(\V3/V4/V1/overflow ));
 AND2_X1 \V3/V4/V1/V1/HA1/_0_  (.A1(\V3/V4/V1/V1/w2 ),
    .A2(\V3/V4/V1/V1/w1 ),
    .ZN(\V3/V4/V1/V1/w4 ));
 XOR2_X2 \V3/V4/V1/V1/HA1/_1_  (.A(\V3/V4/V1/V1/w2 ),
    .B(\V3/V4/V1/V1/w1 ),
    .Z(\V3/v4 [1]));
 AND2_X1 \V3/V4/V1/V1/HA2/_0_  (.A1(\V3/V4/V1/V1/w4 ),
    .A2(\V3/V4/V1/V1/w3 ),
    .ZN(\V3/V4/V1/v1 [3]));
 XOR2_X2 \V3/V4/V1/V1/HA2/_1_  (.A(\V3/V4/V1/V1/w4 ),
    .B(\V3/V4/V1/V1/w3 ),
    .Z(\V3/V4/V1/v1 [2]));
 AND2_X1 \V3/V4/V1/V1/_0_  (.A1(A[8]),
    .A2(B[24]),
    .ZN(\V3/v4 [0]));
 AND2_X1 \V3/V4/V1/V1/_1_  (.A1(A[8]),
    .A2(B[25]),
    .ZN(\V3/V4/V1/V1/w1 ));
 AND2_X1 \V3/V4/V1/V1/_2_  (.A1(B[24]),
    .A2(A[9]),
    .ZN(\V3/V4/V1/V1/w2 ));
 AND2_X1 \V3/V4/V1/V1/_3_  (.A1(B[25]),
    .A2(A[9]),
    .ZN(\V3/V4/V1/V1/w3 ));
 AND2_X1 \V3/V4/V1/V2/HA1/_0_  (.A1(\V3/V4/V1/V2/w2 ),
    .A2(\V3/V4/V1/V2/w1 ),
    .ZN(\V3/V4/V1/V2/w4 ));
 XOR2_X2 \V3/V4/V1/V2/HA1/_1_  (.A(\V3/V4/V1/V2/w2 ),
    .B(\V3/V4/V1/V2/w1 ),
    .Z(\V3/V4/V1/v2 [1]));
 AND2_X1 \V3/V4/V1/V2/HA2/_0_  (.A1(\V3/V4/V1/V2/w4 ),
    .A2(\V3/V4/V1/V2/w3 ),
    .ZN(\V3/V4/V1/v2 [3]));
 XOR2_X2 \V3/V4/V1/V2/HA2/_1_  (.A(\V3/V4/V1/V2/w4 ),
    .B(\V3/V4/V1/V2/w3 ),
    .Z(\V3/V4/V1/v2 [2]));
 AND2_X1 \V3/V4/V1/V2/_0_  (.A1(A[10]),
    .A2(B[24]),
    .ZN(\V3/V4/V1/v2 [0]));
 AND2_X1 \V3/V4/V1/V2/_1_  (.A1(A[10]),
    .A2(B[25]),
    .ZN(\V3/V4/V1/V2/w1 ));
 AND2_X1 \V3/V4/V1/V2/_2_  (.A1(B[24]),
    .A2(A[11]),
    .ZN(\V3/V4/V1/V2/w2 ));
 AND2_X1 \V3/V4/V1/V2/_3_  (.A1(B[25]),
    .A2(A[11]),
    .ZN(\V3/V4/V1/V2/w3 ));
 AND2_X1 \V3/V4/V1/V3/HA1/_0_  (.A1(\V3/V4/V1/V3/w2 ),
    .A2(\V3/V4/V1/V3/w1 ),
    .ZN(\V3/V4/V1/V3/w4 ));
 XOR2_X2 \V3/V4/V1/V3/HA1/_1_  (.A(\V3/V4/V1/V3/w2 ),
    .B(\V3/V4/V1/V3/w1 ),
    .Z(\V3/V4/V1/v3 [1]));
 AND2_X1 \V3/V4/V1/V3/HA2/_0_  (.A1(\V3/V4/V1/V3/w4 ),
    .A2(\V3/V4/V1/V3/w3 ),
    .ZN(\V3/V4/V1/v3 [3]));
 XOR2_X2 \V3/V4/V1/V3/HA2/_1_  (.A(\V3/V4/V1/V3/w4 ),
    .B(\V3/V4/V1/V3/w3 ),
    .Z(\V3/V4/V1/v3 [2]));
 AND2_X1 \V3/V4/V1/V3/_0_  (.A1(A[8]),
    .A2(B[26]),
    .ZN(\V3/V4/V1/v3 [0]));
 AND2_X1 \V3/V4/V1/V3/_1_  (.A1(A[8]),
    .A2(B[27]),
    .ZN(\V3/V4/V1/V3/w1 ));
 AND2_X1 \V3/V4/V1/V3/_2_  (.A1(B[26]),
    .A2(A[9]),
    .ZN(\V3/V4/V1/V3/w2 ));
 AND2_X1 \V3/V4/V1/V3/_3_  (.A1(B[27]),
    .A2(A[9]),
    .ZN(\V3/V4/V1/V3/w3 ));
 AND2_X1 \V3/V4/V1/V4/HA1/_0_  (.A1(\V3/V4/V1/V4/w2 ),
    .A2(\V3/V4/V1/V4/w1 ),
    .ZN(\V3/V4/V1/V4/w4 ));
 XOR2_X2 \V3/V4/V1/V4/HA1/_1_  (.A(\V3/V4/V1/V4/w2 ),
    .B(\V3/V4/V1/V4/w1 ),
    .Z(\V3/V4/V1/v4 [1]));
 AND2_X1 \V3/V4/V1/V4/HA2/_0_  (.A1(\V3/V4/V1/V4/w4 ),
    .A2(\V3/V4/V1/V4/w3 ),
    .ZN(\V3/V4/V1/v4 [3]));
 XOR2_X2 \V3/V4/V1/V4/HA2/_1_  (.A(\V3/V4/V1/V4/w4 ),
    .B(\V3/V4/V1/V4/w3 ),
    .Z(\V3/V4/V1/v4 [2]));
 AND2_X1 \V3/V4/V1/V4/_0_  (.A1(A[10]),
    .A2(B[26]),
    .ZN(\V3/V4/V1/v4 [0]));
 AND2_X1 \V3/V4/V1/V4/_1_  (.A1(A[10]),
    .A2(B[27]),
    .ZN(\V3/V4/V1/V4/w1 ));
 AND2_X1 \V3/V4/V1/V4/_2_  (.A1(B[26]),
    .A2(A[11]),
    .ZN(\V3/V4/V1/V4/w2 ));
 AND2_X1 \V3/V4/V1/V4/_3_  (.A1(B[27]),
    .A2(A[11]),
    .ZN(\V3/V4/V1/V4/w3 ));
 OR2_X1 \V3/V4/V1/_0_  (.A1(\V3/V4/V1/c1 ),
    .A2(\V3/V4/V1/c2 ),
    .ZN(\V3/V4/V1/c3 ));
 AND2_X1 \V3/V4/V2/A1/M1/M1/_0_  (.A1(\V3/V4/V2/v2 [0]),
    .A2(\V3/V4/V2/v3 [0]),
    .ZN(\V3/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M1/M1/_1_  (.A(\V3/V4/V2/v2 [0]),
    .B(\V3/V4/V2/v3 [0]),
    .Z(\V3/V4/V2/A1/M1/s1 ));
 AND2_X1 \V3/V4/V2/A1/M1/M2/_0_  (.A1(\V3/V4/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M1/M2/_1_  (.A(\V3/V4/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/V2/s1 [0]));
 OR2_X1 \V3/V4/V2/A1/M1/_0_  (.A1(\V3/V4/V2/A1/M1/c1 ),
    .A2(\V3/V4/V2/A1/M1/c2 ),
    .ZN(\V3/V4/V2/A1/c1 ));
 AND2_X1 \V3/V4/V2/A1/M2/M1/_0_  (.A1(\V3/V4/V2/v2 [1]),
    .A2(\V3/V4/V2/v3 [1]),
    .ZN(\V3/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M2/M1/_1_  (.A(\V3/V4/V2/v2 [1]),
    .B(\V3/V4/V2/v3 [1]),
    .Z(\V3/V4/V2/A1/M2/s1 ));
 AND2_X1 \V3/V4/V2/A1/M2/M2/_0_  (.A1(\V3/V4/V2/A1/M2/s1 ),
    .A2(\V3/V4/V2/A1/c1 ),
    .ZN(\V3/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M2/M2/_1_  (.A(\V3/V4/V2/A1/M2/s1 ),
    .B(\V3/V4/V2/A1/c1 ),
    .Z(\V3/V4/V2/s1 [1]));
 OR2_X1 \V3/V4/V2/A1/M2/_0_  (.A1(\V3/V4/V2/A1/M2/c1 ),
    .A2(\V3/V4/V2/A1/M2/c2 ),
    .ZN(\V3/V4/V2/A1/c2 ));
 AND2_X1 \V3/V4/V2/A1/M3/M1/_0_  (.A1(\V3/V4/V2/v2 [2]),
    .A2(\V3/V4/V2/v3 [2]),
    .ZN(\V3/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M3/M1/_1_  (.A(\V3/V4/V2/v2 [2]),
    .B(\V3/V4/V2/v3 [2]),
    .Z(\V3/V4/V2/A1/M3/s1 ));
 AND2_X1 \V3/V4/V2/A1/M3/M2/_0_  (.A1(\V3/V4/V2/A1/M3/s1 ),
    .A2(\V3/V4/V2/A1/c2 ),
    .ZN(\V3/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M3/M2/_1_  (.A(\V3/V4/V2/A1/M3/s1 ),
    .B(\V3/V4/V2/A1/c2 ),
    .Z(\V3/V4/V2/s1 [2]));
 OR2_X1 \V3/V4/V2/A1/M3/_0_  (.A1(\V3/V4/V2/A1/M3/c1 ),
    .A2(\V3/V4/V2/A1/M3/c2 ),
    .ZN(\V3/V4/V2/A1/c3 ));
 AND2_X1 \V3/V4/V2/A1/M4/M1/_0_  (.A1(\V3/V4/V2/v2 [3]),
    .A2(\V3/V4/V2/v3 [3]),
    .ZN(\V3/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M4/M1/_1_  (.A(\V3/V4/V2/v2 [3]),
    .B(\V3/V4/V2/v3 [3]),
    .Z(\V3/V4/V2/A1/M4/s1 ));
 AND2_X1 \V3/V4/V2/A1/M4/M2/_0_  (.A1(\V3/V4/V2/A1/M4/s1 ),
    .A2(\V3/V4/V2/A1/c3 ),
    .ZN(\V3/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M4/M2/_1_  (.A(\V3/V4/V2/A1/M4/s1 ),
    .B(\V3/V4/V2/A1/c3 ),
    .Z(\V3/V4/V2/s1 [3]));
 OR2_X1 \V3/V4/V2/A1/M4/_0_  (.A1(\V3/V4/V2/A1/M4/c1 ),
    .A2(\V3/V4/V2/A1/M4/c2 ),
    .ZN(\V3/V4/V2/c1 ));
 AND2_X1 \V3/V4/V2/A2/M1/M1/_0_  (.A1(\V3/V4/V2/s1 [0]),
    .A2(\V3/V4/V2/v1 [2]),
    .ZN(\V3/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M1/M1/_1_  (.A(\V3/V4/V2/s1 [0]),
    .B(\V3/V4/V2/v1 [2]),
    .Z(\V3/V4/V2/A2/M1/s1 ));
 AND2_X1 \V3/V4/V2/A2/M1/M2/_0_  (.A1(\V3/V4/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M1/M2/_1_  (.A(\V3/V4/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v2 [2]));
 OR2_X1 \V3/V4/V2/A2/M1/_0_  (.A1(\V3/V4/V2/A2/M1/c1 ),
    .A2(\V3/V4/V2/A2/M1/c2 ),
    .ZN(\V3/V4/V2/A2/c1 ));
 AND2_X1 \V3/V4/V2/A2/M2/M1/_0_  (.A1(\V3/V4/V2/s1 [1]),
    .A2(\V3/V4/V2/v1 [3]),
    .ZN(\V3/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M2/M1/_1_  (.A(\V3/V4/V2/s1 [1]),
    .B(\V3/V4/V2/v1 [3]),
    .Z(\V3/V4/V2/A2/M2/s1 ));
 AND2_X1 \V3/V4/V2/A2/M2/M2/_0_  (.A1(\V3/V4/V2/A2/M2/s1 ),
    .A2(\V3/V4/V2/A2/c1 ),
    .ZN(\V3/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M2/M2/_1_  (.A(\V3/V4/V2/A2/M2/s1 ),
    .B(\V3/V4/V2/A2/c1 ),
    .Z(\V3/V4/v2 [3]));
 OR2_X1 \V3/V4/V2/A2/M2/_0_  (.A1(\V3/V4/V2/A2/M2/c1 ),
    .A2(\V3/V4/V2/A2/M2/c2 ),
    .ZN(\V3/V4/V2/A2/c2 ));
 AND2_X1 \V3/V4/V2/A2/M3/M1/_0_  (.A1(\V3/V4/V2/s1 [2]),
    .A2(ground),
    .ZN(\V3/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M3/M1/_1_  (.A(\V3/V4/V2/s1 [2]),
    .B(ground),
    .Z(\V3/V4/V2/A2/M3/s1 ));
 AND2_X1 \V3/V4/V2/A2/M3/M2/_0_  (.A1(\V3/V4/V2/A2/M3/s1 ),
    .A2(\V3/V4/V2/A2/c2 ),
    .ZN(\V3/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M3/M2/_1_  (.A(\V3/V4/V2/A2/M3/s1 ),
    .B(\V3/V4/V2/A2/c2 ),
    .Z(\V3/V4/V2/s2 [2]));
 OR2_X1 \V3/V4/V2/A2/M3/_0_  (.A1(\V3/V4/V2/A2/M3/c1 ),
    .A2(\V3/V4/V2/A2/M3/c2 ),
    .ZN(\V3/V4/V2/A2/c3 ));
 AND2_X1 \V3/V4/V2/A2/M4/M1/_0_  (.A1(\V3/V4/V2/s1 [3]),
    .A2(ground),
    .ZN(\V3/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M4/M1/_1_  (.A(\V3/V4/V2/s1 [3]),
    .B(ground),
    .Z(\V3/V4/V2/A2/M4/s1 ));
 AND2_X1 \V3/V4/V2/A2/M4/M2/_0_  (.A1(\V3/V4/V2/A2/M4/s1 ),
    .A2(\V3/V4/V2/A2/c3 ),
    .ZN(\V3/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M4/M2/_1_  (.A(\V3/V4/V2/A2/M4/s1 ),
    .B(\V3/V4/V2/A2/c3 ),
    .Z(\V3/V4/V2/s2 [3]));
 OR2_X1 \V3/V4/V2/A2/M4/_0_  (.A1(\V3/V4/V2/A2/M4/c1 ),
    .A2(\V3/V4/V2/A2/M4/c2 ),
    .ZN(\V3/V4/V2/c2 ));
 AND2_X1 \V3/V4/V2/A3/M1/M1/_0_  (.A1(\V3/V4/V2/v4 [0]),
    .A2(\V3/V4/V2/s2 [2]),
    .ZN(\V3/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M1/M1/_1_  (.A(\V3/V4/V2/v4 [0]),
    .B(\V3/V4/V2/s2 [2]),
    .Z(\V3/V4/V2/A3/M1/s1 ));
 AND2_X1 \V3/V4/V2/A3/M1/M2/_0_  (.A1(\V3/V4/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M1/M2/_1_  (.A(\V3/V4/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v2 [4]));
 OR2_X1 \V3/V4/V2/A3/M1/_0_  (.A1(\V3/V4/V2/A3/M1/c1 ),
    .A2(\V3/V4/V2/A3/M1/c2 ),
    .ZN(\V3/V4/V2/A3/c1 ));
 AND2_X1 \V3/V4/V2/A3/M2/M1/_0_  (.A1(\V3/V4/V2/v4 [1]),
    .A2(\V3/V4/V2/s2 [3]),
    .ZN(\V3/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M2/M1/_1_  (.A(\V3/V4/V2/v4 [1]),
    .B(\V3/V4/V2/s2 [3]),
    .Z(\V3/V4/V2/A3/M2/s1 ));
 AND2_X1 \V3/V4/V2/A3/M2/M2/_0_  (.A1(\V3/V4/V2/A3/M2/s1 ),
    .A2(\V3/V4/V2/A3/c1 ),
    .ZN(\V3/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M2/M2/_1_  (.A(\V3/V4/V2/A3/M2/s1 ),
    .B(\V3/V4/V2/A3/c1 ),
    .Z(\V3/V4/v2 [5]));
 OR2_X1 \V3/V4/V2/A3/M2/_0_  (.A1(\V3/V4/V2/A3/M2/c1 ),
    .A2(\V3/V4/V2/A3/M2/c2 ),
    .ZN(\V3/V4/V2/A3/c2 ));
 AND2_X1 \V3/V4/V2/A3/M3/M1/_0_  (.A1(\V3/V4/V2/v4 [2]),
    .A2(\V3/V4/V2/c3 ),
    .ZN(\V3/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M3/M1/_1_  (.A(\V3/V4/V2/v4 [2]),
    .B(\V3/V4/V2/c3 ),
    .Z(\V3/V4/V2/A3/M3/s1 ));
 AND2_X1 \V3/V4/V2/A3/M3/M2/_0_  (.A1(\V3/V4/V2/A3/M3/s1 ),
    .A2(\V3/V4/V2/A3/c2 ),
    .ZN(\V3/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M3/M2/_1_  (.A(\V3/V4/V2/A3/M3/s1 ),
    .B(\V3/V4/V2/A3/c2 ),
    .Z(\V3/V4/v2 [6]));
 OR2_X1 \V3/V4/V2/A3/M3/_0_  (.A1(\V3/V4/V2/A3/M3/c1 ),
    .A2(\V3/V4/V2/A3/M3/c2 ),
    .ZN(\V3/V4/V2/A3/c3 ));
 AND2_X1 \V3/V4/V2/A3/M4/M1/_0_  (.A1(\V3/V4/V2/v4 [3]),
    .A2(ground),
    .ZN(\V3/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M4/M1/_1_  (.A(\V3/V4/V2/v4 [3]),
    .B(ground),
    .Z(\V3/V4/V2/A3/M4/s1 ));
 AND2_X1 \V3/V4/V2/A3/M4/M2/_0_  (.A1(\V3/V4/V2/A3/M4/s1 ),
    .A2(\V3/V4/V2/A3/c3 ),
    .ZN(\V3/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M4/M2/_1_  (.A(\V3/V4/V2/A3/M4/s1 ),
    .B(\V3/V4/V2/A3/c3 ),
    .Z(\V3/V4/v2 [7]));
 OR2_X1 \V3/V4/V2/A3/M4/_0_  (.A1(\V3/V4/V2/A3/M4/c1 ),
    .A2(\V3/V4/V2/A3/M4/c2 ),
    .ZN(\V3/V4/V2/overflow ));
 AND2_X1 \V3/V4/V2/V1/HA1/_0_  (.A1(\V3/V4/V2/V1/w2 ),
    .A2(\V3/V4/V2/V1/w1 ),
    .ZN(\V3/V4/V2/V1/w4 ));
 XOR2_X2 \V3/V4/V2/V1/HA1/_1_  (.A(\V3/V4/V2/V1/w2 ),
    .B(\V3/V4/V2/V1/w1 ),
    .Z(\V3/V4/v2 [1]));
 AND2_X1 \V3/V4/V2/V1/HA2/_0_  (.A1(\V3/V4/V2/V1/w4 ),
    .A2(\V3/V4/V2/V1/w3 ),
    .ZN(\V3/V4/V2/v1 [3]));
 XOR2_X2 \V3/V4/V2/V1/HA2/_1_  (.A(\V3/V4/V2/V1/w4 ),
    .B(\V3/V4/V2/V1/w3 ),
    .Z(\V3/V4/V2/v1 [2]));
 AND2_X1 \V3/V4/V2/V1/_0_  (.A1(A[12]),
    .A2(B[24]),
    .ZN(\V3/V4/v2 [0]));
 AND2_X1 \V3/V4/V2/V1/_1_  (.A1(A[12]),
    .A2(B[25]),
    .ZN(\V3/V4/V2/V1/w1 ));
 AND2_X1 \V3/V4/V2/V1/_2_  (.A1(B[24]),
    .A2(A[13]),
    .ZN(\V3/V4/V2/V1/w2 ));
 AND2_X1 \V3/V4/V2/V1/_3_  (.A1(B[25]),
    .A2(A[13]),
    .ZN(\V3/V4/V2/V1/w3 ));
 AND2_X1 \V3/V4/V2/V2/HA1/_0_  (.A1(\V3/V4/V2/V2/w2 ),
    .A2(\V3/V4/V2/V2/w1 ),
    .ZN(\V3/V4/V2/V2/w4 ));
 XOR2_X2 \V3/V4/V2/V2/HA1/_1_  (.A(\V3/V4/V2/V2/w2 ),
    .B(\V3/V4/V2/V2/w1 ),
    .Z(\V3/V4/V2/v2 [1]));
 AND2_X1 \V3/V4/V2/V2/HA2/_0_  (.A1(\V3/V4/V2/V2/w4 ),
    .A2(\V3/V4/V2/V2/w3 ),
    .ZN(\V3/V4/V2/v2 [3]));
 XOR2_X2 \V3/V4/V2/V2/HA2/_1_  (.A(\V3/V4/V2/V2/w4 ),
    .B(\V3/V4/V2/V2/w3 ),
    .Z(\V3/V4/V2/v2 [2]));
 AND2_X1 \V3/V4/V2/V2/_0_  (.A1(A[14]),
    .A2(B[24]),
    .ZN(\V3/V4/V2/v2 [0]));
 AND2_X1 \V3/V4/V2/V2/_1_  (.A1(A[14]),
    .A2(B[25]),
    .ZN(\V3/V4/V2/V2/w1 ));
 AND2_X1 \V3/V4/V2/V2/_2_  (.A1(B[24]),
    .A2(A[15]),
    .ZN(\V3/V4/V2/V2/w2 ));
 AND2_X1 \V3/V4/V2/V2/_3_  (.A1(B[25]),
    .A2(A[15]),
    .ZN(\V3/V4/V2/V2/w3 ));
 AND2_X1 \V3/V4/V2/V3/HA1/_0_  (.A1(\V3/V4/V2/V3/w2 ),
    .A2(\V3/V4/V2/V3/w1 ),
    .ZN(\V3/V4/V2/V3/w4 ));
 XOR2_X2 \V3/V4/V2/V3/HA1/_1_  (.A(\V3/V4/V2/V3/w2 ),
    .B(\V3/V4/V2/V3/w1 ),
    .Z(\V3/V4/V2/v3 [1]));
 AND2_X1 \V3/V4/V2/V3/HA2/_0_  (.A1(\V3/V4/V2/V3/w4 ),
    .A2(\V3/V4/V2/V3/w3 ),
    .ZN(\V3/V4/V2/v3 [3]));
 XOR2_X2 \V3/V4/V2/V3/HA2/_1_  (.A(\V3/V4/V2/V3/w4 ),
    .B(\V3/V4/V2/V3/w3 ),
    .Z(\V3/V4/V2/v3 [2]));
 AND2_X1 \V3/V4/V2/V3/_0_  (.A1(A[12]),
    .A2(B[26]),
    .ZN(\V3/V4/V2/v3 [0]));
 AND2_X1 \V3/V4/V2/V3/_1_  (.A1(A[12]),
    .A2(B[27]),
    .ZN(\V3/V4/V2/V3/w1 ));
 AND2_X1 \V3/V4/V2/V3/_2_  (.A1(B[26]),
    .A2(A[13]),
    .ZN(\V3/V4/V2/V3/w2 ));
 AND2_X1 \V3/V4/V2/V3/_3_  (.A1(B[27]),
    .A2(A[13]),
    .ZN(\V3/V4/V2/V3/w3 ));
 AND2_X1 \V3/V4/V2/V4/HA1/_0_  (.A1(\V3/V4/V2/V4/w2 ),
    .A2(\V3/V4/V2/V4/w1 ),
    .ZN(\V3/V4/V2/V4/w4 ));
 XOR2_X2 \V3/V4/V2/V4/HA1/_1_  (.A(\V3/V4/V2/V4/w2 ),
    .B(\V3/V4/V2/V4/w1 ),
    .Z(\V3/V4/V2/v4 [1]));
 AND2_X1 \V3/V4/V2/V4/HA2/_0_  (.A1(\V3/V4/V2/V4/w4 ),
    .A2(\V3/V4/V2/V4/w3 ),
    .ZN(\V3/V4/V2/v4 [3]));
 XOR2_X2 \V3/V4/V2/V4/HA2/_1_  (.A(\V3/V4/V2/V4/w4 ),
    .B(\V3/V4/V2/V4/w3 ),
    .Z(\V3/V4/V2/v4 [2]));
 AND2_X1 \V3/V4/V2/V4/_0_  (.A1(A[14]),
    .A2(B[26]),
    .ZN(\V3/V4/V2/v4 [0]));
 AND2_X1 \V3/V4/V2/V4/_1_  (.A1(A[14]),
    .A2(B[27]),
    .ZN(\V3/V4/V2/V4/w1 ));
 AND2_X1 \V3/V4/V2/V4/_2_  (.A1(B[26]),
    .A2(A[15]),
    .ZN(\V3/V4/V2/V4/w2 ));
 AND2_X1 \V3/V4/V2/V4/_3_  (.A1(B[27]),
    .A2(A[15]),
    .ZN(\V3/V4/V2/V4/w3 ));
 OR2_X1 \V3/V4/V2/_0_  (.A1(\V3/V4/V2/c1 ),
    .A2(\V3/V4/V2/c2 ),
    .ZN(\V3/V4/V2/c3 ));
 AND2_X1 \V3/V4/V3/A1/M1/M1/_0_  (.A1(\V3/V4/V3/v2 [0]),
    .A2(\V3/V4/V3/v3 [0]),
    .ZN(\V3/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M1/M1/_1_  (.A(\V3/V4/V3/v2 [0]),
    .B(\V3/V4/V3/v3 [0]),
    .Z(\V3/V4/V3/A1/M1/s1 ));
 AND2_X1 \V3/V4/V3/A1/M1/M2/_0_  (.A1(\V3/V4/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M1/M2/_1_  (.A(\V3/V4/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/V3/s1 [0]));
 OR2_X1 \V3/V4/V3/A1/M1/_0_  (.A1(\V3/V4/V3/A1/M1/c1 ),
    .A2(\V3/V4/V3/A1/M1/c2 ),
    .ZN(\V3/V4/V3/A1/c1 ));
 AND2_X1 \V3/V4/V3/A1/M2/M1/_0_  (.A1(\V3/V4/V3/v2 [1]),
    .A2(\V3/V4/V3/v3 [1]),
    .ZN(\V3/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M2/M1/_1_  (.A(\V3/V4/V3/v2 [1]),
    .B(\V3/V4/V3/v3 [1]),
    .Z(\V3/V4/V3/A1/M2/s1 ));
 AND2_X1 \V3/V4/V3/A1/M2/M2/_0_  (.A1(\V3/V4/V3/A1/M2/s1 ),
    .A2(\V3/V4/V3/A1/c1 ),
    .ZN(\V3/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M2/M2/_1_  (.A(\V3/V4/V3/A1/M2/s1 ),
    .B(\V3/V4/V3/A1/c1 ),
    .Z(\V3/V4/V3/s1 [1]));
 OR2_X1 \V3/V4/V3/A1/M2/_0_  (.A1(\V3/V4/V3/A1/M2/c1 ),
    .A2(\V3/V4/V3/A1/M2/c2 ),
    .ZN(\V3/V4/V3/A1/c2 ));
 AND2_X1 \V3/V4/V3/A1/M3/M1/_0_  (.A1(\V3/V4/V3/v2 [2]),
    .A2(\V3/V4/V3/v3 [2]),
    .ZN(\V3/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M3/M1/_1_  (.A(\V3/V4/V3/v2 [2]),
    .B(\V3/V4/V3/v3 [2]),
    .Z(\V3/V4/V3/A1/M3/s1 ));
 AND2_X1 \V3/V4/V3/A1/M3/M2/_0_  (.A1(\V3/V4/V3/A1/M3/s1 ),
    .A2(\V3/V4/V3/A1/c2 ),
    .ZN(\V3/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M3/M2/_1_  (.A(\V3/V4/V3/A1/M3/s1 ),
    .B(\V3/V4/V3/A1/c2 ),
    .Z(\V3/V4/V3/s1 [2]));
 OR2_X1 \V3/V4/V3/A1/M3/_0_  (.A1(\V3/V4/V3/A1/M3/c1 ),
    .A2(\V3/V4/V3/A1/M3/c2 ),
    .ZN(\V3/V4/V3/A1/c3 ));
 AND2_X1 \V3/V4/V3/A1/M4/M1/_0_  (.A1(\V3/V4/V3/v2 [3]),
    .A2(\V3/V4/V3/v3 [3]),
    .ZN(\V3/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M4/M1/_1_  (.A(\V3/V4/V3/v2 [3]),
    .B(\V3/V4/V3/v3 [3]),
    .Z(\V3/V4/V3/A1/M4/s1 ));
 AND2_X1 \V3/V4/V3/A1/M4/M2/_0_  (.A1(\V3/V4/V3/A1/M4/s1 ),
    .A2(\V3/V4/V3/A1/c3 ),
    .ZN(\V3/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M4/M2/_1_  (.A(\V3/V4/V3/A1/M4/s1 ),
    .B(\V3/V4/V3/A1/c3 ),
    .Z(\V3/V4/V3/s1 [3]));
 OR2_X1 \V3/V4/V3/A1/M4/_0_  (.A1(\V3/V4/V3/A1/M4/c1 ),
    .A2(\V3/V4/V3/A1/M4/c2 ),
    .ZN(\V3/V4/V3/c1 ));
 AND2_X1 \V3/V4/V3/A2/M1/M1/_0_  (.A1(\V3/V4/V3/s1 [0]),
    .A2(\V3/V4/V3/v1 [2]),
    .ZN(\V3/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M1/M1/_1_  (.A(\V3/V4/V3/s1 [0]),
    .B(\V3/V4/V3/v1 [2]),
    .Z(\V3/V4/V3/A2/M1/s1 ));
 AND2_X1 \V3/V4/V3/A2/M1/M2/_0_  (.A1(\V3/V4/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M1/M2/_1_  (.A(\V3/V4/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v3 [2]));
 OR2_X1 \V3/V4/V3/A2/M1/_0_  (.A1(\V3/V4/V3/A2/M1/c1 ),
    .A2(\V3/V4/V3/A2/M1/c2 ),
    .ZN(\V3/V4/V3/A2/c1 ));
 AND2_X1 \V3/V4/V3/A2/M2/M1/_0_  (.A1(\V3/V4/V3/s1 [1]),
    .A2(\V3/V4/V3/v1 [3]),
    .ZN(\V3/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M2/M1/_1_  (.A(\V3/V4/V3/s1 [1]),
    .B(\V3/V4/V3/v1 [3]),
    .Z(\V3/V4/V3/A2/M2/s1 ));
 AND2_X1 \V3/V4/V3/A2/M2/M2/_0_  (.A1(\V3/V4/V3/A2/M2/s1 ),
    .A2(\V3/V4/V3/A2/c1 ),
    .ZN(\V3/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M2/M2/_1_  (.A(\V3/V4/V3/A2/M2/s1 ),
    .B(\V3/V4/V3/A2/c1 ),
    .Z(\V3/V4/v3 [3]));
 OR2_X1 \V3/V4/V3/A2/M2/_0_  (.A1(\V3/V4/V3/A2/M2/c1 ),
    .A2(\V3/V4/V3/A2/M2/c2 ),
    .ZN(\V3/V4/V3/A2/c2 ));
 AND2_X1 \V3/V4/V3/A2/M3/M1/_0_  (.A1(\V3/V4/V3/s1 [2]),
    .A2(ground),
    .ZN(\V3/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M3/M1/_1_  (.A(\V3/V4/V3/s1 [2]),
    .B(ground),
    .Z(\V3/V4/V3/A2/M3/s1 ));
 AND2_X1 \V3/V4/V3/A2/M3/M2/_0_  (.A1(\V3/V4/V3/A2/M3/s1 ),
    .A2(\V3/V4/V3/A2/c2 ),
    .ZN(\V3/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M3/M2/_1_  (.A(\V3/V4/V3/A2/M3/s1 ),
    .B(\V3/V4/V3/A2/c2 ),
    .Z(\V3/V4/V3/s2 [2]));
 OR2_X1 \V3/V4/V3/A2/M3/_0_  (.A1(\V3/V4/V3/A2/M3/c1 ),
    .A2(\V3/V4/V3/A2/M3/c2 ),
    .ZN(\V3/V4/V3/A2/c3 ));
 AND2_X1 \V3/V4/V3/A2/M4/M1/_0_  (.A1(\V3/V4/V3/s1 [3]),
    .A2(ground),
    .ZN(\V3/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M4/M1/_1_  (.A(\V3/V4/V3/s1 [3]),
    .B(ground),
    .Z(\V3/V4/V3/A2/M4/s1 ));
 AND2_X1 \V3/V4/V3/A2/M4/M2/_0_  (.A1(\V3/V4/V3/A2/M4/s1 ),
    .A2(\V3/V4/V3/A2/c3 ),
    .ZN(\V3/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M4/M2/_1_  (.A(\V3/V4/V3/A2/M4/s1 ),
    .B(\V3/V4/V3/A2/c3 ),
    .Z(\V3/V4/V3/s2 [3]));
 OR2_X1 \V3/V4/V3/A2/M4/_0_  (.A1(\V3/V4/V3/A2/M4/c1 ),
    .A2(\V3/V4/V3/A2/M4/c2 ),
    .ZN(\V3/V4/V3/c2 ));
 AND2_X1 \V3/V4/V3/A3/M1/M1/_0_  (.A1(\V3/V4/V3/v4 [0]),
    .A2(\V3/V4/V3/s2 [2]),
    .ZN(\V3/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M1/M1/_1_  (.A(\V3/V4/V3/v4 [0]),
    .B(\V3/V4/V3/s2 [2]),
    .Z(\V3/V4/V3/A3/M1/s1 ));
 AND2_X1 \V3/V4/V3/A3/M1/M2/_0_  (.A1(\V3/V4/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M1/M2/_1_  (.A(\V3/V4/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v3 [4]));
 OR2_X1 \V3/V4/V3/A3/M1/_0_  (.A1(\V3/V4/V3/A3/M1/c1 ),
    .A2(\V3/V4/V3/A3/M1/c2 ),
    .ZN(\V3/V4/V3/A3/c1 ));
 AND2_X1 \V3/V4/V3/A3/M2/M1/_0_  (.A1(\V3/V4/V3/v4 [1]),
    .A2(\V3/V4/V3/s2 [3]),
    .ZN(\V3/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M2/M1/_1_  (.A(\V3/V4/V3/v4 [1]),
    .B(\V3/V4/V3/s2 [3]),
    .Z(\V3/V4/V3/A3/M2/s1 ));
 AND2_X1 \V3/V4/V3/A3/M2/M2/_0_  (.A1(\V3/V4/V3/A3/M2/s1 ),
    .A2(\V3/V4/V3/A3/c1 ),
    .ZN(\V3/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M2/M2/_1_  (.A(\V3/V4/V3/A3/M2/s1 ),
    .B(\V3/V4/V3/A3/c1 ),
    .Z(\V3/V4/v3 [5]));
 OR2_X1 \V3/V4/V3/A3/M2/_0_  (.A1(\V3/V4/V3/A3/M2/c1 ),
    .A2(\V3/V4/V3/A3/M2/c2 ),
    .ZN(\V3/V4/V3/A3/c2 ));
 AND2_X1 \V3/V4/V3/A3/M3/M1/_0_  (.A1(\V3/V4/V3/v4 [2]),
    .A2(\V3/V4/V3/c3 ),
    .ZN(\V3/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M3/M1/_1_  (.A(\V3/V4/V3/v4 [2]),
    .B(\V3/V4/V3/c3 ),
    .Z(\V3/V4/V3/A3/M3/s1 ));
 AND2_X1 \V3/V4/V3/A3/M3/M2/_0_  (.A1(\V3/V4/V3/A3/M3/s1 ),
    .A2(\V3/V4/V3/A3/c2 ),
    .ZN(\V3/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M3/M2/_1_  (.A(\V3/V4/V3/A3/M3/s1 ),
    .B(\V3/V4/V3/A3/c2 ),
    .Z(\V3/V4/v3 [6]));
 OR2_X1 \V3/V4/V3/A3/M3/_0_  (.A1(\V3/V4/V3/A3/M3/c1 ),
    .A2(\V3/V4/V3/A3/M3/c2 ),
    .ZN(\V3/V4/V3/A3/c3 ));
 AND2_X1 \V3/V4/V3/A3/M4/M1/_0_  (.A1(\V3/V4/V3/v4 [3]),
    .A2(ground),
    .ZN(\V3/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M4/M1/_1_  (.A(\V3/V4/V3/v4 [3]),
    .B(ground),
    .Z(\V3/V4/V3/A3/M4/s1 ));
 AND2_X1 \V3/V4/V3/A3/M4/M2/_0_  (.A1(\V3/V4/V3/A3/M4/s1 ),
    .A2(\V3/V4/V3/A3/c3 ),
    .ZN(\V3/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M4/M2/_1_  (.A(\V3/V4/V3/A3/M4/s1 ),
    .B(\V3/V4/V3/A3/c3 ),
    .Z(\V3/V4/v3 [7]));
 OR2_X1 \V3/V4/V3/A3/M4/_0_  (.A1(\V3/V4/V3/A3/M4/c1 ),
    .A2(\V3/V4/V3/A3/M4/c2 ),
    .ZN(\V3/V4/V3/overflow ));
 AND2_X1 \V3/V4/V3/V1/HA1/_0_  (.A1(\V3/V4/V3/V1/w2 ),
    .A2(\V3/V4/V3/V1/w1 ),
    .ZN(\V3/V4/V3/V1/w4 ));
 XOR2_X2 \V3/V4/V3/V1/HA1/_1_  (.A(\V3/V4/V3/V1/w2 ),
    .B(\V3/V4/V3/V1/w1 ),
    .Z(\V3/V4/v3 [1]));
 AND2_X1 \V3/V4/V3/V1/HA2/_0_  (.A1(\V3/V4/V3/V1/w4 ),
    .A2(\V3/V4/V3/V1/w3 ),
    .ZN(\V3/V4/V3/v1 [3]));
 XOR2_X2 \V3/V4/V3/V1/HA2/_1_  (.A(\V3/V4/V3/V1/w4 ),
    .B(\V3/V4/V3/V1/w3 ),
    .Z(\V3/V4/V3/v1 [2]));
 AND2_X1 \V3/V4/V3/V1/_0_  (.A1(A[8]),
    .A2(B[28]),
    .ZN(\V3/V4/v3 [0]));
 AND2_X1 \V3/V4/V3/V1/_1_  (.A1(A[8]),
    .A2(B[29]),
    .ZN(\V3/V4/V3/V1/w1 ));
 AND2_X1 \V3/V4/V3/V1/_2_  (.A1(B[28]),
    .A2(A[9]),
    .ZN(\V3/V4/V3/V1/w2 ));
 AND2_X1 \V3/V4/V3/V1/_3_  (.A1(B[29]),
    .A2(A[9]),
    .ZN(\V3/V4/V3/V1/w3 ));
 AND2_X1 \V3/V4/V3/V2/HA1/_0_  (.A1(\V3/V4/V3/V2/w2 ),
    .A2(\V3/V4/V3/V2/w1 ),
    .ZN(\V3/V4/V3/V2/w4 ));
 XOR2_X2 \V3/V4/V3/V2/HA1/_1_  (.A(\V3/V4/V3/V2/w2 ),
    .B(\V3/V4/V3/V2/w1 ),
    .Z(\V3/V4/V3/v2 [1]));
 AND2_X1 \V3/V4/V3/V2/HA2/_0_  (.A1(\V3/V4/V3/V2/w4 ),
    .A2(\V3/V4/V3/V2/w3 ),
    .ZN(\V3/V4/V3/v2 [3]));
 XOR2_X2 \V3/V4/V3/V2/HA2/_1_  (.A(\V3/V4/V3/V2/w4 ),
    .B(\V3/V4/V3/V2/w3 ),
    .Z(\V3/V4/V3/v2 [2]));
 AND2_X1 \V3/V4/V3/V2/_0_  (.A1(A[10]),
    .A2(B[28]),
    .ZN(\V3/V4/V3/v2 [0]));
 AND2_X1 \V3/V4/V3/V2/_1_  (.A1(A[10]),
    .A2(B[29]),
    .ZN(\V3/V4/V3/V2/w1 ));
 AND2_X1 \V3/V4/V3/V2/_2_  (.A1(B[28]),
    .A2(A[11]),
    .ZN(\V3/V4/V3/V2/w2 ));
 AND2_X1 \V3/V4/V3/V2/_3_  (.A1(B[29]),
    .A2(A[11]),
    .ZN(\V3/V4/V3/V2/w3 ));
 AND2_X1 \V3/V4/V3/V3/HA1/_0_  (.A1(\V3/V4/V3/V3/w2 ),
    .A2(\V3/V4/V3/V3/w1 ),
    .ZN(\V3/V4/V3/V3/w4 ));
 XOR2_X2 \V3/V4/V3/V3/HA1/_1_  (.A(\V3/V4/V3/V3/w2 ),
    .B(\V3/V4/V3/V3/w1 ),
    .Z(\V3/V4/V3/v3 [1]));
 AND2_X1 \V3/V4/V3/V3/HA2/_0_  (.A1(\V3/V4/V3/V3/w4 ),
    .A2(\V3/V4/V3/V3/w3 ),
    .ZN(\V3/V4/V3/v3 [3]));
 XOR2_X2 \V3/V4/V3/V3/HA2/_1_  (.A(\V3/V4/V3/V3/w4 ),
    .B(\V3/V4/V3/V3/w3 ),
    .Z(\V3/V4/V3/v3 [2]));
 AND2_X1 \V3/V4/V3/V3/_0_  (.A1(A[8]),
    .A2(B[30]),
    .ZN(\V3/V4/V3/v3 [0]));
 AND2_X1 \V3/V4/V3/V3/_1_  (.A1(A[8]),
    .A2(B[31]),
    .ZN(\V3/V4/V3/V3/w1 ));
 AND2_X1 \V3/V4/V3/V3/_2_  (.A1(B[30]),
    .A2(A[9]),
    .ZN(\V3/V4/V3/V3/w2 ));
 AND2_X1 \V3/V4/V3/V3/_3_  (.A1(B[31]),
    .A2(A[9]),
    .ZN(\V3/V4/V3/V3/w3 ));
 AND2_X1 \V3/V4/V3/V4/HA1/_0_  (.A1(\V3/V4/V3/V4/w2 ),
    .A2(\V3/V4/V3/V4/w1 ),
    .ZN(\V3/V4/V3/V4/w4 ));
 XOR2_X2 \V3/V4/V3/V4/HA1/_1_  (.A(\V3/V4/V3/V4/w2 ),
    .B(\V3/V4/V3/V4/w1 ),
    .Z(\V3/V4/V3/v4 [1]));
 AND2_X1 \V3/V4/V3/V4/HA2/_0_  (.A1(\V3/V4/V3/V4/w4 ),
    .A2(\V3/V4/V3/V4/w3 ),
    .ZN(\V3/V4/V3/v4 [3]));
 XOR2_X2 \V3/V4/V3/V4/HA2/_1_  (.A(\V3/V4/V3/V4/w4 ),
    .B(\V3/V4/V3/V4/w3 ),
    .Z(\V3/V4/V3/v4 [2]));
 AND2_X1 \V3/V4/V3/V4/_0_  (.A1(A[10]),
    .A2(B[30]),
    .ZN(\V3/V4/V3/v4 [0]));
 AND2_X1 \V3/V4/V3/V4/_1_  (.A1(A[10]),
    .A2(B[31]),
    .ZN(\V3/V4/V3/V4/w1 ));
 AND2_X1 \V3/V4/V3/V4/_2_  (.A1(B[30]),
    .A2(A[11]),
    .ZN(\V3/V4/V3/V4/w2 ));
 AND2_X1 \V3/V4/V3/V4/_3_  (.A1(B[31]),
    .A2(A[11]),
    .ZN(\V3/V4/V3/V4/w3 ));
 OR2_X1 \V3/V4/V3/_0_  (.A1(\V3/V4/V3/c1 ),
    .A2(\V3/V4/V3/c2 ),
    .ZN(\V3/V4/V3/c3 ));
 AND2_X1 \V3/V4/V4/A1/M1/M1/_0_  (.A1(\V3/V4/V4/v2 [0]),
    .A2(\V3/V4/V4/v3 [0]),
    .ZN(\V3/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M1/M1/_1_  (.A(\V3/V4/V4/v2 [0]),
    .B(\V3/V4/V4/v3 [0]),
    .Z(\V3/V4/V4/A1/M1/s1 ));
 AND2_X1 \V3/V4/V4/A1/M1/M2/_0_  (.A1(\V3/V4/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M1/M2/_1_  (.A(\V3/V4/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/V4/s1 [0]));
 OR2_X1 \V3/V4/V4/A1/M1/_0_  (.A1(\V3/V4/V4/A1/M1/c1 ),
    .A2(\V3/V4/V4/A1/M1/c2 ),
    .ZN(\V3/V4/V4/A1/c1 ));
 AND2_X1 \V3/V4/V4/A1/M2/M1/_0_  (.A1(\V3/V4/V4/v2 [1]),
    .A2(\V3/V4/V4/v3 [1]),
    .ZN(\V3/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M2/M1/_1_  (.A(\V3/V4/V4/v2 [1]),
    .B(\V3/V4/V4/v3 [1]),
    .Z(\V3/V4/V4/A1/M2/s1 ));
 AND2_X1 \V3/V4/V4/A1/M2/M2/_0_  (.A1(\V3/V4/V4/A1/M2/s1 ),
    .A2(\V3/V4/V4/A1/c1 ),
    .ZN(\V3/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M2/M2/_1_  (.A(\V3/V4/V4/A1/M2/s1 ),
    .B(\V3/V4/V4/A1/c1 ),
    .Z(\V3/V4/V4/s1 [1]));
 OR2_X1 \V3/V4/V4/A1/M2/_0_  (.A1(\V3/V4/V4/A1/M2/c1 ),
    .A2(\V3/V4/V4/A1/M2/c2 ),
    .ZN(\V3/V4/V4/A1/c2 ));
 AND2_X1 \V3/V4/V4/A1/M3/M1/_0_  (.A1(\V3/V4/V4/v2 [2]),
    .A2(\V3/V4/V4/v3 [2]),
    .ZN(\V3/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M3/M1/_1_  (.A(\V3/V4/V4/v2 [2]),
    .B(\V3/V4/V4/v3 [2]),
    .Z(\V3/V4/V4/A1/M3/s1 ));
 AND2_X1 \V3/V4/V4/A1/M3/M2/_0_  (.A1(\V3/V4/V4/A1/M3/s1 ),
    .A2(\V3/V4/V4/A1/c2 ),
    .ZN(\V3/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M3/M2/_1_  (.A(\V3/V4/V4/A1/M3/s1 ),
    .B(\V3/V4/V4/A1/c2 ),
    .Z(\V3/V4/V4/s1 [2]));
 OR2_X1 \V3/V4/V4/A1/M3/_0_  (.A1(\V3/V4/V4/A1/M3/c1 ),
    .A2(\V3/V4/V4/A1/M3/c2 ),
    .ZN(\V3/V4/V4/A1/c3 ));
 AND2_X1 \V3/V4/V4/A1/M4/M1/_0_  (.A1(\V3/V4/V4/v2 [3]),
    .A2(\V3/V4/V4/v3 [3]),
    .ZN(\V3/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M4/M1/_1_  (.A(\V3/V4/V4/v2 [3]),
    .B(\V3/V4/V4/v3 [3]),
    .Z(\V3/V4/V4/A1/M4/s1 ));
 AND2_X1 \V3/V4/V4/A1/M4/M2/_0_  (.A1(\V3/V4/V4/A1/M4/s1 ),
    .A2(\V3/V4/V4/A1/c3 ),
    .ZN(\V3/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M4/M2/_1_  (.A(\V3/V4/V4/A1/M4/s1 ),
    .B(\V3/V4/V4/A1/c3 ),
    .Z(\V3/V4/V4/s1 [3]));
 OR2_X1 \V3/V4/V4/A1/M4/_0_  (.A1(\V3/V4/V4/A1/M4/c1 ),
    .A2(\V3/V4/V4/A1/M4/c2 ),
    .ZN(\V3/V4/V4/c1 ));
 AND2_X1 \V3/V4/V4/A2/M1/M1/_0_  (.A1(\V3/V4/V4/s1 [0]),
    .A2(\V3/V4/V4/v1 [2]),
    .ZN(\V3/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M1/M1/_1_  (.A(\V3/V4/V4/s1 [0]),
    .B(\V3/V4/V4/v1 [2]),
    .Z(\V3/V4/V4/A2/M1/s1 ));
 AND2_X1 \V3/V4/V4/A2/M1/M2/_0_  (.A1(\V3/V4/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M1/M2/_1_  (.A(\V3/V4/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v4 [2]));
 OR2_X1 \V3/V4/V4/A2/M1/_0_  (.A1(\V3/V4/V4/A2/M1/c1 ),
    .A2(\V3/V4/V4/A2/M1/c2 ),
    .ZN(\V3/V4/V4/A2/c1 ));
 AND2_X1 \V3/V4/V4/A2/M2/M1/_0_  (.A1(\V3/V4/V4/s1 [1]),
    .A2(\V3/V4/V4/v1 [3]),
    .ZN(\V3/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M2/M1/_1_  (.A(\V3/V4/V4/s1 [1]),
    .B(\V3/V4/V4/v1 [3]),
    .Z(\V3/V4/V4/A2/M2/s1 ));
 AND2_X1 \V3/V4/V4/A2/M2/M2/_0_  (.A1(\V3/V4/V4/A2/M2/s1 ),
    .A2(\V3/V4/V4/A2/c1 ),
    .ZN(\V3/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M2/M2/_1_  (.A(\V3/V4/V4/A2/M2/s1 ),
    .B(\V3/V4/V4/A2/c1 ),
    .Z(\V3/V4/v4 [3]));
 OR2_X1 \V3/V4/V4/A2/M2/_0_  (.A1(\V3/V4/V4/A2/M2/c1 ),
    .A2(\V3/V4/V4/A2/M2/c2 ),
    .ZN(\V3/V4/V4/A2/c2 ));
 AND2_X1 \V3/V4/V4/A2/M3/M1/_0_  (.A1(\V3/V4/V4/s1 [2]),
    .A2(ground),
    .ZN(\V3/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M3/M1/_1_  (.A(\V3/V4/V4/s1 [2]),
    .B(ground),
    .Z(\V3/V4/V4/A2/M3/s1 ));
 AND2_X1 \V3/V4/V4/A2/M3/M2/_0_  (.A1(\V3/V4/V4/A2/M3/s1 ),
    .A2(\V3/V4/V4/A2/c2 ),
    .ZN(\V3/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M3/M2/_1_  (.A(\V3/V4/V4/A2/M3/s1 ),
    .B(\V3/V4/V4/A2/c2 ),
    .Z(\V3/V4/V4/s2 [2]));
 OR2_X1 \V3/V4/V4/A2/M3/_0_  (.A1(\V3/V4/V4/A2/M3/c1 ),
    .A2(\V3/V4/V4/A2/M3/c2 ),
    .ZN(\V3/V4/V4/A2/c3 ));
 AND2_X1 \V3/V4/V4/A2/M4/M1/_0_  (.A1(\V3/V4/V4/s1 [3]),
    .A2(ground),
    .ZN(\V3/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M4/M1/_1_  (.A(\V3/V4/V4/s1 [3]),
    .B(ground),
    .Z(\V3/V4/V4/A2/M4/s1 ));
 AND2_X1 \V3/V4/V4/A2/M4/M2/_0_  (.A1(\V3/V4/V4/A2/M4/s1 ),
    .A2(\V3/V4/V4/A2/c3 ),
    .ZN(\V3/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M4/M2/_1_  (.A(\V3/V4/V4/A2/M4/s1 ),
    .B(\V3/V4/V4/A2/c3 ),
    .Z(\V3/V4/V4/s2 [3]));
 OR2_X1 \V3/V4/V4/A2/M4/_0_  (.A1(\V3/V4/V4/A2/M4/c1 ),
    .A2(\V3/V4/V4/A2/M4/c2 ),
    .ZN(\V3/V4/V4/c2 ));
 AND2_X1 \V3/V4/V4/A3/M1/M1/_0_  (.A1(\V3/V4/V4/v4 [0]),
    .A2(\V3/V4/V4/s2 [2]),
    .ZN(\V3/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M1/M1/_1_  (.A(\V3/V4/V4/v4 [0]),
    .B(\V3/V4/V4/s2 [2]),
    .Z(\V3/V4/V4/A3/M1/s1 ));
 AND2_X1 \V3/V4/V4/A3/M1/M2/_0_  (.A1(\V3/V4/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V3/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M1/M2/_1_  (.A(\V3/V4/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V3/V4/v4 [4]));
 OR2_X1 \V3/V4/V4/A3/M1/_0_  (.A1(\V3/V4/V4/A3/M1/c1 ),
    .A2(\V3/V4/V4/A3/M1/c2 ),
    .ZN(\V3/V4/V4/A3/c1 ));
 AND2_X1 \V3/V4/V4/A3/M2/M1/_0_  (.A1(\V3/V4/V4/v4 [1]),
    .A2(\V3/V4/V4/s2 [3]),
    .ZN(\V3/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M2/M1/_1_  (.A(\V3/V4/V4/v4 [1]),
    .B(\V3/V4/V4/s2 [3]),
    .Z(\V3/V4/V4/A3/M2/s1 ));
 AND2_X1 \V3/V4/V4/A3/M2/M2/_0_  (.A1(\V3/V4/V4/A3/M2/s1 ),
    .A2(\V3/V4/V4/A3/c1 ),
    .ZN(\V3/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M2/M2/_1_  (.A(\V3/V4/V4/A3/M2/s1 ),
    .B(\V3/V4/V4/A3/c1 ),
    .Z(\V3/V4/v4 [5]));
 OR2_X1 \V3/V4/V4/A3/M2/_0_  (.A1(\V3/V4/V4/A3/M2/c1 ),
    .A2(\V3/V4/V4/A3/M2/c2 ),
    .ZN(\V3/V4/V4/A3/c2 ));
 AND2_X1 \V3/V4/V4/A3/M3/M1/_0_  (.A1(\V3/V4/V4/v4 [2]),
    .A2(\V3/V4/V4/c3 ),
    .ZN(\V3/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M3/M1/_1_  (.A(\V3/V4/V4/v4 [2]),
    .B(\V3/V4/V4/c3 ),
    .Z(\V3/V4/V4/A3/M3/s1 ));
 AND2_X1 \V3/V4/V4/A3/M3/M2/_0_  (.A1(\V3/V4/V4/A3/M3/s1 ),
    .A2(\V3/V4/V4/A3/c2 ),
    .ZN(\V3/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M3/M2/_1_  (.A(\V3/V4/V4/A3/M3/s1 ),
    .B(\V3/V4/V4/A3/c2 ),
    .Z(\V3/V4/v4 [6]));
 OR2_X1 \V3/V4/V4/A3/M3/_0_  (.A1(\V3/V4/V4/A3/M3/c1 ),
    .A2(\V3/V4/V4/A3/M3/c2 ),
    .ZN(\V3/V4/V4/A3/c3 ));
 AND2_X1 \V3/V4/V4/A3/M4/M1/_0_  (.A1(\V3/V4/V4/v4 [3]),
    .A2(ground),
    .ZN(\V3/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M4/M1/_1_  (.A(\V3/V4/V4/v4 [3]),
    .B(ground),
    .Z(\V3/V4/V4/A3/M4/s1 ));
 AND2_X1 \V3/V4/V4/A3/M4/M2/_0_  (.A1(\V3/V4/V4/A3/M4/s1 ),
    .A2(\V3/V4/V4/A3/c3 ),
    .ZN(\V3/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M4/M2/_1_  (.A(\V3/V4/V4/A3/M4/s1 ),
    .B(\V3/V4/V4/A3/c3 ),
    .Z(\V3/V4/v4 [7]));
 OR2_X1 \V3/V4/V4/A3/M4/_0_  (.A1(\V3/V4/V4/A3/M4/c1 ),
    .A2(\V3/V4/V4/A3/M4/c2 ),
    .ZN(\V3/V4/V4/overflow ));
 AND2_X1 \V3/V4/V4/V1/HA1/_0_  (.A1(\V3/V4/V4/V1/w2 ),
    .A2(\V3/V4/V4/V1/w1 ),
    .ZN(\V3/V4/V4/V1/w4 ));
 XOR2_X2 \V3/V4/V4/V1/HA1/_1_  (.A(\V3/V4/V4/V1/w2 ),
    .B(\V3/V4/V4/V1/w1 ),
    .Z(\V3/V4/v4 [1]));
 AND2_X1 \V3/V4/V4/V1/HA2/_0_  (.A1(\V3/V4/V4/V1/w4 ),
    .A2(\V3/V4/V4/V1/w3 ),
    .ZN(\V3/V4/V4/v1 [3]));
 XOR2_X2 \V3/V4/V4/V1/HA2/_1_  (.A(\V3/V4/V4/V1/w4 ),
    .B(\V3/V4/V4/V1/w3 ),
    .Z(\V3/V4/V4/v1 [2]));
 AND2_X1 \V3/V4/V4/V1/_0_  (.A1(A[12]),
    .A2(B[28]),
    .ZN(\V3/V4/v4 [0]));
 AND2_X1 \V3/V4/V4/V1/_1_  (.A1(A[12]),
    .A2(B[29]),
    .ZN(\V3/V4/V4/V1/w1 ));
 AND2_X1 \V3/V4/V4/V1/_2_  (.A1(B[28]),
    .A2(A[13]),
    .ZN(\V3/V4/V4/V1/w2 ));
 AND2_X1 \V3/V4/V4/V1/_3_  (.A1(B[29]),
    .A2(A[13]),
    .ZN(\V3/V4/V4/V1/w3 ));
 AND2_X1 \V3/V4/V4/V2/HA1/_0_  (.A1(\V3/V4/V4/V2/w2 ),
    .A2(\V3/V4/V4/V2/w1 ),
    .ZN(\V3/V4/V4/V2/w4 ));
 XOR2_X2 \V3/V4/V4/V2/HA1/_1_  (.A(\V3/V4/V4/V2/w2 ),
    .B(\V3/V4/V4/V2/w1 ),
    .Z(\V3/V4/V4/v2 [1]));
 AND2_X1 \V3/V4/V4/V2/HA2/_0_  (.A1(\V3/V4/V4/V2/w4 ),
    .A2(\V3/V4/V4/V2/w3 ),
    .ZN(\V3/V4/V4/v2 [3]));
 XOR2_X2 \V3/V4/V4/V2/HA2/_1_  (.A(\V3/V4/V4/V2/w4 ),
    .B(\V3/V4/V4/V2/w3 ),
    .Z(\V3/V4/V4/v2 [2]));
 AND2_X1 \V3/V4/V4/V2/_0_  (.A1(A[14]),
    .A2(B[28]),
    .ZN(\V3/V4/V4/v2 [0]));
 AND2_X1 \V3/V4/V4/V2/_1_  (.A1(A[14]),
    .A2(B[29]),
    .ZN(\V3/V4/V4/V2/w1 ));
 AND2_X1 \V3/V4/V4/V2/_2_  (.A1(B[28]),
    .A2(A[15]),
    .ZN(\V3/V4/V4/V2/w2 ));
 AND2_X1 \V3/V4/V4/V2/_3_  (.A1(B[29]),
    .A2(A[15]),
    .ZN(\V3/V4/V4/V2/w3 ));
 AND2_X1 \V3/V4/V4/V3/HA1/_0_  (.A1(\V3/V4/V4/V3/w2 ),
    .A2(\V3/V4/V4/V3/w1 ),
    .ZN(\V3/V4/V4/V3/w4 ));
 XOR2_X2 \V3/V4/V4/V3/HA1/_1_  (.A(\V3/V4/V4/V3/w2 ),
    .B(\V3/V4/V4/V3/w1 ),
    .Z(\V3/V4/V4/v3 [1]));
 AND2_X1 \V3/V4/V4/V3/HA2/_0_  (.A1(\V3/V4/V4/V3/w4 ),
    .A2(\V3/V4/V4/V3/w3 ),
    .ZN(\V3/V4/V4/v3 [3]));
 XOR2_X2 \V3/V4/V4/V3/HA2/_1_  (.A(\V3/V4/V4/V3/w4 ),
    .B(\V3/V4/V4/V3/w3 ),
    .Z(\V3/V4/V4/v3 [2]));
 AND2_X1 \V3/V4/V4/V3/_0_  (.A1(A[12]),
    .A2(B[30]),
    .ZN(\V3/V4/V4/v3 [0]));
 AND2_X1 \V3/V4/V4/V3/_1_  (.A1(A[12]),
    .A2(B[31]),
    .ZN(\V3/V4/V4/V3/w1 ));
 AND2_X1 \V3/V4/V4/V3/_2_  (.A1(B[30]),
    .A2(A[13]),
    .ZN(\V3/V4/V4/V3/w2 ));
 AND2_X1 \V3/V4/V4/V3/_3_  (.A1(B[31]),
    .A2(A[13]),
    .ZN(\V3/V4/V4/V3/w3 ));
 AND2_X1 \V3/V4/V4/V4/HA1/_0_  (.A1(\V3/V4/V4/V4/w2 ),
    .A2(\V3/V4/V4/V4/w1 ),
    .ZN(\V3/V4/V4/V4/w4 ));
 XOR2_X2 \V3/V4/V4/V4/HA1/_1_  (.A(\V3/V4/V4/V4/w2 ),
    .B(\V3/V4/V4/V4/w1 ),
    .Z(\V3/V4/V4/v4 [1]));
 AND2_X1 \V3/V4/V4/V4/HA2/_0_  (.A1(\V3/V4/V4/V4/w4 ),
    .A2(\V3/V4/V4/V4/w3 ),
    .ZN(\V3/V4/V4/v4 [3]));
 XOR2_X2 \V3/V4/V4/V4/HA2/_1_  (.A(\V3/V4/V4/V4/w4 ),
    .B(\V3/V4/V4/V4/w3 ),
    .Z(\V3/V4/V4/v4 [2]));
 AND2_X1 \V3/V4/V4/V4/_0_  (.A1(A[14]),
    .A2(B[30]),
    .ZN(\V3/V4/V4/v4 [0]));
 AND2_X1 \V3/V4/V4/V4/_1_  (.A1(A[14]),
    .A2(B[31]),
    .ZN(\V3/V4/V4/V4/w1 ));
 AND2_X1 \V3/V4/V4/V4/_2_  (.A1(B[30]),
    .A2(A[15]),
    .ZN(\V3/V4/V4/V4/w2 ));
 AND2_X1 \V3/V4/V4/V4/_3_  (.A1(B[31]),
    .A2(A[15]),
    .ZN(\V3/V4/V4/V4/w3 ));
 OR2_X1 \V3/V4/V4/_0_  (.A1(\V3/V4/V4/c1 ),
    .A2(\V3/V4/V4/c2 ),
    .ZN(\V3/V4/V4/c3 ));
 OR2_X1 \V3/V4/_0_  (.A1(\V3/V4/c1 ),
    .A2(\V3/V4/c2 ),
    .ZN(\V3/V4/c3 ));
 OR2_X2 \V3/_0_  (.A1(\V3/c1 ),
    .A2(\V3/c2 ),
    .ZN(\V3/c3 ));
 AND2_X1 \V4/A1/A1/A1/M1/M1/_0_  (.A1(\V4/v2 [0]),
    .A2(\V4/v3 [0]),
    .ZN(\V4/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M1/M1/_1_  (.A(\V4/v2 [0]),
    .B(\V4/v3 [0]),
    .Z(\V4/A1/A1/A1/M1/s1 ));
 AND2_X1 \V4/A1/A1/A1/M1/M2/_0_  (.A1(\V4/A1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M1/M2/_1_  (.A(\V4/A1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/s1 [0]));
 OR2_X1 \V4/A1/A1/A1/M1/_0_  (.A1(\V4/A1/A1/A1/M1/c1 ),
    .A2(\V4/A1/A1/A1/M1/c2 ),
    .ZN(\V4/A1/A1/A1/c1 ));
 AND2_X1 \V4/A1/A1/A1/M2/M1/_0_  (.A1(\V4/v2 [1]),
    .A2(\V4/v3 [1]),
    .ZN(\V4/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M2/M1/_1_  (.A(\V4/v2 [1]),
    .B(\V4/v3 [1]),
    .Z(\V4/A1/A1/A1/M2/s1 ));
 AND2_X1 \V4/A1/A1/A1/M2/M2/_0_  (.A1(\V4/A1/A1/A1/M2/s1 ),
    .A2(\V4/A1/A1/A1/c1 ),
    .ZN(\V4/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M2/M2/_1_  (.A(\V4/A1/A1/A1/M2/s1 ),
    .B(\V4/A1/A1/A1/c1 ),
    .Z(\V4/s1 [1]));
 OR2_X1 \V4/A1/A1/A1/M2/_0_  (.A1(\V4/A1/A1/A1/M2/c1 ),
    .A2(\V4/A1/A1/A1/M2/c2 ),
    .ZN(\V4/A1/A1/A1/c2 ));
 AND2_X1 \V4/A1/A1/A1/M3/M1/_0_  (.A1(\V4/v2 [2]),
    .A2(\V4/v3 [2]),
    .ZN(\V4/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M3/M1/_1_  (.A(\V4/v2 [2]),
    .B(\V4/v3 [2]),
    .Z(\V4/A1/A1/A1/M3/s1 ));
 AND2_X1 \V4/A1/A1/A1/M3/M2/_0_  (.A1(\V4/A1/A1/A1/M3/s1 ),
    .A2(\V4/A1/A1/A1/c2 ),
    .ZN(\V4/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M3/M2/_1_  (.A(\V4/A1/A1/A1/M3/s1 ),
    .B(\V4/A1/A1/A1/c2 ),
    .Z(\V4/s1 [2]));
 OR2_X1 \V4/A1/A1/A1/M3/_0_  (.A1(\V4/A1/A1/A1/M3/c1 ),
    .A2(\V4/A1/A1/A1/M3/c2 ),
    .ZN(\V4/A1/A1/A1/c3 ));
 AND2_X1 \V4/A1/A1/A1/M4/M1/_0_  (.A1(\V4/v2 [3]),
    .A2(\V4/v3 [3]),
    .ZN(\V4/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M4/M1/_1_  (.A(\V4/v2 [3]),
    .B(\V4/v3 [3]),
    .Z(\V4/A1/A1/A1/M4/s1 ));
 AND2_X1 \V4/A1/A1/A1/M4/M2/_0_  (.A1(\V4/A1/A1/A1/M4/s1 ),
    .A2(\V4/A1/A1/A1/c3 ),
    .ZN(\V4/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M4/M2/_1_  (.A(\V4/A1/A1/A1/M4/s1 ),
    .B(\V4/A1/A1/A1/c3 ),
    .Z(\V4/s1 [3]));
 OR2_X1 \V4/A1/A1/A1/M4/_0_  (.A1(\V4/A1/A1/A1/M4/c1 ),
    .A2(\V4/A1/A1/A1/M4/c2 ),
    .ZN(\V4/A1/A1/c1 ));
 AND2_X1 \V4/A1/A1/A2/M1/M1/_0_  (.A1(\V4/v2 [4]),
    .A2(\V4/v3 [4]),
    .ZN(\V4/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M1/M1/_1_  (.A(\V4/v2 [4]),
    .B(\V4/v3 [4]),
    .Z(\V4/A1/A1/A2/M1/s1 ));
 AND2_X1 \V4/A1/A1/A2/M1/M2/_0_  (.A1(\V4/A1/A1/A2/M1/s1 ),
    .A2(\V4/A1/A1/c1 ),
    .ZN(\V4/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M1/M2/_1_  (.A(\V4/A1/A1/A2/M1/s1 ),
    .B(\V4/A1/A1/c1 ),
    .Z(\V4/s1 [4]));
 OR2_X1 \V4/A1/A1/A2/M1/_0_  (.A1(\V4/A1/A1/A2/M1/c1 ),
    .A2(\V4/A1/A1/A2/M1/c2 ),
    .ZN(\V4/A1/A1/A2/c1 ));
 AND2_X1 \V4/A1/A1/A2/M2/M1/_0_  (.A1(\V4/v2 [5]),
    .A2(\V4/v3 [5]),
    .ZN(\V4/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M2/M1/_1_  (.A(\V4/v2 [5]),
    .B(\V4/v3 [5]),
    .Z(\V4/A1/A1/A2/M2/s1 ));
 AND2_X1 \V4/A1/A1/A2/M2/M2/_0_  (.A1(\V4/A1/A1/A2/M2/s1 ),
    .A2(\V4/A1/A1/A2/c1 ),
    .ZN(\V4/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M2/M2/_1_  (.A(\V4/A1/A1/A2/M2/s1 ),
    .B(\V4/A1/A1/A2/c1 ),
    .Z(\V4/s1 [5]));
 OR2_X1 \V4/A1/A1/A2/M2/_0_  (.A1(\V4/A1/A1/A2/M2/c1 ),
    .A2(\V4/A1/A1/A2/M2/c2 ),
    .ZN(\V4/A1/A1/A2/c2 ));
 AND2_X1 \V4/A1/A1/A2/M3/M1/_0_  (.A1(\V4/v2 [6]),
    .A2(\V4/v3 [6]),
    .ZN(\V4/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M3/M1/_1_  (.A(\V4/v2 [6]),
    .B(\V4/v3 [6]),
    .Z(\V4/A1/A1/A2/M3/s1 ));
 AND2_X1 \V4/A1/A1/A2/M3/M2/_0_  (.A1(\V4/A1/A1/A2/M3/s1 ),
    .A2(\V4/A1/A1/A2/c2 ),
    .ZN(\V4/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M3/M2/_1_  (.A(\V4/A1/A1/A2/M3/s1 ),
    .B(\V4/A1/A1/A2/c2 ),
    .Z(\V4/s1 [6]));
 OR2_X1 \V4/A1/A1/A2/M3/_0_  (.A1(\V4/A1/A1/A2/M3/c1 ),
    .A2(\V4/A1/A1/A2/M3/c2 ),
    .ZN(\V4/A1/A1/A2/c3 ));
 AND2_X1 \V4/A1/A1/A2/M4/M1/_0_  (.A1(\V4/v2 [7]),
    .A2(\V4/v3 [7]),
    .ZN(\V4/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M4/M1/_1_  (.A(\V4/v2 [7]),
    .B(\V4/v3 [7]),
    .Z(\V4/A1/A1/A2/M4/s1 ));
 AND2_X1 \V4/A1/A1/A2/M4/M2/_0_  (.A1(\V4/A1/A1/A2/M4/s1 ),
    .A2(\V4/A1/A1/A2/c3 ),
    .ZN(\V4/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M4/M2/_1_  (.A(\V4/A1/A1/A2/M4/s1 ),
    .B(\V4/A1/A1/A2/c3 ),
    .Z(\V4/s1 [7]));
 OR2_X1 \V4/A1/A1/A2/M4/_0_  (.A1(\V4/A1/A1/A2/M4/c1 ),
    .A2(\V4/A1/A1/A2/M4/c2 ),
    .ZN(\V4/A1/c1 ));
 AND2_X1 \V4/A1/A2/A1/M1/M1/_0_  (.A1(\V4/v2 [8]),
    .A2(\V4/v3 [8]),
    .ZN(\V4/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M1/M1/_1_  (.A(\V4/v2 [8]),
    .B(\V4/v3 [8]),
    .Z(\V4/A1/A2/A1/M1/s1 ));
 AND2_X1 \V4/A1/A2/A1/M1/M2/_0_  (.A1(\V4/A1/A2/A1/M1/s1 ),
    .A2(\V4/A1/c1 ),
    .ZN(\V4/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M1/M2/_1_  (.A(\V4/A1/A2/A1/M1/s1 ),
    .B(\V4/A1/c1 ),
    .Z(\V4/s1 [8]));
 OR2_X1 \V4/A1/A2/A1/M1/_0_  (.A1(\V4/A1/A2/A1/M1/c1 ),
    .A2(\V4/A1/A2/A1/M1/c2 ),
    .ZN(\V4/A1/A2/A1/c1 ));
 AND2_X1 \V4/A1/A2/A1/M2/M1/_0_  (.A1(\V4/v2 [9]),
    .A2(\V4/v3 [9]),
    .ZN(\V4/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M2/M1/_1_  (.A(\V4/v2 [9]),
    .B(\V4/v3 [9]),
    .Z(\V4/A1/A2/A1/M2/s1 ));
 AND2_X1 \V4/A1/A2/A1/M2/M2/_0_  (.A1(\V4/A1/A2/A1/M2/s1 ),
    .A2(\V4/A1/A2/A1/c1 ),
    .ZN(\V4/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M2/M2/_1_  (.A(\V4/A1/A2/A1/M2/s1 ),
    .B(\V4/A1/A2/A1/c1 ),
    .Z(\V4/s1 [9]));
 OR2_X1 \V4/A1/A2/A1/M2/_0_  (.A1(\V4/A1/A2/A1/M2/c1 ),
    .A2(\V4/A1/A2/A1/M2/c2 ),
    .ZN(\V4/A1/A2/A1/c2 ));
 AND2_X1 \V4/A1/A2/A1/M3/M1/_0_  (.A1(\V4/v2 [10]),
    .A2(\V4/v3 [10]),
    .ZN(\V4/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M3/M1/_1_  (.A(\V4/v2 [10]),
    .B(\V4/v3 [10]),
    .Z(\V4/A1/A2/A1/M3/s1 ));
 AND2_X1 \V4/A1/A2/A1/M3/M2/_0_  (.A1(\V4/A1/A2/A1/M3/s1 ),
    .A2(\V4/A1/A2/A1/c2 ),
    .ZN(\V4/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M3/M2/_1_  (.A(\V4/A1/A2/A1/M3/s1 ),
    .B(\V4/A1/A2/A1/c2 ),
    .Z(\V4/s1 [10]));
 OR2_X1 \V4/A1/A2/A1/M3/_0_  (.A1(\V4/A1/A2/A1/M3/c1 ),
    .A2(\V4/A1/A2/A1/M3/c2 ),
    .ZN(\V4/A1/A2/A1/c3 ));
 AND2_X1 \V4/A1/A2/A1/M4/M1/_0_  (.A1(\V4/v2 [11]),
    .A2(\V4/v3 [11]),
    .ZN(\V4/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M4/M1/_1_  (.A(\V4/v2 [11]),
    .B(\V4/v3 [11]),
    .Z(\V4/A1/A2/A1/M4/s1 ));
 AND2_X1 \V4/A1/A2/A1/M4/M2/_0_  (.A1(\V4/A1/A2/A1/M4/s1 ),
    .A2(\V4/A1/A2/A1/c3 ),
    .ZN(\V4/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M4/M2/_1_  (.A(\V4/A1/A2/A1/M4/s1 ),
    .B(\V4/A1/A2/A1/c3 ),
    .Z(\V4/s1 [11]));
 OR2_X1 \V4/A1/A2/A1/M4/_0_  (.A1(\V4/A1/A2/A1/M4/c1 ),
    .A2(\V4/A1/A2/A1/M4/c2 ),
    .ZN(\V4/A1/A2/c1 ));
 AND2_X1 \V4/A1/A2/A2/M1/M1/_0_  (.A1(\V4/v2 [12]),
    .A2(\V4/v3 [12]),
    .ZN(\V4/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M1/M1/_1_  (.A(\V4/v2 [12]),
    .B(\V4/v3 [12]),
    .Z(\V4/A1/A2/A2/M1/s1 ));
 AND2_X1 \V4/A1/A2/A2/M1/M2/_0_  (.A1(\V4/A1/A2/A2/M1/s1 ),
    .A2(\V4/A1/A2/c1 ),
    .ZN(\V4/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M1/M2/_1_  (.A(\V4/A1/A2/A2/M1/s1 ),
    .B(\V4/A1/A2/c1 ),
    .Z(\V4/s1 [12]));
 OR2_X1 \V4/A1/A2/A2/M1/_0_  (.A1(\V4/A1/A2/A2/M1/c1 ),
    .A2(\V4/A1/A2/A2/M1/c2 ),
    .ZN(\V4/A1/A2/A2/c1 ));
 AND2_X1 \V4/A1/A2/A2/M2/M1/_0_  (.A1(\V4/v2 [13]),
    .A2(\V4/v3 [13]),
    .ZN(\V4/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M2/M1/_1_  (.A(\V4/v2 [13]),
    .B(\V4/v3 [13]),
    .Z(\V4/A1/A2/A2/M2/s1 ));
 AND2_X1 \V4/A1/A2/A2/M2/M2/_0_  (.A1(\V4/A1/A2/A2/M2/s1 ),
    .A2(\V4/A1/A2/A2/c1 ),
    .ZN(\V4/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M2/M2/_1_  (.A(\V4/A1/A2/A2/M2/s1 ),
    .B(\V4/A1/A2/A2/c1 ),
    .Z(\V4/s1 [13]));
 OR2_X1 \V4/A1/A2/A2/M2/_0_  (.A1(\V4/A1/A2/A2/M2/c1 ),
    .A2(\V4/A1/A2/A2/M2/c2 ),
    .ZN(\V4/A1/A2/A2/c2 ));
 AND2_X1 \V4/A1/A2/A2/M3/M1/_0_  (.A1(\V4/v2 [14]),
    .A2(\V4/v3 [14]),
    .ZN(\V4/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M3/M1/_1_  (.A(\V4/v2 [14]),
    .B(\V4/v3 [14]),
    .Z(\V4/A1/A2/A2/M3/s1 ));
 AND2_X1 \V4/A1/A2/A2/M3/M2/_0_  (.A1(\V4/A1/A2/A2/M3/s1 ),
    .A2(\V4/A1/A2/A2/c2 ),
    .ZN(\V4/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M3/M2/_1_  (.A(\V4/A1/A2/A2/M3/s1 ),
    .B(\V4/A1/A2/A2/c2 ),
    .Z(\V4/s1 [14]));
 OR2_X1 \V4/A1/A2/A2/M3/_0_  (.A1(\V4/A1/A2/A2/M3/c1 ),
    .A2(\V4/A1/A2/A2/M3/c2 ),
    .ZN(\V4/A1/A2/A2/c3 ));
 AND2_X1 \V4/A1/A2/A2/M4/M1/_0_  (.A1(\V4/v2 [15]),
    .A2(\V4/v3 [15]),
    .ZN(\V4/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M4/M1/_1_  (.A(\V4/v2 [15]),
    .B(\V4/v3 [15]),
    .Z(\V4/A1/A2/A2/M4/s1 ));
 AND2_X1 \V4/A1/A2/A2/M4/M2/_0_  (.A1(\V4/A1/A2/A2/M4/s1 ),
    .A2(\V4/A1/A2/A2/c3 ),
    .ZN(\V4/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M4/M2/_1_  (.A(\V4/A1/A2/A2/M4/s1 ),
    .B(\V4/A1/A2/A2/c3 ),
    .Z(\V4/s1 [15]));
 OR2_X1 \V4/A1/A2/A2/M4/_0_  (.A1(\V4/A1/A2/A2/M4/c1 ),
    .A2(\V4/A1/A2/A2/M4/c2 ),
    .ZN(\V4/c1 ));
 AND2_X1 \V4/A2/A1/A1/M1/M1/_0_  (.A1(\V4/s1 [0]),
    .A2(\V4/v1 [8]),
    .ZN(\V4/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M1/M1/_1_  (.A(\V4/s1 [0]),
    .B(\V4/v1 [8]),
    .Z(\V4/A2/A1/A1/M1/s1 ));
 AND2_X1 \V4/A2/A1/A1/M1/M2/_0_  (.A1(\V4/A2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M1/M2/_1_  (.A(\V4/A2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v4[8]));
 OR2_X1 \V4/A2/A1/A1/M1/_0_  (.A1(\V4/A2/A1/A1/M1/c1 ),
    .A2(\V4/A2/A1/A1/M1/c2 ),
    .ZN(\V4/A2/A1/A1/c1 ));
 AND2_X1 \V4/A2/A1/A1/M2/M1/_0_  (.A1(\V4/s1 [1]),
    .A2(\V4/v1 [9]),
    .ZN(\V4/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M2/M1/_1_  (.A(\V4/s1 [1]),
    .B(\V4/v1 [9]),
    .Z(\V4/A2/A1/A1/M2/s1 ));
 AND2_X1 \V4/A2/A1/A1/M2/M2/_0_  (.A1(\V4/A2/A1/A1/M2/s1 ),
    .A2(\V4/A2/A1/A1/c1 ),
    .ZN(\V4/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M2/M2/_1_  (.A(\V4/A2/A1/A1/M2/s1 ),
    .B(\V4/A2/A1/A1/c1 ),
    .Z(v4[9]));
 OR2_X1 \V4/A2/A1/A1/M2/_0_  (.A1(\V4/A2/A1/A1/M2/c1 ),
    .A2(\V4/A2/A1/A1/M2/c2 ),
    .ZN(\V4/A2/A1/A1/c2 ));
 AND2_X1 \V4/A2/A1/A1/M3/M1/_0_  (.A1(\V4/s1 [2]),
    .A2(\V4/v1 [10]),
    .ZN(\V4/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M3/M1/_1_  (.A(\V4/s1 [2]),
    .B(\V4/v1 [10]),
    .Z(\V4/A2/A1/A1/M3/s1 ));
 AND2_X1 \V4/A2/A1/A1/M3/M2/_0_  (.A1(\V4/A2/A1/A1/M3/s1 ),
    .A2(\V4/A2/A1/A1/c2 ),
    .ZN(\V4/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M3/M2/_1_  (.A(\V4/A2/A1/A1/M3/s1 ),
    .B(\V4/A2/A1/A1/c2 ),
    .Z(v4[10]));
 OR2_X1 \V4/A2/A1/A1/M3/_0_  (.A1(\V4/A2/A1/A1/M3/c1 ),
    .A2(\V4/A2/A1/A1/M3/c2 ),
    .ZN(\V4/A2/A1/A1/c3 ));
 AND2_X1 \V4/A2/A1/A1/M4/M1/_0_  (.A1(\V4/s1 [3]),
    .A2(\V4/v1 [11]),
    .ZN(\V4/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M4/M1/_1_  (.A(\V4/s1 [3]),
    .B(\V4/v1 [11]),
    .Z(\V4/A2/A1/A1/M4/s1 ));
 AND2_X1 \V4/A2/A1/A1/M4/M2/_0_  (.A1(\V4/A2/A1/A1/M4/s1 ),
    .A2(\V4/A2/A1/A1/c3 ),
    .ZN(\V4/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M4/M2/_1_  (.A(\V4/A2/A1/A1/M4/s1 ),
    .B(\V4/A2/A1/A1/c3 ),
    .Z(v4[11]));
 OR2_X1 \V4/A2/A1/A1/M4/_0_  (.A1(\V4/A2/A1/A1/M4/c1 ),
    .A2(\V4/A2/A1/A1/M4/c2 ),
    .ZN(\V4/A2/A1/c1 ));
 AND2_X1 \V4/A2/A1/A2/M1/M1/_0_  (.A1(\V4/s1 [4]),
    .A2(\V4/v1 [12]),
    .ZN(\V4/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M1/M1/_1_  (.A(\V4/s1 [4]),
    .B(\V4/v1 [12]),
    .Z(\V4/A2/A1/A2/M1/s1 ));
 AND2_X1 \V4/A2/A1/A2/M1/M2/_0_  (.A1(\V4/A2/A1/A2/M1/s1 ),
    .A2(\V4/A2/A1/c1 ),
    .ZN(\V4/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M1/M2/_1_  (.A(\V4/A2/A1/A2/M1/s1 ),
    .B(\V4/A2/A1/c1 ),
    .Z(v4[12]));
 OR2_X1 \V4/A2/A1/A2/M1/_0_  (.A1(\V4/A2/A1/A2/M1/c1 ),
    .A2(\V4/A2/A1/A2/M1/c2 ),
    .ZN(\V4/A2/A1/A2/c1 ));
 AND2_X1 \V4/A2/A1/A2/M2/M1/_0_  (.A1(\V4/s1 [5]),
    .A2(\V4/v1 [13]),
    .ZN(\V4/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M2/M1/_1_  (.A(\V4/s1 [5]),
    .B(\V4/v1 [13]),
    .Z(\V4/A2/A1/A2/M2/s1 ));
 AND2_X1 \V4/A2/A1/A2/M2/M2/_0_  (.A1(\V4/A2/A1/A2/M2/s1 ),
    .A2(\V4/A2/A1/A2/c1 ),
    .ZN(\V4/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M2/M2/_1_  (.A(\V4/A2/A1/A2/M2/s1 ),
    .B(\V4/A2/A1/A2/c1 ),
    .Z(v4[13]));
 OR2_X1 \V4/A2/A1/A2/M2/_0_  (.A1(\V4/A2/A1/A2/M2/c1 ),
    .A2(\V4/A2/A1/A2/M2/c2 ),
    .ZN(\V4/A2/A1/A2/c2 ));
 AND2_X1 \V4/A2/A1/A2/M3/M1/_0_  (.A1(\V4/s1 [6]),
    .A2(\V4/v1 [14]),
    .ZN(\V4/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M3/M1/_1_  (.A(\V4/s1 [6]),
    .B(\V4/v1 [14]),
    .Z(\V4/A2/A1/A2/M3/s1 ));
 AND2_X1 \V4/A2/A1/A2/M3/M2/_0_  (.A1(\V4/A2/A1/A2/M3/s1 ),
    .A2(\V4/A2/A1/A2/c2 ),
    .ZN(\V4/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M3/M2/_1_  (.A(\V4/A2/A1/A2/M3/s1 ),
    .B(\V4/A2/A1/A2/c2 ),
    .Z(v4[14]));
 OR2_X1 \V4/A2/A1/A2/M3/_0_  (.A1(\V4/A2/A1/A2/M3/c1 ),
    .A2(\V4/A2/A1/A2/M3/c2 ),
    .ZN(\V4/A2/A1/A2/c3 ));
 AND2_X1 \V4/A2/A1/A2/M4/M1/_0_  (.A1(\V4/s1 [7]),
    .A2(\V4/v1 [15]),
    .ZN(\V4/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M4/M1/_1_  (.A(\V4/s1 [7]),
    .B(\V4/v1 [15]),
    .Z(\V4/A2/A1/A2/M4/s1 ));
 AND2_X1 \V4/A2/A1/A2/M4/M2/_0_  (.A1(\V4/A2/A1/A2/M4/s1 ),
    .A2(\V4/A2/A1/A2/c3 ),
    .ZN(\V4/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M4/M2/_1_  (.A(\V4/A2/A1/A2/M4/s1 ),
    .B(\V4/A2/A1/A2/c3 ),
    .Z(v4[15]));
 OR2_X1 \V4/A2/A1/A2/M4/_0_  (.A1(\V4/A2/A1/A2/M4/c1 ),
    .A2(\V4/A2/A1/A2/M4/c2 ),
    .ZN(\V4/A2/c1 ));
 AND2_X1 \V4/A2/A2/A1/M1/M1/_0_  (.A1(\V4/s1 [8]),
    .A2(ground),
    .ZN(\V4/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M1/M1/_1_  (.A(\V4/s1 [8]),
    .B(ground),
    .Z(\V4/A2/A2/A1/M1/s1 ));
 AND2_X1 \V4/A2/A2/A1/M1/M2/_0_  (.A1(\V4/A2/A2/A1/M1/s1 ),
    .A2(\V4/A2/c1 ),
    .ZN(\V4/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M1/M2/_1_  (.A(\V4/A2/A2/A1/M1/s1 ),
    .B(\V4/A2/c1 ),
    .Z(\V4/s2 [8]));
 OR2_X1 \V4/A2/A2/A1/M1/_0_  (.A1(\V4/A2/A2/A1/M1/c1 ),
    .A2(\V4/A2/A2/A1/M1/c2 ),
    .ZN(\V4/A2/A2/A1/c1 ));
 AND2_X1 \V4/A2/A2/A1/M2/M1/_0_  (.A1(\V4/s1 [9]),
    .A2(ground),
    .ZN(\V4/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M2/M1/_1_  (.A(\V4/s1 [9]),
    .B(ground),
    .Z(\V4/A2/A2/A1/M2/s1 ));
 AND2_X1 \V4/A2/A2/A1/M2/M2/_0_  (.A1(\V4/A2/A2/A1/M2/s1 ),
    .A2(\V4/A2/A2/A1/c1 ),
    .ZN(\V4/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M2/M2/_1_  (.A(\V4/A2/A2/A1/M2/s1 ),
    .B(\V4/A2/A2/A1/c1 ),
    .Z(\V4/s2 [9]));
 OR2_X1 \V4/A2/A2/A1/M2/_0_  (.A1(\V4/A2/A2/A1/M2/c1 ),
    .A2(\V4/A2/A2/A1/M2/c2 ),
    .ZN(\V4/A2/A2/A1/c2 ));
 AND2_X1 \V4/A2/A2/A1/M3/M1/_0_  (.A1(\V4/s1 [10]),
    .A2(ground),
    .ZN(\V4/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M3/M1/_1_  (.A(\V4/s1 [10]),
    .B(ground),
    .Z(\V4/A2/A2/A1/M3/s1 ));
 AND2_X1 \V4/A2/A2/A1/M3/M2/_0_  (.A1(\V4/A2/A2/A1/M3/s1 ),
    .A2(\V4/A2/A2/A1/c2 ),
    .ZN(\V4/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M3/M2/_1_  (.A(\V4/A2/A2/A1/M3/s1 ),
    .B(\V4/A2/A2/A1/c2 ),
    .Z(\V4/s2 [10]));
 OR2_X1 \V4/A2/A2/A1/M3/_0_  (.A1(\V4/A2/A2/A1/M3/c1 ),
    .A2(\V4/A2/A2/A1/M3/c2 ),
    .ZN(\V4/A2/A2/A1/c3 ));
 AND2_X1 \V4/A2/A2/A1/M4/M1/_0_  (.A1(\V4/s1 [11]),
    .A2(ground),
    .ZN(\V4/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M4/M1/_1_  (.A(\V4/s1 [11]),
    .B(ground),
    .Z(\V4/A2/A2/A1/M4/s1 ));
 AND2_X1 \V4/A2/A2/A1/M4/M2/_0_  (.A1(\V4/A2/A2/A1/M4/s1 ),
    .A2(\V4/A2/A2/A1/c3 ),
    .ZN(\V4/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M4/M2/_1_  (.A(\V4/A2/A2/A1/M4/s1 ),
    .B(\V4/A2/A2/A1/c3 ),
    .Z(\V4/s2 [11]));
 OR2_X1 \V4/A2/A2/A1/M4/_0_  (.A1(\V4/A2/A2/A1/M4/c1 ),
    .A2(\V4/A2/A2/A1/M4/c2 ),
    .ZN(\V4/A2/A2/c1 ));
 AND2_X1 \V4/A2/A2/A2/M1/M1/_0_  (.A1(\V4/s1 [12]),
    .A2(ground),
    .ZN(\V4/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M1/M1/_1_  (.A(\V4/s1 [12]),
    .B(ground),
    .Z(\V4/A2/A2/A2/M1/s1 ));
 AND2_X1 \V4/A2/A2/A2/M1/M2/_0_  (.A1(\V4/A2/A2/A2/M1/s1 ),
    .A2(\V4/A2/A2/c1 ),
    .ZN(\V4/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M1/M2/_1_  (.A(\V4/A2/A2/A2/M1/s1 ),
    .B(\V4/A2/A2/c1 ),
    .Z(\V4/s2 [12]));
 OR2_X1 \V4/A2/A2/A2/M1/_0_  (.A1(\V4/A2/A2/A2/M1/c1 ),
    .A2(\V4/A2/A2/A2/M1/c2 ),
    .ZN(\V4/A2/A2/A2/c1 ));
 AND2_X1 \V4/A2/A2/A2/M2/M1/_0_  (.A1(\V4/s1 [13]),
    .A2(ground),
    .ZN(\V4/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M2/M1/_1_  (.A(\V4/s1 [13]),
    .B(ground),
    .Z(\V4/A2/A2/A2/M2/s1 ));
 AND2_X1 \V4/A2/A2/A2/M2/M2/_0_  (.A1(\V4/A2/A2/A2/M2/s1 ),
    .A2(\V4/A2/A2/A2/c1 ),
    .ZN(\V4/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M2/M2/_1_  (.A(\V4/A2/A2/A2/M2/s1 ),
    .B(\V4/A2/A2/A2/c1 ),
    .Z(\V4/s2 [13]));
 OR2_X1 \V4/A2/A2/A2/M2/_0_  (.A1(\V4/A2/A2/A2/M2/c1 ),
    .A2(\V4/A2/A2/A2/M2/c2 ),
    .ZN(\V4/A2/A2/A2/c2 ));
 AND2_X1 \V4/A2/A2/A2/M3/M1/_0_  (.A1(\V4/s1 [14]),
    .A2(ground),
    .ZN(\V4/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M3/M1/_1_  (.A(\V4/s1 [14]),
    .B(ground),
    .Z(\V4/A2/A2/A2/M3/s1 ));
 AND2_X1 \V4/A2/A2/A2/M3/M2/_0_  (.A1(\V4/A2/A2/A2/M3/s1 ),
    .A2(\V4/A2/A2/A2/c2 ),
    .ZN(\V4/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M3/M2/_1_  (.A(\V4/A2/A2/A2/M3/s1 ),
    .B(\V4/A2/A2/A2/c2 ),
    .Z(\V4/s2 [14]));
 OR2_X1 \V4/A2/A2/A2/M3/_0_  (.A1(\V4/A2/A2/A2/M3/c1 ),
    .A2(\V4/A2/A2/A2/M3/c2 ),
    .ZN(\V4/A2/A2/A2/c3 ));
 AND2_X1 \V4/A2/A2/A2/M4/M1/_0_  (.A1(\V4/s1 [15]),
    .A2(ground),
    .ZN(\V4/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M4/M1/_1_  (.A(\V4/s1 [15]),
    .B(ground),
    .Z(\V4/A2/A2/A2/M4/s1 ));
 AND2_X1 \V4/A2/A2/A2/M4/M2/_0_  (.A1(\V4/A2/A2/A2/M4/s1 ),
    .A2(\V4/A2/A2/A2/c3 ),
    .ZN(\V4/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M4/M2/_1_  (.A(\V4/A2/A2/A2/M4/s1 ),
    .B(\V4/A2/A2/A2/c3 ),
    .Z(\V4/s2 [15]));
 OR2_X1 \V4/A2/A2/A2/M4/_0_  (.A1(\V4/A2/A2/A2/M4/c1 ),
    .A2(\V4/A2/A2/A2/M4/c2 ),
    .ZN(\V4/c2 ));
 AND2_X1 \V4/A3/A1/A1/M1/M1/_0_  (.A1(\V4/v4 [0]),
    .A2(\V4/s2 [8]),
    .ZN(\V4/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M1/M1/_1_  (.A(\V4/v4 [0]),
    .B(\V4/s2 [8]),
    .Z(\V4/A3/A1/A1/M1/s1 ));
 AND2_X1 \V4/A3/A1/A1/M1/M2/_0_  (.A1(\V4/A3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M1/M2/_1_  (.A(\V4/A3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(v4[16]));
 OR2_X1 \V4/A3/A1/A1/M1/_0_  (.A1(\V4/A3/A1/A1/M1/c1 ),
    .A2(\V4/A3/A1/A1/M1/c2 ),
    .ZN(\V4/A3/A1/A1/c1 ));
 AND2_X1 \V4/A3/A1/A1/M2/M1/_0_  (.A1(\V4/v4 [1]),
    .A2(\V4/s2 [9]),
    .ZN(\V4/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M2/M1/_1_  (.A(\V4/v4 [1]),
    .B(\V4/s2 [9]),
    .Z(\V4/A3/A1/A1/M2/s1 ));
 AND2_X1 \V4/A3/A1/A1/M2/M2/_0_  (.A1(\V4/A3/A1/A1/M2/s1 ),
    .A2(\V4/A3/A1/A1/c1 ),
    .ZN(\V4/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M2/M2/_1_  (.A(\V4/A3/A1/A1/M2/s1 ),
    .B(\V4/A3/A1/A1/c1 ),
    .Z(v4[17]));
 OR2_X1 \V4/A3/A1/A1/M2/_0_  (.A1(\V4/A3/A1/A1/M2/c1 ),
    .A2(\V4/A3/A1/A1/M2/c2 ),
    .ZN(\V4/A3/A1/A1/c2 ));
 AND2_X1 \V4/A3/A1/A1/M3/M1/_0_  (.A1(\V4/v4 [2]),
    .A2(\V4/s2 [10]),
    .ZN(\V4/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M3/M1/_1_  (.A(\V4/v4 [2]),
    .B(\V4/s2 [10]),
    .Z(\V4/A3/A1/A1/M3/s1 ));
 AND2_X1 \V4/A3/A1/A1/M3/M2/_0_  (.A1(\V4/A3/A1/A1/M3/s1 ),
    .A2(\V4/A3/A1/A1/c2 ),
    .ZN(\V4/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M3/M2/_1_  (.A(\V4/A3/A1/A1/M3/s1 ),
    .B(\V4/A3/A1/A1/c2 ),
    .Z(v4[18]));
 OR2_X1 \V4/A3/A1/A1/M3/_0_  (.A1(\V4/A3/A1/A1/M3/c1 ),
    .A2(\V4/A3/A1/A1/M3/c2 ),
    .ZN(\V4/A3/A1/A1/c3 ));
 AND2_X1 \V4/A3/A1/A1/M4/M1/_0_  (.A1(\V4/v4 [3]),
    .A2(\V4/s2 [11]),
    .ZN(\V4/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M4/M1/_1_  (.A(\V4/v4 [3]),
    .B(\V4/s2 [11]),
    .Z(\V4/A3/A1/A1/M4/s1 ));
 AND2_X1 \V4/A3/A1/A1/M4/M2/_0_  (.A1(\V4/A3/A1/A1/M4/s1 ),
    .A2(\V4/A3/A1/A1/c3 ),
    .ZN(\V4/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M4/M2/_1_  (.A(\V4/A3/A1/A1/M4/s1 ),
    .B(\V4/A3/A1/A1/c3 ),
    .Z(v4[19]));
 OR2_X1 \V4/A3/A1/A1/M4/_0_  (.A1(\V4/A3/A1/A1/M4/c1 ),
    .A2(\V4/A3/A1/A1/M4/c2 ),
    .ZN(\V4/A3/A1/c1 ));
 AND2_X1 \V4/A3/A1/A2/M1/M1/_0_  (.A1(\V4/v4 [4]),
    .A2(\V4/s2 [12]),
    .ZN(\V4/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M1/M1/_1_  (.A(\V4/v4 [4]),
    .B(\V4/s2 [12]),
    .Z(\V4/A3/A1/A2/M1/s1 ));
 AND2_X1 \V4/A3/A1/A2/M1/M2/_0_  (.A1(\V4/A3/A1/A2/M1/s1 ),
    .A2(\V4/A3/A1/c1 ),
    .ZN(\V4/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M1/M2/_1_  (.A(\V4/A3/A1/A2/M1/s1 ),
    .B(\V4/A3/A1/c1 ),
    .Z(v4[20]));
 OR2_X1 \V4/A3/A1/A2/M1/_0_  (.A1(\V4/A3/A1/A2/M1/c1 ),
    .A2(\V4/A3/A1/A2/M1/c2 ),
    .ZN(\V4/A3/A1/A2/c1 ));
 AND2_X1 \V4/A3/A1/A2/M2/M1/_0_  (.A1(\V4/v4 [5]),
    .A2(\V4/s2 [13]),
    .ZN(\V4/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M2/M1/_1_  (.A(\V4/v4 [5]),
    .B(\V4/s2 [13]),
    .Z(\V4/A3/A1/A2/M2/s1 ));
 AND2_X1 \V4/A3/A1/A2/M2/M2/_0_  (.A1(\V4/A3/A1/A2/M2/s1 ),
    .A2(\V4/A3/A1/A2/c1 ),
    .ZN(\V4/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M2/M2/_1_  (.A(\V4/A3/A1/A2/M2/s1 ),
    .B(\V4/A3/A1/A2/c1 ),
    .Z(v4[21]));
 OR2_X1 \V4/A3/A1/A2/M2/_0_  (.A1(\V4/A3/A1/A2/M2/c1 ),
    .A2(\V4/A3/A1/A2/M2/c2 ),
    .ZN(\V4/A3/A1/A2/c2 ));
 AND2_X1 \V4/A3/A1/A2/M3/M1/_0_  (.A1(\V4/v4 [6]),
    .A2(\V4/s2 [14]),
    .ZN(\V4/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M3/M1/_1_  (.A(\V4/v4 [6]),
    .B(\V4/s2 [14]),
    .Z(\V4/A3/A1/A2/M3/s1 ));
 AND2_X1 \V4/A3/A1/A2/M3/M2/_0_  (.A1(\V4/A3/A1/A2/M3/s1 ),
    .A2(\V4/A3/A1/A2/c2 ),
    .ZN(\V4/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M3/M2/_1_  (.A(\V4/A3/A1/A2/M3/s1 ),
    .B(\V4/A3/A1/A2/c2 ),
    .Z(v4[22]));
 OR2_X1 \V4/A3/A1/A2/M3/_0_  (.A1(\V4/A3/A1/A2/M3/c1 ),
    .A2(\V4/A3/A1/A2/M3/c2 ),
    .ZN(\V4/A3/A1/A2/c3 ));
 AND2_X1 \V4/A3/A1/A2/M4/M1/_0_  (.A1(\V4/v4 [7]),
    .A2(\V4/s2 [15]),
    .ZN(\V4/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M4/M1/_1_  (.A(\V4/v4 [7]),
    .B(\V4/s2 [15]),
    .Z(\V4/A3/A1/A2/M4/s1 ));
 AND2_X1 \V4/A3/A1/A2/M4/M2/_0_  (.A1(\V4/A3/A1/A2/M4/s1 ),
    .A2(\V4/A3/A1/A2/c3 ),
    .ZN(\V4/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M4/M2/_1_  (.A(\V4/A3/A1/A2/M4/s1 ),
    .B(\V4/A3/A1/A2/c3 ),
    .Z(v4[23]));
 OR2_X1 \V4/A3/A1/A2/M4/_0_  (.A1(\V4/A3/A1/A2/M4/c1 ),
    .A2(\V4/A3/A1/A2/M4/c2 ),
    .ZN(\V4/A3/c1 ));
 AND2_X1 \V4/A3/A2/A1/M1/M1/_0_  (.A1(\V4/v4 [8]),
    .A2(\V4/c3 ),
    .ZN(\V4/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M1/M1/_1_  (.A(\V4/v4 [8]),
    .B(\V4/c3 ),
    .Z(\V4/A3/A2/A1/M1/s1 ));
 AND2_X1 \V4/A3/A2/A1/M1/M2/_0_  (.A1(\V4/A3/A2/A1/M1/s1 ),
    .A2(\V4/A3/c1 ),
    .ZN(\V4/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M1/M2/_1_  (.A(\V4/A3/A2/A1/M1/s1 ),
    .B(\V4/A3/c1 ),
    .Z(v4[24]));
 OR2_X1 \V4/A3/A2/A1/M1/_0_  (.A1(\V4/A3/A2/A1/M1/c1 ),
    .A2(\V4/A3/A2/A1/M1/c2 ),
    .ZN(\V4/A3/A2/A1/c1 ));
 AND2_X1 \V4/A3/A2/A1/M2/M1/_0_  (.A1(\V4/v4 [9]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M2/M1/_1_  (.A(\V4/v4 [9]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M2/s1 ));
 AND2_X1 \V4/A3/A2/A1/M2/M2/_0_  (.A1(\V4/A3/A2/A1/M2/s1 ),
    .A2(\V4/A3/A2/A1/c1 ),
    .ZN(\V4/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M2/M2/_1_  (.A(\V4/A3/A2/A1/M2/s1 ),
    .B(\V4/A3/A2/A1/c1 ),
    .Z(v4[25]));
 OR2_X1 \V4/A3/A2/A1/M2/_0_  (.A1(\V4/A3/A2/A1/M2/c1 ),
    .A2(\V4/A3/A2/A1/M2/c2 ),
    .ZN(\V4/A3/A2/A1/c2 ));
 AND2_X1 \V4/A3/A2/A1/M3/M1/_0_  (.A1(\V4/v4 [10]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M3/M1/_1_  (.A(\V4/v4 [10]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M3/s1 ));
 AND2_X1 \V4/A3/A2/A1/M3/M2/_0_  (.A1(\V4/A3/A2/A1/M3/s1 ),
    .A2(\V4/A3/A2/A1/c2 ),
    .ZN(\V4/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M3/M2/_1_  (.A(\V4/A3/A2/A1/M3/s1 ),
    .B(\V4/A3/A2/A1/c2 ),
    .Z(v4[26]));
 OR2_X1 \V4/A3/A2/A1/M3/_0_  (.A1(\V4/A3/A2/A1/M3/c1 ),
    .A2(\V4/A3/A2/A1/M3/c2 ),
    .ZN(\V4/A3/A2/A1/c3 ));
 AND2_X1 \V4/A3/A2/A1/M4/M1/_0_  (.A1(\V4/v4 [11]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M4/c1 ));
 XOR2_X1 \V4/A3/A2/A1/M4/M1/_1_  (.A(\V4/v4 [11]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M4/s1 ));
 AND2_X1 \V4/A3/A2/A1/M4/M2/_0_  (.A1(\V4/A3/A2/A1/M4/s1 ),
    .A2(\V4/A3/A2/A1/c3 ),
    .ZN(\V4/A3/A2/A1/M4/c2 ));
 XOR2_X1 \V4/A3/A2/A1/M4/M2/_1_  (.A(\V4/A3/A2/A1/M4/s1 ),
    .B(\V4/A3/A2/A1/c3 ),
    .Z(v4[27]));
 OR2_X1 \V4/A3/A2/A1/M4/_0_  (.A1(\V4/A3/A2/A1/M4/c1 ),
    .A2(\V4/A3/A2/A1/M4/c2 ),
    .ZN(\V4/A3/A2/c1 ));
 AND2_X1 \V4/A3/A2/A2/M1/M1/_0_  (.A1(\V4/v4 [12]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M1/M1/_1_  (.A(\V4/v4 [12]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M1/s1 ));
 AND2_X1 \V4/A3/A2/A2/M1/M2/_0_  (.A1(\V4/A3/A2/A2/M1/s1 ),
    .A2(\V4/A3/A2/c1 ),
    .ZN(\V4/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M1/M2/_1_  (.A(\V4/A3/A2/A2/M1/s1 ),
    .B(\V4/A3/A2/c1 ),
    .Z(v4[28]));
 OR2_X1 \V4/A3/A2/A2/M1/_0_  (.A1(\V4/A3/A2/A2/M1/c1 ),
    .A2(\V4/A3/A2/A2/M1/c2 ),
    .ZN(\V4/A3/A2/A2/c1 ));
 AND2_X1 \V4/A3/A2/A2/M2/M1/_0_  (.A1(\V4/v4 [13]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M2/M1/_1_  (.A(\V4/v4 [13]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M2/s1 ));
 AND2_X1 \V4/A3/A2/A2/M2/M2/_0_  (.A1(\V4/A3/A2/A2/M2/s1 ),
    .A2(\V4/A3/A2/A2/c1 ),
    .ZN(\V4/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M2/M2/_1_  (.A(\V4/A3/A2/A2/M2/s1 ),
    .B(\V4/A3/A2/A2/c1 ),
    .Z(v4[29]));
 OR2_X1 \V4/A3/A2/A2/M2/_0_  (.A1(\V4/A3/A2/A2/M2/c1 ),
    .A2(\V4/A3/A2/A2/M2/c2 ),
    .ZN(\V4/A3/A2/A2/c2 ));
 AND2_X1 \V4/A3/A2/A2/M3/M1/_0_  (.A1(\V4/v4 [14]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M3/c1 ));
 XOR2_X1 \V4/A3/A2/A2/M3/M1/_1_  (.A(\V4/v4 [14]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M3/s1 ));
 AND2_X1 \V4/A3/A2/A2/M3/M2/_0_  (.A1(\V4/A3/A2/A2/M3/s1 ),
    .A2(\V4/A3/A2/A2/c2 ),
    .ZN(\V4/A3/A2/A2/M3/c2 ));
 XOR2_X1 \V4/A3/A2/A2/M3/M2/_1_  (.A(\V4/A3/A2/A2/M3/s1 ),
    .B(\V4/A3/A2/A2/c2 ),
    .Z(v4[30]));
 OR2_X1 \V4/A3/A2/A2/M3/_0_  (.A1(\V4/A3/A2/A2/M3/c1 ),
    .A2(\V4/A3/A2/A2/M3/c2 ),
    .ZN(\V4/A3/A2/A2/c3 ));
 AND2_X1 \V4/A3/A2/A2/M4/M1/_0_  (.A1(\V4/v4 [15]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M4/M1/_1_  (.A(\V4/v4 [15]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M4/s1 ));
 AND2_X1 \V4/A3/A2/A2/M4/M2/_0_  (.A1(\V4/A3/A2/A2/M4/s1 ),
    .A2(\V4/A3/A2/A2/c3 ),
    .ZN(\V4/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M4/M2/_1_  (.A(\V4/A3/A2/A2/M4/s1 ),
    .B(\V4/A3/A2/A2/c3 ),
    .Z(v4[31]));
 OR2_X1 \V4/A3/A2/A2/M4/_0_  (.A1(\V4/A3/A2/A2/M4/c1 ),
    .A2(\V4/A3/A2/A2/M4/c2 ),
    .ZN(\V4/overflow ));
 AND2_X1 \V4/V1/A1/A1/M1/M1/_0_  (.A1(\V4/V1/v2 [0]),
    .A2(\V4/V1/v3 [0]),
    .ZN(\V4/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M1/M1/_1_  (.A(\V4/V1/v2 [0]),
    .B(\V4/V1/v3 [0]),
    .Z(\V4/V1/A1/A1/M1/s1 ));
 AND2_X1 \V4/V1/A1/A1/M1/M2/_0_  (.A1(\V4/V1/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M1/M2/_1_  (.A(\V4/V1/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/s1 [0]));
 OR2_X1 \V4/V1/A1/A1/M1/_0_  (.A1(\V4/V1/A1/A1/M1/c1 ),
    .A2(\V4/V1/A1/A1/M1/c2 ),
    .ZN(\V4/V1/A1/A1/c1 ));
 AND2_X1 \V4/V1/A1/A1/M2/M1/_0_  (.A1(\V4/V1/v2 [1]),
    .A2(\V4/V1/v3 [1]),
    .ZN(\V4/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M2/M1/_1_  (.A(\V4/V1/v2 [1]),
    .B(\V4/V1/v3 [1]),
    .Z(\V4/V1/A1/A1/M2/s1 ));
 AND2_X1 \V4/V1/A1/A1/M2/M2/_0_  (.A1(\V4/V1/A1/A1/M2/s1 ),
    .A2(\V4/V1/A1/A1/c1 ),
    .ZN(\V4/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M2/M2/_1_  (.A(\V4/V1/A1/A1/M2/s1 ),
    .B(\V4/V1/A1/A1/c1 ),
    .Z(\V4/V1/s1 [1]));
 OR2_X1 \V4/V1/A1/A1/M2/_0_  (.A1(\V4/V1/A1/A1/M2/c1 ),
    .A2(\V4/V1/A1/A1/M2/c2 ),
    .ZN(\V4/V1/A1/A1/c2 ));
 AND2_X1 \V4/V1/A1/A1/M3/M1/_0_  (.A1(\V4/V1/v2 [2]),
    .A2(\V4/V1/v3 [2]),
    .ZN(\V4/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M3/M1/_1_  (.A(\V4/V1/v2 [2]),
    .B(\V4/V1/v3 [2]),
    .Z(\V4/V1/A1/A1/M3/s1 ));
 AND2_X1 \V4/V1/A1/A1/M3/M2/_0_  (.A1(\V4/V1/A1/A1/M3/s1 ),
    .A2(\V4/V1/A1/A1/c2 ),
    .ZN(\V4/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M3/M2/_1_  (.A(\V4/V1/A1/A1/M3/s1 ),
    .B(\V4/V1/A1/A1/c2 ),
    .Z(\V4/V1/s1 [2]));
 OR2_X1 \V4/V1/A1/A1/M3/_0_  (.A1(\V4/V1/A1/A1/M3/c1 ),
    .A2(\V4/V1/A1/A1/M3/c2 ),
    .ZN(\V4/V1/A1/A1/c3 ));
 AND2_X1 \V4/V1/A1/A1/M4/M1/_0_  (.A1(\V4/V1/v2 [3]),
    .A2(\V4/V1/v3 [3]),
    .ZN(\V4/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M4/M1/_1_  (.A(\V4/V1/v2 [3]),
    .B(\V4/V1/v3 [3]),
    .Z(\V4/V1/A1/A1/M4/s1 ));
 AND2_X1 \V4/V1/A1/A1/M4/M2/_0_  (.A1(\V4/V1/A1/A1/M4/s1 ),
    .A2(\V4/V1/A1/A1/c3 ),
    .ZN(\V4/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M4/M2/_1_  (.A(\V4/V1/A1/A1/M4/s1 ),
    .B(\V4/V1/A1/A1/c3 ),
    .Z(\V4/V1/s1 [3]));
 OR2_X1 \V4/V1/A1/A1/M4/_0_  (.A1(\V4/V1/A1/A1/M4/c1 ),
    .A2(\V4/V1/A1/A1/M4/c2 ),
    .ZN(\V4/V1/A1/c1 ));
 AND2_X1 \V4/V1/A1/A2/M1/M1/_0_  (.A1(\V4/V1/v2 [4]),
    .A2(\V4/V1/v3 [4]),
    .ZN(\V4/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M1/M1/_1_  (.A(\V4/V1/v2 [4]),
    .B(\V4/V1/v3 [4]),
    .Z(\V4/V1/A1/A2/M1/s1 ));
 AND2_X1 \V4/V1/A1/A2/M1/M2/_0_  (.A1(\V4/V1/A1/A2/M1/s1 ),
    .A2(\V4/V1/A1/c1 ),
    .ZN(\V4/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M1/M2/_1_  (.A(\V4/V1/A1/A2/M1/s1 ),
    .B(\V4/V1/A1/c1 ),
    .Z(\V4/V1/s1 [4]));
 OR2_X1 \V4/V1/A1/A2/M1/_0_  (.A1(\V4/V1/A1/A2/M1/c1 ),
    .A2(\V4/V1/A1/A2/M1/c2 ),
    .ZN(\V4/V1/A1/A2/c1 ));
 AND2_X1 \V4/V1/A1/A2/M2/M1/_0_  (.A1(\V4/V1/v2 [5]),
    .A2(\V4/V1/v3 [5]),
    .ZN(\V4/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M2/M1/_1_  (.A(\V4/V1/v2 [5]),
    .B(\V4/V1/v3 [5]),
    .Z(\V4/V1/A1/A2/M2/s1 ));
 AND2_X1 \V4/V1/A1/A2/M2/M2/_0_  (.A1(\V4/V1/A1/A2/M2/s1 ),
    .A2(\V4/V1/A1/A2/c1 ),
    .ZN(\V4/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M2/M2/_1_  (.A(\V4/V1/A1/A2/M2/s1 ),
    .B(\V4/V1/A1/A2/c1 ),
    .Z(\V4/V1/s1 [5]));
 OR2_X1 \V4/V1/A1/A2/M2/_0_  (.A1(\V4/V1/A1/A2/M2/c1 ),
    .A2(\V4/V1/A1/A2/M2/c2 ),
    .ZN(\V4/V1/A1/A2/c2 ));
 AND2_X1 \V4/V1/A1/A2/M3/M1/_0_  (.A1(\V4/V1/v2 [6]),
    .A2(\V4/V1/v3 [6]),
    .ZN(\V4/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M3/M1/_1_  (.A(\V4/V1/v2 [6]),
    .B(\V4/V1/v3 [6]),
    .Z(\V4/V1/A1/A2/M3/s1 ));
 AND2_X1 \V4/V1/A1/A2/M3/M2/_0_  (.A1(\V4/V1/A1/A2/M3/s1 ),
    .A2(\V4/V1/A1/A2/c2 ),
    .ZN(\V4/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M3/M2/_1_  (.A(\V4/V1/A1/A2/M3/s1 ),
    .B(\V4/V1/A1/A2/c2 ),
    .Z(\V4/V1/s1 [6]));
 OR2_X1 \V4/V1/A1/A2/M3/_0_  (.A1(\V4/V1/A1/A2/M3/c1 ),
    .A2(\V4/V1/A1/A2/M3/c2 ),
    .ZN(\V4/V1/A1/A2/c3 ));
 AND2_X1 \V4/V1/A1/A2/M4/M1/_0_  (.A1(\V4/V1/v2 [7]),
    .A2(\V4/V1/v3 [7]),
    .ZN(\V4/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M4/M1/_1_  (.A(\V4/V1/v2 [7]),
    .B(\V4/V1/v3 [7]),
    .Z(\V4/V1/A1/A2/M4/s1 ));
 AND2_X1 \V4/V1/A1/A2/M4/M2/_0_  (.A1(\V4/V1/A1/A2/M4/s1 ),
    .A2(\V4/V1/A1/A2/c3 ),
    .ZN(\V4/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M4/M2/_1_  (.A(\V4/V1/A1/A2/M4/s1 ),
    .B(\V4/V1/A1/A2/c3 ),
    .Z(\V4/V1/s1 [7]));
 OR2_X1 \V4/V1/A1/A2/M4/_0_  (.A1(\V4/V1/A1/A2/M4/c1 ),
    .A2(\V4/V1/A1/A2/M4/c2 ),
    .ZN(\V4/V1/c1 ));
 AND2_X1 \V4/V1/A2/A1/M1/M1/_0_  (.A1(\V4/V1/s1 [0]),
    .A2(\V4/V1/v1 [4]),
    .ZN(\V4/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M1/M1/_1_  (.A(\V4/V1/s1 [0]),
    .B(\V4/V1/v1 [4]),
    .Z(\V4/V1/A2/A1/M1/s1 ));
 AND2_X1 \V4/V1/A2/A1/M1/M2/_0_  (.A1(\V4/V1/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M1/M2/_1_  (.A(\V4/V1/A2/A1/M1/s1 ),
    .B(ground),
    .Z(v4[4]));
 OR2_X1 \V4/V1/A2/A1/M1/_0_  (.A1(\V4/V1/A2/A1/M1/c1 ),
    .A2(\V4/V1/A2/A1/M1/c2 ),
    .ZN(\V4/V1/A2/A1/c1 ));
 AND2_X1 \V4/V1/A2/A1/M2/M1/_0_  (.A1(\V4/V1/s1 [1]),
    .A2(\V4/V1/v1 [5]),
    .ZN(\V4/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M2/M1/_1_  (.A(\V4/V1/s1 [1]),
    .B(\V4/V1/v1 [5]),
    .Z(\V4/V1/A2/A1/M2/s1 ));
 AND2_X1 \V4/V1/A2/A1/M2/M2/_0_  (.A1(\V4/V1/A2/A1/M2/s1 ),
    .A2(\V4/V1/A2/A1/c1 ),
    .ZN(\V4/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M2/M2/_1_  (.A(\V4/V1/A2/A1/M2/s1 ),
    .B(\V4/V1/A2/A1/c1 ),
    .Z(v4[5]));
 OR2_X1 \V4/V1/A2/A1/M2/_0_  (.A1(\V4/V1/A2/A1/M2/c1 ),
    .A2(\V4/V1/A2/A1/M2/c2 ),
    .ZN(\V4/V1/A2/A1/c2 ));
 AND2_X1 \V4/V1/A2/A1/M3/M1/_0_  (.A1(\V4/V1/s1 [2]),
    .A2(\V4/V1/v1 [6]),
    .ZN(\V4/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M3/M1/_1_  (.A(\V4/V1/s1 [2]),
    .B(\V4/V1/v1 [6]),
    .Z(\V4/V1/A2/A1/M3/s1 ));
 AND2_X1 \V4/V1/A2/A1/M3/M2/_0_  (.A1(\V4/V1/A2/A1/M3/s1 ),
    .A2(\V4/V1/A2/A1/c2 ),
    .ZN(\V4/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M3/M2/_1_  (.A(\V4/V1/A2/A1/M3/s1 ),
    .B(\V4/V1/A2/A1/c2 ),
    .Z(v4[6]));
 OR2_X1 \V4/V1/A2/A1/M3/_0_  (.A1(\V4/V1/A2/A1/M3/c1 ),
    .A2(\V4/V1/A2/A1/M3/c2 ),
    .ZN(\V4/V1/A2/A1/c3 ));
 AND2_X1 \V4/V1/A2/A1/M4/M1/_0_  (.A1(\V4/V1/s1 [3]),
    .A2(\V4/V1/v1 [7]),
    .ZN(\V4/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M4/M1/_1_  (.A(\V4/V1/s1 [3]),
    .B(\V4/V1/v1 [7]),
    .Z(\V4/V1/A2/A1/M4/s1 ));
 AND2_X1 \V4/V1/A2/A1/M4/M2/_0_  (.A1(\V4/V1/A2/A1/M4/s1 ),
    .A2(\V4/V1/A2/A1/c3 ),
    .ZN(\V4/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M4/M2/_1_  (.A(\V4/V1/A2/A1/M4/s1 ),
    .B(\V4/V1/A2/A1/c3 ),
    .Z(v4[7]));
 OR2_X1 \V4/V1/A2/A1/M4/_0_  (.A1(\V4/V1/A2/A1/M4/c1 ),
    .A2(\V4/V1/A2/A1/M4/c2 ),
    .ZN(\V4/V1/A2/c1 ));
 AND2_X1 \V4/V1/A2/A2/M1/M1/_0_  (.A1(\V4/V1/s1 [4]),
    .A2(ground),
    .ZN(\V4/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M1/M1/_1_  (.A(\V4/V1/s1 [4]),
    .B(ground),
    .Z(\V4/V1/A2/A2/M1/s1 ));
 AND2_X1 \V4/V1/A2/A2/M1/M2/_0_  (.A1(\V4/V1/A2/A2/M1/s1 ),
    .A2(\V4/V1/A2/c1 ),
    .ZN(\V4/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M1/M2/_1_  (.A(\V4/V1/A2/A2/M1/s1 ),
    .B(\V4/V1/A2/c1 ),
    .Z(\V4/V1/s2 [4]));
 OR2_X1 \V4/V1/A2/A2/M1/_0_  (.A1(\V4/V1/A2/A2/M1/c1 ),
    .A2(\V4/V1/A2/A2/M1/c2 ),
    .ZN(\V4/V1/A2/A2/c1 ));
 AND2_X1 \V4/V1/A2/A2/M2/M1/_0_  (.A1(\V4/V1/s1 [5]),
    .A2(ground),
    .ZN(\V4/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M2/M1/_1_  (.A(\V4/V1/s1 [5]),
    .B(ground),
    .Z(\V4/V1/A2/A2/M2/s1 ));
 AND2_X1 \V4/V1/A2/A2/M2/M2/_0_  (.A1(\V4/V1/A2/A2/M2/s1 ),
    .A2(\V4/V1/A2/A2/c1 ),
    .ZN(\V4/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M2/M2/_1_  (.A(\V4/V1/A2/A2/M2/s1 ),
    .B(\V4/V1/A2/A2/c1 ),
    .Z(\V4/V1/s2 [5]));
 OR2_X1 \V4/V1/A2/A2/M2/_0_  (.A1(\V4/V1/A2/A2/M2/c1 ),
    .A2(\V4/V1/A2/A2/M2/c2 ),
    .ZN(\V4/V1/A2/A2/c2 ));
 AND2_X1 \V4/V1/A2/A2/M3/M1/_0_  (.A1(\V4/V1/s1 [6]),
    .A2(ground),
    .ZN(\V4/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M3/M1/_1_  (.A(\V4/V1/s1 [6]),
    .B(ground),
    .Z(\V4/V1/A2/A2/M3/s1 ));
 AND2_X1 \V4/V1/A2/A2/M3/M2/_0_  (.A1(\V4/V1/A2/A2/M3/s1 ),
    .A2(\V4/V1/A2/A2/c2 ),
    .ZN(\V4/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M3/M2/_1_  (.A(\V4/V1/A2/A2/M3/s1 ),
    .B(\V4/V1/A2/A2/c2 ),
    .Z(\V4/V1/s2 [6]));
 OR2_X1 \V4/V1/A2/A2/M3/_0_  (.A1(\V4/V1/A2/A2/M3/c1 ),
    .A2(\V4/V1/A2/A2/M3/c2 ),
    .ZN(\V4/V1/A2/A2/c3 ));
 AND2_X1 \V4/V1/A2/A2/M4/M1/_0_  (.A1(\V4/V1/s1 [7]),
    .A2(ground),
    .ZN(\V4/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M4/M1/_1_  (.A(\V4/V1/s1 [7]),
    .B(ground),
    .Z(\V4/V1/A2/A2/M4/s1 ));
 AND2_X1 \V4/V1/A2/A2/M4/M2/_0_  (.A1(\V4/V1/A2/A2/M4/s1 ),
    .A2(\V4/V1/A2/A2/c3 ),
    .ZN(\V4/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M4/M2/_1_  (.A(\V4/V1/A2/A2/M4/s1 ),
    .B(\V4/V1/A2/A2/c3 ),
    .Z(\V4/V1/s2 [7]));
 OR2_X1 \V4/V1/A2/A2/M4/_0_  (.A1(\V4/V1/A2/A2/M4/c1 ),
    .A2(\V4/V1/A2/A2/M4/c2 ),
    .ZN(\V4/V1/c2 ));
 AND2_X1 \V4/V1/A3/A1/M1/M1/_0_  (.A1(\V4/V1/v4 [0]),
    .A2(\V4/V1/s2 [4]),
    .ZN(\V4/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M1/M1/_1_  (.A(\V4/V1/v4 [0]),
    .B(\V4/V1/s2 [4]),
    .Z(\V4/V1/A3/A1/M1/s1 ));
 AND2_X1 \V4/V1/A3/A1/M1/M2/_0_  (.A1(\V4/V1/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M1/M2/_1_  (.A(\V4/V1/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v1 [8]));
 OR2_X1 \V4/V1/A3/A1/M1/_0_  (.A1(\V4/V1/A3/A1/M1/c1 ),
    .A2(\V4/V1/A3/A1/M1/c2 ),
    .ZN(\V4/V1/A3/A1/c1 ));
 AND2_X1 \V4/V1/A3/A1/M2/M1/_0_  (.A1(\V4/V1/v4 [1]),
    .A2(\V4/V1/s2 [5]),
    .ZN(\V4/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M2/M1/_1_  (.A(\V4/V1/v4 [1]),
    .B(\V4/V1/s2 [5]),
    .Z(\V4/V1/A3/A1/M2/s1 ));
 AND2_X1 \V4/V1/A3/A1/M2/M2/_0_  (.A1(\V4/V1/A3/A1/M2/s1 ),
    .A2(\V4/V1/A3/A1/c1 ),
    .ZN(\V4/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M2/M2/_1_  (.A(\V4/V1/A3/A1/M2/s1 ),
    .B(\V4/V1/A3/A1/c1 ),
    .Z(\V4/v1 [9]));
 OR2_X1 \V4/V1/A3/A1/M2/_0_  (.A1(\V4/V1/A3/A1/M2/c1 ),
    .A2(\V4/V1/A3/A1/M2/c2 ),
    .ZN(\V4/V1/A3/A1/c2 ));
 AND2_X1 \V4/V1/A3/A1/M3/M1/_0_  (.A1(\V4/V1/v4 [2]),
    .A2(\V4/V1/s2 [6]),
    .ZN(\V4/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M3/M1/_1_  (.A(\V4/V1/v4 [2]),
    .B(\V4/V1/s2 [6]),
    .Z(\V4/V1/A3/A1/M3/s1 ));
 AND2_X1 \V4/V1/A3/A1/M3/M2/_0_  (.A1(\V4/V1/A3/A1/M3/s1 ),
    .A2(\V4/V1/A3/A1/c2 ),
    .ZN(\V4/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M3/M2/_1_  (.A(\V4/V1/A3/A1/M3/s1 ),
    .B(\V4/V1/A3/A1/c2 ),
    .Z(\V4/v1 [10]));
 OR2_X1 \V4/V1/A3/A1/M3/_0_  (.A1(\V4/V1/A3/A1/M3/c1 ),
    .A2(\V4/V1/A3/A1/M3/c2 ),
    .ZN(\V4/V1/A3/A1/c3 ));
 AND2_X1 \V4/V1/A3/A1/M4/M1/_0_  (.A1(\V4/V1/v4 [3]),
    .A2(\V4/V1/s2 [7]),
    .ZN(\V4/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M4/M1/_1_  (.A(\V4/V1/v4 [3]),
    .B(\V4/V1/s2 [7]),
    .Z(\V4/V1/A3/A1/M4/s1 ));
 AND2_X1 \V4/V1/A3/A1/M4/M2/_0_  (.A1(\V4/V1/A3/A1/M4/s1 ),
    .A2(\V4/V1/A3/A1/c3 ),
    .ZN(\V4/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M4/M2/_1_  (.A(\V4/V1/A3/A1/M4/s1 ),
    .B(\V4/V1/A3/A1/c3 ),
    .Z(\V4/v1 [11]));
 OR2_X1 \V4/V1/A3/A1/M4/_0_  (.A1(\V4/V1/A3/A1/M4/c1 ),
    .A2(\V4/V1/A3/A1/M4/c2 ),
    .ZN(\V4/V1/A3/c1 ));
 AND2_X1 \V4/V1/A3/A2/M1/M1/_0_  (.A1(\V4/V1/v4 [4]),
    .A2(\V4/V1/c3 ),
    .ZN(\V4/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M1/M1/_1_  (.A(\V4/V1/v4 [4]),
    .B(\V4/V1/c3 ),
    .Z(\V4/V1/A3/A2/M1/s1 ));
 AND2_X1 \V4/V1/A3/A2/M1/M2/_0_  (.A1(\V4/V1/A3/A2/M1/s1 ),
    .A2(\V4/V1/A3/c1 ),
    .ZN(\V4/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M1/M2/_1_  (.A(\V4/V1/A3/A2/M1/s1 ),
    .B(\V4/V1/A3/c1 ),
    .Z(\V4/v1 [12]));
 OR2_X1 \V4/V1/A3/A2/M1/_0_  (.A1(\V4/V1/A3/A2/M1/c1 ),
    .A2(\V4/V1/A3/A2/M1/c2 ),
    .ZN(\V4/V1/A3/A2/c1 ));
 AND2_X1 \V4/V1/A3/A2/M2/M1/_0_  (.A1(\V4/V1/v4 [5]),
    .A2(ground),
    .ZN(\V4/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M2/M1/_1_  (.A(\V4/V1/v4 [5]),
    .B(ground),
    .Z(\V4/V1/A3/A2/M2/s1 ));
 AND2_X1 \V4/V1/A3/A2/M2/M2/_0_  (.A1(\V4/V1/A3/A2/M2/s1 ),
    .A2(\V4/V1/A3/A2/c1 ),
    .ZN(\V4/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M2/M2/_1_  (.A(\V4/V1/A3/A2/M2/s1 ),
    .B(\V4/V1/A3/A2/c1 ),
    .Z(\V4/v1 [13]));
 OR2_X1 \V4/V1/A3/A2/M2/_0_  (.A1(\V4/V1/A3/A2/M2/c1 ),
    .A2(\V4/V1/A3/A2/M2/c2 ),
    .ZN(\V4/V1/A3/A2/c2 ));
 AND2_X1 \V4/V1/A3/A2/M3/M1/_0_  (.A1(\V4/V1/v4 [6]),
    .A2(ground),
    .ZN(\V4/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M3/M1/_1_  (.A(\V4/V1/v4 [6]),
    .B(ground),
    .Z(\V4/V1/A3/A2/M3/s1 ));
 AND2_X1 \V4/V1/A3/A2/M3/M2/_0_  (.A1(\V4/V1/A3/A2/M3/s1 ),
    .A2(\V4/V1/A3/A2/c2 ),
    .ZN(\V4/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M3/M2/_1_  (.A(\V4/V1/A3/A2/M3/s1 ),
    .B(\V4/V1/A3/A2/c2 ),
    .Z(\V4/v1 [14]));
 OR2_X1 \V4/V1/A3/A2/M3/_0_  (.A1(\V4/V1/A3/A2/M3/c1 ),
    .A2(\V4/V1/A3/A2/M3/c2 ),
    .ZN(\V4/V1/A3/A2/c3 ));
 AND2_X1 \V4/V1/A3/A2/M4/M1/_0_  (.A1(\V4/V1/v4 [7]),
    .A2(ground),
    .ZN(\V4/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M4/M1/_1_  (.A(\V4/V1/v4 [7]),
    .B(ground),
    .Z(\V4/V1/A3/A2/M4/s1 ));
 AND2_X1 \V4/V1/A3/A2/M4/M2/_0_  (.A1(\V4/V1/A3/A2/M4/s1 ),
    .A2(\V4/V1/A3/A2/c3 ),
    .ZN(\V4/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M4/M2/_1_  (.A(\V4/V1/A3/A2/M4/s1 ),
    .B(\V4/V1/A3/A2/c3 ),
    .Z(\V4/v1 [15]));
 OR2_X1 \V4/V1/A3/A2/M4/_0_  (.A1(\V4/V1/A3/A2/M4/c1 ),
    .A2(\V4/V1/A3/A2/M4/c2 ),
    .ZN(\V4/V1/overflow ));
 AND2_X1 \V4/V1/V1/A1/M1/M1/_0_  (.A1(\V4/V1/V1/v2 [0]),
    .A2(\V4/V1/V1/v3 [0]),
    .ZN(\V4/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M1/M1/_1_  (.A(\V4/V1/V1/v2 [0]),
    .B(\V4/V1/V1/v3 [0]),
    .Z(\V4/V1/V1/A1/M1/s1 ));
 AND2_X1 \V4/V1/V1/A1/M1/M2/_0_  (.A1(\V4/V1/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M1/M2/_1_  (.A(\V4/V1/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/V1/s1 [0]));
 OR2_X1 \V4/V1/V1/A1/M1/_0_  (.A1(\V4/V1/V1/A1/M1/c1 ),
    .A2(\V4/V1/V1/A1/M1/c2 ),
    .ZN(\V4/V1/V1/A1/c1 ));
 AND2_X1 \V4/V1/V1/A1/M2/M1/_0_  (.A1(\V4/V1/V1/v2 [1]),
    .A2(\V4/V1/V1/v3 [1]),
    .ZN(\V4/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M2/M1/_1_  (.A(\V4/V1/V1/v2 [1]),
    .B(\V4/V1/V1/v3 [1]),
    .Z(\V4/V1/V1/A1/M2/s1 ));
 AND2_X1 \V4/V1/V1/A1/M2/M2/_0_  (.A1(\V4/V1/V1/A1/M2/s1 ),
    .A2(\V4/V1/V1/A1/c1 ),
    .ZN(\V4/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M2/M2/_1_  (.A(\V4/V1/V1/A1/M2/s1 ),
    .B(\V4/V1/V1/A1/c1 ),
    .Z(\V4/V1/V1/s1 [1]));
 OR2_X1 \V4/V1/V1/A1/M2/_0_  (.A1(\V4/V1/V1/A1/M2/c1 ),
    .A2(\V4/V1/V1/A1/M2/c2 ),
    .ZN(\V4/V1/V1/A1/c2 ));
 AND2_X1 \V4/V1/V1/A1/M3/M1/_0_  (.A1(\V4/V1/V1/v2 [2]),
    .A2(\V4/V1/V1/v3 [2]),
    .ZN(\V4/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M3/M1/_1_  (.A(\V4/V1/V1/v2 [2]),
    .B(\V4/V1/V1/v3 [2]),
    .Z(\V4/V1/V1/A1/M3/s1 ));
 AND2_X1 \V4/V1/V1/A1/M3/M2/_0_  (.A1(\V4/V1/V1/A1/M3/s1 ),
    .A2(\V4/V1/V1/A1/c2 ),
    .ZN(\V4/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M3/M2/_1_  (.A(\V4/V1/V1/A1/M3/s1 ),
    .B(\V4/V1/V1/A1/c2 ),
    .Z(\V4/V1/V1/s1 [2]));
 OR2_X1 \V4/V1/V1/A1/M3/_0_  (.A1(\V4/V1/V1/A1/M3/c1 ),
    .A2(\V4/V1/V1/A1/M3/c2 ),
    .ZN(\V4/V1/V1/A1/c3 ));
 AND2_X1 \V4/V1/V1/A1/M4/M1/_0_  (.A1(\V4/V1/V1/v2 [3]),
    .A2(\V4/V1/V1/v3 [3]),
    .ZN(\V4/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M4/M1/_1_  (.A(\V4/V1/V1/v2 [3]),
    .B(\V4/V1/V1/v3 [3]),
    .Z(\V4/V1/V1/A1/M4/s1 ));
 AND2_X1 \V4/V1/V1/A1/M4/M2/_0_  (.A1(\V4/V1/V1/A1/M4/s1 ),
    .A2(\V4/V1/V1/A1/c3 ),
    .ZN(\V4/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M4/M2/_1_  (.A(\V4/V1/V1/A1/M4/s1 ),
    .B(\V4/V1/V1/A1/c3 ),
    .Z(\V4/V1/V1/s1 [3]));
 OR2_X1 \V4/V1/V1/A1/M4/_0_  (.A1(\V4/V1/V1/A1/M4/c1 ),
    .A2(\V4/V1/V1/A1/M4/c2 ),
    .ZN(\V4/V1/V1/c1 ));
 AND2_X1 \V4/V1/V1/A2/M1/M1/_0_  (.A1(\V4/V1/V1/s1 [0]),
    .A2(\V4/V1/V1/v1 [2]),
    .ZN(\V4/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M1/M1/_1_  (.A(\V4/V1/V1/s1 [0]),
    .B(\V4/V1/V1/v1 [2]),
    .Z(\V4/V1/V1/A2/M1/s1 ));
 AND2_X1 \V4/V1/V1/A2/M1/M2/_0_  (.A1(\V4/V1/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M1/M2/_1_  (.A(\V4/V1/V1/A2/M1/s1 ),
    .B(ground),
    .Z(v4[2]));
 OR2_X1 \V4/V1/V1/A2/M1/_0_  (.A1(\V4/V1/V1/A2/M1/c1 ),
    .A2(\V4/V1/V1/A2/M1/c2 ),
    .ZN(\V4/V1/V1/A2/c1 ));
 AND2_X1 \V4/V1/V1/A2/M2/M1/_0_  (.A1(\V4/V1/V1/s1 [1]),
    .A2(\V4/V1/V1/v1 [3]),
    .ZN(\V4/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M2/M1/_1_  (.A(\V4/V1/V1/s1 [1]),
    .B(\V4/V1/V1/v1 [3]),
    .Z(\V4/V1/V1/A2/M2/s1 ));
 AND2_X1 \V4/V1/V1/A2/M2/M2/_0_  (.A1(\V4/V1/V1/A2/M2/s1 ),
    .A2(\V4/V1/V1/A2/c1 ),
    .ZN(\V4/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M2/M2/_1_  (.A(\V4/V1/V1/A2/M2/s1 ),
    .B(\V4/V1/V1/A2/c1 ),
    .Z(v4[3]));
 OR2_X1 \V4/V1/V1/A2/M2/_0_  (.A1(\V4/V1/V1/A2/M2/c1 ),
    .A2(\V4/V1/V1/A2/M2/c2 ),
    .ZN(\V4/V1/V1/A2/c2 ));
 AND2_X1 \V4/V1/V1/A2/M3/M1/_0_  (.A1(\V4/V1/V1/s1 [2]),
    .A2(ground),
    .ZN(\V4/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M3/M1/_1_  (.A(\V4/V1/V1/s1 [2]),
    .B(ground),
    .Z(\V4/V1/V1/A2/M3/s1 ));
 AND2_X1 \V4/V1/V1/A2/M3/M2/_0_  (.A1(\V4/V1/V1/A2/M3/s1 ),
    .A2(\V4/V1/V1/A2/c2 ),
    .ZN(\V4/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M3/M2/_1_  (.A(\V4/V1/V1/A2/M3/s1 ),
    .B(\V4/V1/V1/A2/c2 ),
    .Z(\V4/V1/V1/s2 [2]));
 OR2_X1 \V4/V1/V1/A2/M3/_0_  (.A1(\V4/V1/V1/A2/M3/c1 ),
    .A2(\V4/V1/V1/A2/M3/c2 ),
    .ZN(\V4/V1/V1/A2/c3 ));
 AND2_X1 \V4/V1/V1/A2/M4/M1/_0_  (.A1(\V4/V1/V1/s1 [3]),
    .A2(ground),
    .ZN(\V4/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M4/M1/_1_  (.A(\V4/V1/V1/s1 [3]),
    .B(ground),
    .Z(\V4/V1/V1/A2/M4/s1 ));
 AND2_X1 \V4/V1/V1/A2/M4/M2/_0_  (.A1(\V4/V1/V1/A2/M4/s1 ),
    .A2(\V4/V1/V1/A2/c3 ),
    .ZN(\V4/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M4/M2/_1_  (.A(\V4/V1/V1/A2/M4/s1 ),
    .B(\V4/V1/V1/A2/c3 ),
    .Z(\V4/V1/V1/s2 [3]));
 OR2_X1 \V4/V1/V1/A2/M4/_0_  (.A1(\V4/V1/V1/A2/M4/c1 ),
    .A2(\V4/V1/V1/A2/M4/c2 ),
    .ZN(\V4/V1/V1/c2 ));
 AND2_X1 \V4/V1/V1/A3/M1/M1/_0_  (.A1(\V4/V1/V1/v4 [0]),
    .A2(\V4/V1/V1/s2 [2]),
    .ZN(\V4/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M1/M1/_1_  (.A(\V4/V1/V1/v4 [0]),
    .B(\V4/V1/V1/s2 [2]),
    .Z(\V4/V1/V1/A3/M1/s1 ));
 AND2_X1 \V4/V1/V1/A3/M1/M2/_0_  (.A1(\V4/V1/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M1/M2/_1_  (.A(\V4/V1/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v1 [4]));
 OR2_X1 \V4/V1/V1/A3/M1/_0_  (.A1(\V4/V1/V1/A3/M1/c1 ),
    .A2(\V4/V1/V1/A3/M1/c2 ),
    .ZN(\V4/V1/V1/A3/c1 ));
 AND2_X1 \V4/V1/V1/A3/M2/M1/_0_  (.A1(\V4/V1/V1/v4 [1]),
    .A2(\V4/V1/V1/s2 [3]),
    .ZN(\V4/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M2/M1/_1_  (.A(\V4/V1/V1/v4 [1]),
    .B(\V4/V1/V1/s2 [3]),
    .Z(\V4/V1/V1/A3/M2/s1 ));
 AND2_X1 \V4/V1/V1/A3/M2/M2/_0_  (.A1(\V4/V1/V1/A3/M2/s1 ),
    .A2(\V4/V1/V1/A3/c1 ),
    .ZN(\V4/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M2/M2/_1_  (.A(\V4/V1/V1/A3/M2/s1 ),
    .B(\V4/V1/V1/A3/c1 ),
    .Z(\V4/V1/v1 [5]));
 OR2_X1 \V4/V1/V1/A3/M2/_0_  (.A1(\V4/V1/V1/A3/M2/c1 ),
    .A2(\V4/V1/V1/A3/M2/c2 ),
    .ZN(\V4/V1/V1/A3/c2 ));
 AND2_X1 \V4/V1/V1/A3/M3/M1/_0_  (.A1(\V4/V1/V1/v4 [2]),
    .A2(\V4/V1/V1/c3 ),
    .ZN(\V4/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M3/M1/_1_  (.A(\V4/V1/V1/v4 [2]),
    .B(\V4/V1/V1/c3 ),
    .Z(\V4/V1/V1/A3/M3/s1 ));
 AND2_X1 \V4/V1/V1/A3/M3/M2/_0_  (.A1(\V4/V1/V1/A3/M3/s1 ),
    .A2(\V4/V1/V1/A3/c2 ),
    .ZN(\V4/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M3/M2/_1_  (.A(\V4/V1/V1/A3/M3/s1 ),
    .B(\V4/V1/V1/A3/c2 ),
    .Z(\V4/V1/v1 [6]));
 OR2_X1 \V4/V1/V1/A3/M3/_0_  (.A1(\V4/V1/V1/A3/M3/c1 ),
    .A2(\V4/V1/V1/A3/M3/c2 ),
    .ZN(\V4/V1/V1/A3/c3 ));
 AND2_X1 \V4/V1/V1/A3/M4/M1/_0_  (.A1(\V4/V1/V1/v4 [3]),
    .A2(ground),
    .ZN(\V4/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M4/M1/_1_  (.A(\V4/V1/V1/v4 [3]),
    .B(ground),
    .Z(\V4/V1/V1/A3/M4/s1 ));
 AND2_X1 \V4/V1/V1/A3/M4/M2/_0_  (.A1(\V4/V1/V1/A3/M4/s1 ),
    .A2(\V4/V1/V1/A3/c3 ),
    .ZN(\V4/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M4/M2/_1_  (.A(\V4/V1/V1/A3/M4/s1 ),
    .B(\V4/V1/V1/A3/c3 ),
    .Z(\V4/V1/v1 [7]));
 OR2_X1 \V4/V1/V1/A3/M4/_0_  (.A1(\V4/V1/V1/A3/M4/c1 ),
    .A2(\V4/V1/V1/A3/M4/c2 ),
    .ZN(\V4/V1/V1/overflow ));
 AND2_X1 \V4/V1/V1/V1/HA1/_0_  (.A1(\V4/V1/V1/V1/w2 ),
    .A2(\V4/V1/V1/V1/w1 ),
    .ZN(\V4/V1/V1/V1/w4 ));
 XOR2_X2 \V4/V1/V1/V1/HA1/_1_  (.A(\V4/V1/V1/V1/w2 ),
    .B(\V4/V1/V1/V1/w1 ),
    .Z(v4[1]));
 AND2_X1 \V4/V1/V1/V1/HA2/_0_  (.A1(\V4/V1/V1/V1/w4 ),
    .A2(\V4/V1/V1/V1/w3 ),
    .ZN(\V4/V1/V1/v1 [3]));
 XOR2_X2 \V4/V1/V1/V1/HA2/_1_  (.A(\V4/V1/V1/V1/w4 ),
    .B(\V4/V1/V1/V1/w3 ),
    .Z(\V4/V1/V1/v1 [2]));
 AND2_X1 \V4/V1/V1/V1/_0_  (.A1(A[16]),
    .A2(B[16]),
    .ZN(v4[0]));
 AND2_X1 \V4/V1/V1/V1/_1_  (.A1(A[16]),
    .A2(B[17]),
    .ZN(\V4/V1/V1/V1/w1 ));
 AND2_X1 \V4/V1/V1/V1/_2_  (.A1(B[16]),
    .A2(A[17]),
    .ZN(\V4/V1/V1/V1/w2 ));
 AND2_X1 \V4/V1/V1/V1/_3_  (.A1(B[17]),
    .A2(A[17]),
    .ZN(\V4/V1/V1/V1/w3 ));
 AND2_X1 \V4/V1/V1/V2/HA1/_0_  (.A1(\V4/V1/V1/V2/w2 ),
    .A2(\V4/V1/V1/V2/w1 ),
    .ZN(\V4/V1/V1/V2/w4 ));
 XOR2_X2 \V4/V1/V1/V2/HA1/_1_  (.A(\V4/V1/V1/V2/w2 ),
    .B(\V4/V1/V1/V2/w1 ),
    .Z(\V4/V1/V1/v2 [1]));
 AND2_X1 \V4/V1/V1/V2/HA2/_0_  (.A1(\V4/V1/V1/V2/w4 ),
    .A2(\V4/V1/V1/V2/w3 ),
    .ZN(\V4/V1/V1/v2 [3]));
 XOR2_X2 \V4/V1/V1/V2/HA2/_1_  (.A(\V4/V1/V1/V2/w4 ),
    .B(\V4/V1/V1/V2/w3 ),
    .Z(\V4/V1/V1/v2 [2]));
 AND2_X1 \V4/V1/V1/V2/_0_  (.A1(A[18]),
    .A2(B[16]),
    .ZN(\V4/V1/V1/v2 [0]));
 AND2_X1 \V4/V1/V1/V2/_1_  (.A1(A[18]),
    .A2(B[17]),
    .ZN(\V4/V1/V1/V2/w1 ));
 AND2_X1 \V4/V1/V1/V2/_2_  (.A1(B[16]),
    .A2(A[19]),
    .ZN(\V4/V1/V1/V2/w2 ));
 AND2_X1 \V4/V1/V1/V2/_3_  (.A1(B[17]),
    .A2(A[19]),
    .ZN(\V4/V1/V1/V2/w3 ));
 AND2_X1 \V4/V1/V1/V3/HA1/_0_  (.A1(\V4/V1/V1/V3/w2 ),
    .A2(\V4/V1/V1/V3/w1 ),
    .ZN(\V4/V1/V1/V3/w4 ));
 XOR2_X2 \V4/V1/V1/V3/HA1/_1_  (.A(\V4/V1/V1/V3/w2 ),
    .B(\V4/V1/V1/V3/w1 ),
    .Z(\V4/V1/V1/v3 [1]));
 AND2_X1 \V4/V1/V1/V3/HA2/_0_  (.A1(\V4/V1/V1/V3/w4 ),
    .A2(\V4/V1/V1/V3/w3 ),
    .ZN(\V4/V1/V1/v3 [3]));
 XOR2_X2 \V4/V1/V1/V3/HA2/_1_  (.A(\V4/V1/V1/V3/w4 ),
    .B(\V4/V1/V1/V3/w3 ),
    .Z(\V4/V1/V1/v3 [2]));
 AND2_X1 \V4/V1/V1/V3/_0_  (.A1(A[16]),
    .A2(B[18]),
    .ZN(\V4/V1/V1/v3 [0]));
 AND2_X1 \V4/V1/V1/V3/_1_  (.A1(A[16]),
    .A2(B[19]),
    .ZN(\V4/V1/V1/V3/w1 ));
 AND2_X1 \V4/V1/V1/V3/_2_  (.A1(B[18]),
    .A2(A[17]),
    .ZN(\V4/V1/V1/V3/w2 ));
 AND2_X1 \V4/V1/V1/V3/_3_  (.A1(B[19]),
    .A2(A[17]),
    .ZN(\V4/V1/V1/V3/w3 ));
 AND2_X1 \V4/V1/V1/V4/HA1/_0_  (.A1(\V4/V1/V1/V4/w2 ),
    .A2(\V4/V1/V1/V4/w1 ),
    .ZN(\V4/V1/V1/V4/w4 ));
 XOR2_X2 \V4/V1/V1/V4/HA1/_1_  (.A(\V4/V1/V1/V4/w2 ),
    .B(\V4/V1/V1/V4/w1 ),
    .Z(\V4/V1/V1/v4 [1]));
 AND2_X1 \V4/V1/V1/V4/HA2/_0_  (.A1(\V4/V1/V1/V4/w4 ),
    .A2(\V4/V1/V1/V4/w3 ),
    .ZN(\V4/V1/V1/v4 [3]));
 XOR2_X2 \V4/V1/V1/V4/HA2/_1_  (.A(\V4/V1/V1/V4/w4 ),
    .B(\V4/V1/V1/V4/w3 ),
    .Z(\V4/V1/V1/v4 [2]));
 AND2_X1 \V4/V1/V1/V4/_0_  (.A1(A[18]),
    .A2(B[18]),
    .ZN(\V4/V1/V1/v4 [0]));
 AND2_X1 \V4/V1/V1/V4/_1_  (.A1(A[18]),
    .A2(B[19]),
    .ZN(\V4/V1/V1/V4/w1 ));
 AND2_X1 \V4/V1/V1/V4/_2_  (.A1(B[18]),
    .A2(A[19]),
    .ZN(\V4/V1/V1/V4/w2 ));
 AND2_X1 \V4/V1/V1/V4/_3_  (.A1(B[19]),
    .A2(A[19]),
    .ZN(\V4/V1/V1/V4/w3 ));
 OR2_X1 \V4/V1/V1/_0_  (.A1(\V4/V1/V1/c1 ),
    .A2(\V4/V1/V1/c2 ),
    .ZN(\V4/V1/V1/c3 ));
 AND2_X1 \V4/V1/V2/A1/M1/M1/_0_  (.A1(\V4/V1/V2/v2 [0]),
    .A2(\V4/V1/V2/v3 [0]),
    .ZN(\V4/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M1/M1/_1_  (.A(\V4/V1/V2/v2 [0]),
    .B(\V4/V1/V2/v3 [0]),
    .Z(\V4/V1/V2/A1/M1/s1 ));
 AND2_X1 \V4/V1/V2/A1/M1/M2/_0_  (.A1(\V4/V1/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M1/M2/_1_  (.A(\V4/V1/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/V2/s1 [0]));
 OR2_X1 \V4/V1/V2/A1/M1/_0_  (.A1(\V4/V1/V2/A1/M1/c1 ),
    .A2(\V4/V1/V2/A1/M1/c2 ),
    .ZN(\V4/V1/V2/A1/c1 ));
 AND2_X1 \V4/V1/V2/A1/M2/M1/_0_  (.A1(\V4/V1/V2/v2 [1]),
    .A2(\V4/V1/V2/v3 [1]),
    .ZN(\V4/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M2/M1/_1_  (.A(\V4/V1/V2/v2 [1]),
    .B(\V4/V1/V2/v3 [1]),
    .Z(\V4/V1/V2/A1/M2/s1 ));
 AND2_X1 \V4/V1/V2/A1/M2/M2/_0_  (.A1(\V4/V1/V2/A1/M2/s1 ),
    .A2(\V4/V1/V2/A1/c1 ),
    .ZN(\V4/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M2/M2/_1_  (.A(\V4/V1/V2/A1/M2/s1 ),
    .B(\V4/V1/V2/A1/c1 ),
    .Z(\V4/V1/V2/s1 [1]));
 OR2_X1 \V4/V1/V2/A1/M2/_0_  (.A1(\V4/V1/V2/A1/M2/c1 ),
    .A2(\V4/V1/V2/A1/M2/c2 ),
    .ZN(\V4/V1/V2/A1/c2 ));
 AND2_X1 \V4/V1/V2/A1/M3/M1/_0_  (.A1(\V4/V1/V2/v2 [2]),
    .A2(\V4/V1/V2/v3 [2]),
    .ZN(\V4/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M3/M1/_1_  (.A(\V4/V1/V2/v2 [2]),
    .B(\V4/V1/V2/v3 [2]),
    .Z(\V4/V1/V2/A1/M3/s1 ));
 AND2_X1 \V4/V1/V2/A1/M3/M2/_0_  (.A1(\V4/V1/V2/A1/M3/s1 ),
    .A2(\V4/V1/V2/A1/c2 ),
    .ZN(\V4/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M3/M2/_1_  (.A(\V4/V1/V2/A1/M3/s1 ),
    .B(\V4/V1/V2/A1/c2 ),
    .Z(\V4/V1/V2/s1 [2]));
 OR2_X1 \V4/V1/V2/A1/M3/_0_  (.A1(\V4/V1/V2/A1/M3/c1 ),
    .A2(\V4/V1/V2/A1/M3/c2 ),
    .ZN(\V4/V1/V2/A1/c3 ));
 AND2_X1 \V4/V1/V2/A1/M4/M1/_0_  (.A1(\V4/V1/V2/v2 [3]),
    .A2(\V4/V1/V2/v3 [3]),
    .ZN(\V4/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M4/M1/_1_  (.A(\V4/V1/V2/v2 [3]),
    .B(\V4/V1/V2/v3 [3]),
    .Z(\V4/V1/V2/A1/M4/s1 ));
 AND2_X1 \V4/V1/V2/A1/M4/M2/_0_  (.A1(\V4/V1/V2/A1/M4/s1 ),
    .A2(\V4/V1/V2/A1/c3 ),
    .ZN(\V4/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M4/M2/_1_  (.A(\V4/V1/V2/A1/M4/s1 ),
    .B(\V4/V1/V2/A1/c3 ),
    .Z(\V4/V1/V2/s1 [3]));
 OR2_X1 \V4/V1/V2/A1/M4/_0_  (.A1(\V4/V1/V2/A1/M4/c1 ),
    .A2(\V4/V1/V2/A1/M4/c2 ),
    .ZN(\V4/V1/V2/c1 ));
 AND2_X1 \V4/V1/V2/A2/M1/M1/_0_  (.A1(\V4/V1/V2/s1 [0]),
    .A2(\V4/V1/V2/v1 [2]),
    .ZN(\V4/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M1/M1/_1_  (.A(\V4/V1/V2/s1 [0]),
    .B(\V4/V1/V2/v1 [2]),
    .Z(\V4/V1/V2/A2/M1/s1 ));
 AND2_X1 \V4/V1/V2/A2/M1/M2/_0_  (.A1(\V4/V1/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M1/M2/_1_  (.A(\V4/V1/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v2 [2]));
 OR2_X1 \V4/V1/V2/A2/M1/_0_  (.A1(\V4/V1/V2/A2/M1/c1 ),
    .A2(\V4/V1/V2/A2/M1/c2 ),
    .ZN(\V4/V1/V2/A2/c1 ));
 AND2_X1 \V4/V1/V2/A2/M2/M1/_0_  (.A1(\V4/V1/V2/s1 [1]),
    .A2(\V4/V1/V2/v1 [3]),
    .ZN(\V4/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M2/M1/_1_  (.A(\V4/V1/V2/s1 [1]),
    .B(\V4/V1/V2/v1 [3]),
    .Z(\V4/V1/V2/A2/M2/s1 ));
 AND2_X1 \V4/V1/V2/A2/M2/M2/_0_  (.A1(\V4/V1/V2/A2/M2/s1 ),
    .A2(\V4/V1/V2/A2/c1 ),
    .ZN(\V4/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M2/M2/_1_  (.A(\V4/V1/V2/A2/M2/s1 ),
    .B(\V4/V1/V2/A2/c1 ),
    .Z(\V4/V1/v2 [3]));
 OR2_X1 \V4/V1/V2/A2/M2/_0_  (.A1(\V4/V1/V2/A2/M2/c1 ),
    .A2(\V4/V1/V2/A2/M2/c2 ),
    .ZN(\V4/V1/V2/A2/c2 ));
 AND2_X1 \V4/V1/V2/A2/M3/M1/_0_  (.A1(\V4/V1/V2/s1 [2]),
    .A2(ground),
    .ZN(\V4/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M3/M1/_1_  (.A(\V4/V1/V2/s1 [2]),
    .B(ground),
    .Z(\V4/V1/V2/A2/M3/s1 ));
 AND2_X1 \V4/V1/V2/A2/M3/M2/_0_  (.A1(\V4/V1/V2/A2/M3/s1 ),
    .A2(\V4/V1/V2/A2/c2 ),
    .ZN(\V4/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M3/M2/_1_  (.A(\V4/V1/V2/A2/M3/s1 ),
    .B(\V4/V1/V2/A2/c2 ),
    .Z(\V4/V1/V2/s2 [2]));
 OR2_X1 \V4/V1/V2/A2/M3/_0_  (.A1(\V4/V1/V2/A2/M3/c1 ),
    .A2(\V4/V1/V2/A2/M3/c2 ),
    .ZN(\V4/V1/V2/A2/c3 ));
 AND2_X1 \V4/V1/V2/A2/M4/M1/_0_  (.A1(\V4/V1/V2/s1 [3]),
    .A2(ground),
    .ZN(\V4/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M4/M1/_1_  (.A(\V4/V1/V2/s1 [3]),
    .B(ground),
    .Z(\V4/V1/V2/A2/M4/s1 ));
 AND2_X1 \V4/V1/V2/A2/M4/M2/_0_  (.A1(\V4/V1/V2/A2/M4/s1 ),
    .A2(\V4/V1/V2/A2/c3 ),
    .ZN(\V4/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M4/M2/_1_  (.A(\V4/V1/V2/A2/M4/s1 ),
    .B(\V4/V1/V2/A2/c3 ),
    .Z(\V4/V1/V2/s2 [3]));
 OR2_X1 \V4/V1/V2/A2/M4/_0_  (.A1(\V4/V1/V2/A2/M4/c1 ),
    .A2(\V4/V1/V2/A2/M4/c2 ),
    .ZN(\V4/V1/V2/c2 ));
 AND2_X1 \V4/V1/V2/A3/M1/M1/_0_  (.A1(\V4/V1/V2/v4 [0]),
    .A2(\V4/V1/V2/s2 [2]),
    .ZN(\V4/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M1/M1/_1_  (.A(\V4/V1/V2/v4 [0]),
    .B(\V4/V1/V2/s2 [2]),
    .Z(\V4/V1/V2/A3/M1/s1 ));
 AND2_X1 \V4/V1/V2/A3/M1/M2/_0_  (.A1(\V4/V1/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M1/M2/_1_  (.A(\V4/V1/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v2 [4]));
 OR2_X1 \V4/V1/V2/A3/M1/_0_  (.A1(\V4/V1/V2/A3/M1/c1 ),
    .A2(\V4/V1/V2/A3/M1/c2 ),
    .ZN(\V4/V1/V2/A3/c1 ));
 AND2_X1 \V4/V1/V2/A3/M2/M1/_0_  (.A1(\V4/V1/V2/v4 [1]),
    .A2(\V4/V1/V2/s2 [3]),
    .ZN(\V4/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M2/M1/_1_  (.A(\V4/V1/V2/v4 [1]),
    .B(\V4/V1/V2/s2 [3]),
    .Z(\V4/V1/V2/A3/M2/s1 ));
 AND2_X1 \V4/V1/V2/A3/M2/M2/_0_  (.A1(\V4/V1/V2/A3/M2/s1 ),
    .A2(\V4/V1/V2/A3/c1 ),
    .ZN(\V4/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M2/M2/_1_  (.A(\V4/V1/V2/A3/M2/s1 ),
    .B(\V4/V1/V2/A3/c1 ),
    .Z(\V4/V1/v2 [5]));
 OR2_X1 \V4/V1/V2/A3/M2/_0_  (.A1(\V4/V1/V2/A3/M2/c1 ),
    .A2(\V4/V1/V2/A3/M2/c2 ),
    .ZN(\V4/V1/V2/A3/c2 ));
 AND2_X1 \V4/V1/V2/A3/M3/M1/_0_  (.A1(\V4/V1/V2/v4 [2]),
    .A2(\V4/V1/V2/c3 ),
    .ZN(\V4/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M3/M1/_1_  (.A(\V4/V1/V2/v4 [2]),
    .B(\V4/V1/V2/c3 ),
    .Z(\V4/V1/V2/A3/M3/s1 ));
 AND2_X1 \V4/V1/V2/A3/M3/M2/_0_  (.A1(\V4/V1/V2/A3/M3/s1 ),
    .A2(\V4/V1/V2/A3/c2 ),
    .ZN(\V4/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M3/M2/_1_  (.A(\V4/V1/V2/A3/M3/s1 ),
    .B(\V4/V1/V2/A3/c2 ),
    .Z(\V4/V1/v2 [6]));
 OR2_X1 \V4/V1/V2/A3/M3/_0_  (.A1(\V4/V1/V2/A3/M3/c1 ),
    .A2(\V4/V1/V2/A3/M3/c2 ),
    .ZN(\V4/V1/V2/A3/c3 ));
 AND2_X1 \V4/V1/V2/A3/M4/M1/_0_  (.A1(\V4/V1/V2/v4 [3]),
    .A2(ground),
    .ZN(\V4/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M4/M1/_1_  (.A(\V4/V1/V2/v4 [3]),
    .B(ground),
    .Z(\V4/V1/V2/A3/M4/s1 ));
 AND2_X1 \V4/V1/V2/A3/M4/M2/_0_  (.A1(\V4/V1/V2/A3/M4/s1 ),
    .A2(\V4/V1/V2/A3/c3 ),
    .ZN(\V4/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M4/M2/_1_  (.A(\V4/V1/V2/A3/M4/s1 ),
    .B(\V4/V1/V2/A3/c3 ),
    .Z(\V4/V1/v2 [7]));
 OR2_X1 \V4/V1/V2/A3/M4/_0_  (.A1(\V4/V1/V2/A3/M4/c1 ),
    .A2(\V4/V1/V2/A3/M4/c2 ),
    .ZN(\V4/V1/V2/overflow ));
 AND2_X1 \V4/V1/V2/V1/HA1/_0_  (.A1(\V4/V1/V2/V1/w2 ),
    .A2(\V4/V1/V2/V1/w1 ),
    .ZN(\V4/V1/V2/V1/w4 ));
 XOR2_X2 \V4/V1/V2/V1/HA1/_1_  (.A(\V4/V1/V2/V1/w2 ),
    .B(\V4/V1/V2/V1/w1 ),
    .Z(\V4/V1/v2 [1]));
 AND2_X1 \V4/V1/V2/V1/HA2/_0_  (.A1(\V4/V1/V2/V1/w4 ),
    .A2(\V4/V1/V2/V1/w3 ),
    .ZN(\V4/V1/V2/v1 [3]));
 XOR2_X2 \V4/V1/V2/V1/HA2/_1_  (.A(\V4/V1/V2/V1/w4 ),
    .B(\V4/V1/V2/V1/w3 ),
    .Z(\V4/V1/V2/v1 [2]));
 AND2_X1 \V4/V1/V2/V1/_0_  (.A1(A[20]),
    .A2(B[16]),
    .ZN(\V4/V1/v2 [0]));
 AND2_X1 \V4/V1/V2/V1/_1_  (.A1(A[20]),
    .A2(B[17]),
    .ZN(\V4/V1/V2/V1/w1 ));
 AND2_X1 \V4/V1/V2/V1/_2_  (.A1(B[16]),
    .A2(A[21]),
    .ZN(\V4/V1/V2/V1/w2 ));
 AND2_X1 \V4/V1/V2/V1/_3_  (.A1(B[17]),
    .A2(A[21]),
    .ZN(\V4/V1/V2/V1/w3 ));
 AND2_X1 \V4/V1/V2/V2/HA1/_0_  (.A1(\V4/V1/V2/V2/w2 ),
    .A2(\V4/V1/V2/V2/w1 ),
    .ZN(\V4/V1/V2/V2/w4 ));
 XOR2_X2 \V4/V1/V2/V2/HA1/_1_  (.A(\V4/V1/V2/V2/w2 ),
    .B(\V4/V1/V2/V2/w1 ),
    .Z(\V4/V1/V2/v2 [1]));
 AND2_X1 \V4/V1/V2/V2/HA2/_0_  (.A1(\V4/V1/V2/V2/w4 ),
    .A2(\V4/V1/V2/V2/w3 ),
    .ZN(\V4/V1/V2/v2 [3]));
 XOR2_X2 \V4/V1/V2/V2/HA2/_1_  (.A(\V4/V1/V2/V2/w4 ),
    .B(\V4/V1/V2/V2/w3 ),
    .Z(\V4/V1/V2/v2 [2]));
 AND2_X1 \V4/V1/V2/V2/_0_  (.A1(A[22]),
    .A2(B[16]),
    .ZN(\V4/V1/V2/v2 [0]));
 AND2_X1 \V4/V1/V2/V2/_1_  (.A1(A[22]),
    .A2(B[17]),
    .ZN(\V4/V1/V2/V2/w1 ));
 AND2_X1 \V4/V1/V2/V2/_2_  (.A1(B[16]),
    .A2(A[23]),
    .ZN(\V4/V1/V2/V2/w2 ));
 AND2_X1 \V4/V1/V2/V2/_3_  (.A1(B[17]),
    .A2(A[23]),
    .ZN(\V4/V1/V2/V2/w3 ));
 AND2_X1 \V4/V1/V2/V3/HA1/_0_  (.A1(\V4/V1/V2/V3/w2 ),
    .A2(\V4/V1/V2/V3/w1 ),
    .ZN(\V4/V1/V2/V3/w4 ));
 XOR2_X2 \V4/V1/V2/V3/HA1/_1_  (.A(\V4/V1/V2/V3/w2 ),
    .B(\V4/V1/V2/V3/w1 ),
    .Z(\V4/V1/V2/v3 [1]));
 AND2_X1 \V4/V1/V2/V3/HA2/_0_  (.A1(\V4/V1/V2/V3/w4 ),
    .A2(\V4/V1/V2/V3/w3 ),
    .ZN(\V4/V1/V2/v3 [3]));
 XOR2_X2 \V4/V1/V2/V3/HA2/_1_  (.A(\V4/V1/V2/V3/w4 ),
    .B(\V4/V1/V2/V3/w3 ),
    .Z(\V4/V1/V2/v3 [2]));
 AND2_X1 \V4/V1/V2/V3/_0_  (.A1(A[20]),
    .A2(B[18]),
    .ZN(\V4/V1/V2/v3 [0]));
 AND2_X1 \V4/V1/V2/V3/_1_  (.A1(A[20]),
    .A2(B[19]),
    .ZN(\V4/V1/V2/V3/w1 ));
 AND2_X1 \V4/V1/V2/V3/_2_  (.A1(B[18]),
    .A2(A[21]),
    .ZN(\V4/V1/V2/V3/w2 ));
 AND2_X1 \V4/V1/V2/V3/_3_  (.A1(B[19]),
    .A2(A[21]),
    .ZN(\V4/V1/V2/V3/w3 ));
 AND2_X1 \V4/V1/V2/V4/HA1/_0_  (.A1(\V4/V1/V2/V4/w2 ),
    .A2(\V4/V1/V2/V4/w1 ),
    .ZN(\V4/V1/V2/V4/w4 ));
 XOR2_X2 \V4/V1/V2/V4/HA1/_1_  (.A(\V4/V1/V2/V4/w2 ),
    .B(\V4/V1/V2/V4/w1 ),
    .Z(\V4/V1/V2/v4 [1]));
 AND2_X1 \V4/V1/V2/V4/HA2/_0_  (.A1(\V4/V1/V2/V4/w4 ),
    .A2(\V4/V1/V2/V4/w3 ),
    .ZN(\V4/V1/V2/v4 [3]));
 XOR2_X2 \V4/V1/V2/V4/HA2/_1_  (.A(\V4/V1/V2/V4/w4 ),
    .B(\V4/V1/V2/V4/w3 ),
    .Z(\V4/V1/V2/v4 [2]));
 AND2_X1 \V4/V1/V2/V4/_0_  (.A1(A[22]),
    .A2(B[18]),
    .ZN(\V4/V1/V2/v4 [0]));
 AND2_X1 \V4/V1/V2/V4/_1_  (.A1(A[22]),
    .A2(B[19]),
    .ZN(\V4/V1/V2/V4/w1 ));
 AND2_X1 \V4/V1/V2/V4/_2_  (.A1(B[18]),
    .A2(A[23]),
    .ZN(\V4/V1/V2/V4/w2 ));
 AND2_X1 \V4/V1/V2/V4/_3_  (.A1(B[19]),
    .A2(A[23]),
    .ZN(\V4/V1/V2/V4/w3 ));
 OR2_X1 \V4/V1/V2/_0_  (.A1(\V4/V1/V2/c1 ),
    .A2(\V4/V1/V2/c2 ),
    .ZN(\V4/V1/V2/c3 ));
 AND2_X1 \V4/V1/V3/A1/M1/M1/_0_  (.A1(\V4/V1/V3/v2 [0]),
    .A2(\V4/V1/V3/v3 [0]),
    .ZN(\V4/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M1/M1/_1_  (.A(\V4/V1/V3/v2 [0]),
    .B(\V4/V1/V3/v3 [0]),
    .Z(\V4/V1/V3/A1/M1/s1 ));
 AND2_X1 \V4/V1/V3/A1/M1/M2/_0_  (.A1(\V4/V1/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M1/M2/_1_  (.A(\V4/V1/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/V3/s1 [0]));
 OR2_X1 \V4/V1/V3/A1/M1/_0_  (.A1(\V4/V1/V3/A1/M1/c1 ),
    .A2(\V4/V1/V3/A1/M1/c2 ),
    .ZN(\V4/V1/V3/A1/c1 ));
 AND2_X1 \V4/V1/V3/A1/M2/M1/_0_  (.A1(\V4/V1/V3/v2 [1]),
    .A2(\V4/V1/V3/v3 [1]),
    .ZN(\V4/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M2/M1/_1_  (.A(\V4/V1/V3/v2 [1]),
    .B(\V4/V1/V3/v3 [1]),
    .Z(\V4/V1/V3/A1/M2/s1 ));
 AND2_X1 \V4/V1/V3/A1/M2/M2/_0_  (.A1(\V4/V1/V3/A1/M2/s1 ),
    .A2(\V4/V1/V3/A1/c1 ),
    .ZN(\V4/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M2/M2/_1_  (.A(\V4/V1/V3/A1/M2/s1 ),
    .B(\V4/V1/V3/A1/c1 ),
    .Z(\V4/V1/V3/s1 [1]));
 OR2_X1 \V4/V1/V3/A1/M2/_0_  (.A1(\V4/V1/V3/A1/M2/c1 ),
    .A2(\V4/V1/V3/A1/M2/c2 ),
    .ZN(\V4/V1/V3/A1/c2 ));
 AND2_X1 \V4/V1/V3/A1/M3/M1/_0_  (.A1(\V4/V1/V3/v2 [2]),
    .A2(\V4/V1/V3/v3 [2]),
    .ZN(\V4/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M3/M1/_1_  (.A(\V4/V1/V3/v2 [2]),
    .B(\V4/V1/V3/v3 [2]),
    .Z(\V4/V1/V3/A1/M3/s1 ));
 AND2_X1 \V4/V1/V3/A1/M3/M2/_0_  (.A1(\V4/V1/V3/A1/M3/s1 ),
    .A2(\V4/V1/V3/A1/c2 ),
    .ZN(\V4/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M3/M2/_1_  (.A(\V4/V1/V3/A1/M3/s1 ),
    .B(\V4/V1/V3/A1/c2 ),
    .Z(\V4/V1/V3/s1 [2]));
 OR2_X1 \V4/V1/V3/A1/M3/_0_  (.A1(\V4/V1/V3/A1/M3/c1 ),
    .A2(\V4/V1/V3/A1/M3/c2 ),
    .ZN(\V4/V1/V3/A1/c3 ));
 AND2_X1 \V4/V1/V3/A1/M4/M1/_0_  (.A1(\V4/V1/V3/v2 [3]),
    .A2(\V4/V1/V3/v3 [3]),
    .ZN(\V4/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M4/M1/_1_  (.A(\V4/V1/V3/v2 [3]),
    .B(\V4/V1/V3/v3 [3]),
    .Z(\V4/V1/V3/A1/M4/s1 ));
 AND2_X1 \V4/V1/V3/A1/M4/M2/_0_  (.A1(\V4/V1/V3/A1/M4/s1 ),
    .A2(\V4/V1/V3/A1/c3 ),
    .ZN(\V4/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M4/M2/_1_  (.A(\V4/V1/V3/A1/M4/s1 ),
    .B(\V4/V1/V3/A1/c3 ),
    .Z(\V4/V1/V3/s1 [3]));
 OR2_X1 \V4/V1/V3/A1/M4/_0_  (.A1(\V4/V1/V3/A1/M4/c1 ),
    .A2(\V4/V1/V3/A1/M4/c2 ),
    .ZN(\V4/V1/V3/c1 ));
 AND2_X1 \V4/V1/V3/A2/M1/M1/_0_  (.A1(\V4/V1/V3/s1 [0]),
    .A2(\V4/V1/V3/v1 [2]),
    .ZN(\V4/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M1/M1/_1_  (.A(\V4/V1/V3/s1 [0]),
    .B(\V4/V1/V3/v1 [2]),
    .Z(\V4/V1/V3/A2/M1/s1 ));
 AND2_X1 \V4/V1/V3/A2/M1/M2/_0_  (.A1(\V4/V1/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M1/M2/_1_  (.A(\V4/V1/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v3 [2]));
 OR2_X1 \V4/V1/V3/A2/M1/_0_  (.A1(\V4/V1/V3/A2/M1/c1 ),
    .A2(\V4/V1/V3/A2/M1/c2 ),
    .ZN(\V4/V1/V3/A2/c1 ));
 AND2_X1 \V4/V1/V3/A2/M2/M1/_0_  (.A1(\V4/V1/V3/s1 [1]),
    .A2(\V4/V1/V3/v1 [3]),
    .ZN(\V4/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M2/M1/_1_  (.A(\V4/V1/V3/s1 [1]),
    .B(\V4/V1/V3/v1 [3]),
    .Z(\V4/V1/V3/A2/M2/s1 ));
 AND2_X1 \V4/V1/V3/A2/M2/M2/_0_  (.A1(\V4/V1/V3/A2/M2/s1 ),
    .A2(\V4/V1/V3/A2/c1 ),
    .ZN(\V4/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M2/M2/_1_  (.A(\V4/V1/V3/A2/M2/s1 ),
    .B(\V4/V1/V3/A2/c1 ),
    .Z(\V4/V1/v3 [3]));
 OR2_X1 \V4/V1/V3/A2/M2/_0_  (.A1(\V4/V1/V3/A2/M2/c1 ),
    .A2(\V4/V1/V3/A2/M2/c2 ),
    .ZN(\V4/V1/V3/A2/c2 ));
 AND2_X1 \V4/V1/V3/A2/M3/M1/_0_  (.A1(\V4/V1/V3/s1 [2]),
    .A2(ground),
    .ZN(\V4/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M3/M1/_1_  (.A(\V4/V1/V3/s1 [2]),
    .B(ground),
    .Z(\V4/V1/V3/A2/M3/s1 ));
 AND2_X1 \V4/V1/V3/A2/M3/M2/_0_  (.A1(\V4/V1/V3/A2/M3/s1 ),
    .A2(\V4/V1/V3/A2/c2 ),
    .ZN(\V4/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M3/M2/_1_  (.A(\V4/V1/V3/A2/M3/s1 ),
    .B(\V4/V1/V3/A2/c2 ),
    .Z(\V4/V1/V3/s2 [2]));
 OR2_X1 \V4/V1/V3/A2/M3/_0_  (.A1(\V4/V1/V3/A2/M3/c1 ),
    .A2(\V4/V1/V3/A2/M3/c2 ),
    .ZN(\V4/V1/V3/A2/c3 ));
 AND2_X1 \V4/V1/V3/A2/M4/M1/_0_  (.A1(\V4/V1/V3/s1 [3]),
    .A2(ground),
    .ZN(\V4/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M4/M1/_1_  (.A(\V4/V1/V3/s1 [3]),
    .B(ground),
    .Z(\V4/V1/V3/A2/M4/s1 ));
 AND2_X1 \V4/V1/V3/A2/M4/M2/_0_  (.A1(\V4/V1/V3/A2/M4/s1 ),
    .A2(\V4/V1/V3/A2/c3 ),
    .ZN(\V4/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M4/M2/_1_  (.A(\V4/V1/V3/A2/M4/s1 ),
    .B(\V4/V1/V3/A2/c3 ),
    .Z(\V4/V1/V3/s2 [3]));
 OR2_X1 \V4/V1/V3/A2/M4/_0_  (.A1(\V4/V1/V3/A2/M4/c1 ),
    .A2(\V4/V1/V3/A2/M4/c2 ),
    .ZN(\V4/V1/V3/c2 ));
 AND2_X1 \V4/V1/V3/A3/M1/M1/_0_  (.A1(\V4/V1/V3/v4 [0]),
    .A2(\V4/V1/V3/s2 [2]),
    .ZN(\V4/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M1/M1/_1_  (.A(\V4/V1/V3/v4 [0]),
    .B(\V4/V1/V3/s2 [2]),
    .Z(\V4/V1/V3/A3/M1/s1 ));
 AND2_X1 \V4/V1/V3/A3/M1/M2/_0_  (.A1(\V4/V1/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M1/M2/_1_  (.A(\V4/V1/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v3 [4]));
 OR2_X1 \V4/V1/V3/A3/M1/_0_  (.A1(\V4/V1/V3/A3/M1/c1 ),
    .A2(\V4/V1/V3/A3/M1/c2 ),
    .ZN(\V4/V1/V3/A3/c1 ));
 AND2_X1 \V4/V1/V3/A3/M2/M1/_0_  (.A1(\V4/V1/V3/v4 [1]),
    .A2(\V4/V1/V3/s2 [3]),
    .ZN(\V4/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M2/M1/_1_  (.A(\V4/V1/V3/v4 [1]),
    .B(\V4/V1/V3/s2 [3]),
    .Z(\V4/V1/V3/A3/M2/s1 ));
 AND2_X1 \V4/V1/V3/A3/M2/M2/_0_  (.A1(\V4/V1/V3/A3/M2/s1 ),
    .A2(\V4/V1/V3/A3/c1 ),
    .ZN(\V4/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M2/M2/_1_  (.A(\V4/V1/V3/A3/M2/s1 ),
    .B(\V4/V1/V3/A3/c1 ),
    .Z(\V4/V1/v3 [5]));
 OR2_X1 \V4/V1/V3/A3/M2/_0_  (.A1(\V4/V1/V3/A3/M2/c1 ),
    .A2(\V4/V1/V3/A3/M2/c2 ),
    .ZN(\V4/V1/V3/A3/c2 ));
 AND2_X1 \V4/V1/V3/A3/M3/M1/_0_  (.A1(\V4/V1/V3/v4 [2]),
    .A2(\V4/V1/V3/c3 ),
    .ZN(\V4/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M3/M1/_1_  (.A(\V4/V1/V3/v4 [2]),
    .B(\V4/V1/V3/c3 ),
    .Z(\V4/V1/V3/A3/M3/s1 ));
 AND2_X1 \V4/V1/V3/A3/M3/M2/_0_  (.A1(\V4/V1/V3/A3/M3/s1 ),
    .A2(\V4/V1/V3/A3/c2 ),
    .ZN(\V4/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M3/M2/_1_  (.A(\V4/V1/V3/A3/M3/s1 ),
    .B(\V4/V1/V3/A3/c2 ),
    .Z(\V4/V1/v3 [6]));
 OR2_X1 \V4/V1/V3/A3/M3/_0_  (.A1(\V4/V1/V3/A3/M3/c1 ),
    .A2(\V4/V1/V3/A3/M3/c2 ),
    .ZN(\V4/V1/V3/A3/c3 ));
 AND2_X1 \V4/V1/V3/A3/M4/M1/_0_  (.A1(\V4/V1/V3/v4 [3]),
    .A2(ground),
    .ZN(\V4/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M4/M1/_1_  (.A(\V4/V1/V3/v4 [3]),
    .B(ground),
    .Z(\V4/V1/V3/A3/M4/s1 ));
 AND2_X1 \V4/V1/V3/A3/M4/M2/_0_  (.A1(\V4/V1/V3/A3/M4/s1 ),
    .A2(\V4/V1/V3/A3/c3 ),
    .ZN(\V4/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M4/M2/_1_  (.A(\V4/V1/V3/A3/M4/s1 ),
    .B(\V4/V1/V3/A3/c3 ),
    .Z(\V4/V1/v3 [7]));
 OR2_X1 \V4/V1/V3/A3/M4/_0_  (.A1(\V4/V1/V3/A3/M4/c1 ),
    .A2(\V4/V1/V3/A3/M4/c2 ),
    .ZN(\V4/V1/V3/overflow ));
 AND2_X1 \V4/V1/V3/V1/HA1/_0_  (.A1(\V4/V1/V3/V1/w2 ),
    .A2(\V4/V1/V3/V1/w1 ),
    .ZN(\V4/V1/V3/V1/w4 ));
 XOR2_X2 \V4/V1/V3/V1/HA1/_1_  (.A(\V4/V1/V3/V1/w2 ),
    .B(\V4/V1/V3/V1/w1 ),
    .Z(\V4/V1/v3 [1]));
 AND2_X1 \V4/V1/V3/V1/HA2/_0_  (.A1(\V4/V1/V3/V1/w4 ),
    .A2(\V4/V1/V3/V1/w3 ),
    .ZN(\V4/V1/V3/v1 [3]));
 XOR2_X2 \V4/V1/V3/V1/HA2/_1_  (.A(\V4/V1/V3/V1/w4 ),
    .B(\V4/V1/V3/V1/w3 ),
    .Z(\V4/V1/V3/v1 [2]));
 AND2_X1 \V4/V1/V3/V1/_0_  (.A1(A[16]),
    .A2(B[20]),
    .ZN(\V4/V1/v3 [0]));
 AND2_X1 \V4/V1/V3/V1/_1_  (.A1(A[16]),
    .A2(B[21]),
    .ZN(\V4/V1/V3/V1/w1 ));
 AND2_X1 \V4/V1/V3/V1/_2_  (.A1(B[20]),
    .A2(A[17]),
    .ZN(\V4/V1/V3/V1/w2 ));
 AND2_X1 \V4/V1/V3/V1/_3_  (.A1(B[21]),
    .A2(A[17]),
    .ZN(\V4/V1/V3/V1/w3 ));
 AND2_X1 \V4/V1/V3/V2/HA1/_0_  (.A1(\V4/V1/V3/V2/w2 ),
    .A2(\V4/V1/V3/V2/w1 ),
    .ZN(\V4/V1/V3/V2/w4 ));
 XOR2_X2 \V4/V1/V3/V2/HA1/_1_  (.A(\V4/V1/V3/V2/w2 ),
    .B(\V4/V1/V3/V2/w1 ),
    .Z(\V4/V1/V3/v2 [1]));
 AND2_X1 \V4/V1/V3/V2/HA2/_0_  (.A1(\V4/V1/V3/V2/w4 ),
    .A2(\V4/V1/V3/V2/w3 ),
    .ZN(\V4/V1/V3/v2 [3]));
 XOR2_X2 \V4/V1/V3/V2/HA2/_1_  (.A(\V4/V1/V3/V2/w4 ),
    .B(\V4/V1/V3/V2/w3 ),
    .Z(\V4/V1/V3/v2 [2]));
 AND2_X1 \V4/V1/V3/V2/_0_  (.A1(A[18]),
    .A2(B[20]),
    .ZN(\V4/V1/V3/v2 [0]));
 AND2_X1 \V4/V1/V3/V2/_1_  (.A1(A[18]),
    .A2(B[21]),
    .ZN(\V4/V1/V3/V2/w1 ));
 AND2_X1 \V4/V1/V3/V2/_2_  (.A1(B[20]),
    .A2(A[19]),
    .ZN(\V4/V1/V3/V2/w2 ));
 AND2_X1 \V4/V1/V3/V2/_3_  (.A1(B[21]),
    .A2(A[19]),
    .ZN(\V4/V1/V3/V2/w3 ));
 AND2_X1 \V4/V1/V3/V3/HA1/_0_  (.A1(\V4/V1/V3/V3/w2 ),
    .A2(\V4/V1/V3/V3/w1 ),
    .ZN(\V4/V1/V3/V3/w4 ));
 XOR2_X2 \V4/V1/V3/V3/HA1/_1_  (.A(\V4/V1/V3/V3/w2 ),
    .B(\V4/V1/V3/V3/w1 ),
    .Z(\V4/V1/V3/v3 [1]));
 AND2_X1 \V4/V1/V3/V3/HA2/_0_  (.A1(\V4/V1/V3/V3/w4 ),
    .A2(\V4/V1/V3/V3/w3 ),
    .ZN(\V4/V1/V3/v3 [3]));
 XOR2_X2 \V4/V1/V3/V3/HA2/_1_  (.A(\V4/V1/V3/V3/w4 ),
    .B(\V4/V1/V3/V3/w3 ),
    .Z(\V4/V1/V3/v3 [2]));
 AND2_X1 \V4/V1/V3/V3/_0_  (.A1(A[16]),
    .A2(B[22]),
    .ZN(\V4/V1/V3/v3 [0]));
 AND2_X1 \V4/V1/V3/V3/_1_  (.A1(A[16]),
    .A2(B[23]),
    .ZN(\V4/V1/V3/V3/w1 ));
 AND2_X1 \V4/V1/V3/V3/_2_  (.A1(B[22]),
    .A2(A[17]),
    .ZN(\V4/V1/V3/V3/w2 ));
 AND2_X1 \V4/V1/V3/V3/_3_  (.A1(B[23]),
    .A2(A[17]),
    .ZN(\V4/V1/V3/V3/w3 ));
 AND2_X1 \V4/V1/V3/V4/HA1/_0_  (.A1(\V4/V1/V3/V4/w2 ),
    .A2(\V4/V1/V3/V4/w1 ),
    .ZN(\V4/V1/V3/V4/w4 ));
 XOR2_X2 \V4/V1/V3/V4/HA1/_1_  (.A(\V4/V1/V3/V4/w2 ),
    .B(\V4/V1/V3/V4/w1 ),
    .Z(\V4/V1/V3/v4 [1]));
 AND2_X1 \V4/V1/V3/V4/HA2/_0_  (.A1(\V4/V1/V3/V4/w4 ),
    .A2(\V4/V1/V3/V4/w3 ),
    .ZN(\V4/V1/V3/v4 [3]));
 XOR2_X2 \V4/V1/V3/V4/HA2/_1_  (.A(\V4/V1/V3/V4/w4 ),
    .B(\V4/V1/V3/V4/w3 ),
    .Z(\V4/V1/V3/v4 [2]));
 AND2_X1 \V4/V1/V3/V4/_0_  (.A1(A[18]),
    .A2(B[22]),
    .ZN(\V4/V1/V3/v4 [0]));
 AND2_X1 \V4/V1/V3/V4/_1_  (.A1(A[18]),
    .A2(B[23]),
    .ZN(\V4/V1/V3/V4/w1 ));
 AND2_X1 \V4/V1/V3/V4/_2_  (.A1(B[22]),
    .A2(A[19]),
    .ZN(\V4/V1/V3/V4/w2 ));
 AND2_X1 \V4/V1/V3/V4/_3_  (.A1(B[23]),
    .A2(A[19]),
    .ZN(\V4/V1/V3/V4/w3 ));
 OR2_X1 \V4/V1/V3/_0_  (.A1(\V4/V1/V3/c1 ),
    .A2(\V4/V1/V3/c2 ),
    .ZN(\V4/V1/V3/c3 ));
 AND2_X1 \V4/V1/V4/A1/M1/M1/_0_  (.A1(\V4/V1/V4/v2 [0]),
    .A2(\V4/V1/V4/v3 [0]),
    .ZN(\V4/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M1/M1/_1_  (.A(\V4/V1/V4/v2 [0]),
    .B(\V4/V1/V4/v3 [0]),
    .Z(\V4/V1/V4/A1/M1/s1 ));
 AND2_X1 \V4/V1/V4/A1/M1/M2/_0_  (.A1(\V4/V1/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M1/M2/_1_  (.A(\V4/V1/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/V4/s1 [0]));
 OR2_X1 \V4/V1/V4/A1/M1/_0_  (.A1(\V4/V1/V4/A1/M1/c1 ),
    .A2(\V4/V1/V4/A1/M1/c2 ),
    .ZN(\V4/V1/V4/A1/c1 ));
 AND2_X1 \V4/V1/V4/A1/M2/M1/_0_  (.A1(\V4/V1/V4/v2 [1]),
    .A2(\V4/V1/V4/v3 [1]),
    .ZN(\V4/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M2/M1/_1_  (.A(\V4/V1/V4/v2 [1]),
    .B(\V4/V1/V4/v3 [1]),
    .Z(\V4/V1/V4/A1/M2/s1 ));
 AND2_X1 \V4/V1/V4/A1/M2/M2/_0_  (.A1(\V4/V1/V4/A1/M2/s1 ),
    .A2(\V4/V1/V4/A1/c1 ),
    .ZN(\V4/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M2/M2/_1_  (.A(\V4/V1/V4/A1/M2/s1 ),
    .B(\V4/V1/V4/A1/c1 ),
    .Z(\V4/V1/V4/s1 [1]));
 OR2_X1 \V4/V1/V4/A1/M2/_0_  (.A1(\V4/V1/V4/A1/M2/c1 ),
    .A2(\V4/V1/V4/A1/M2/c2 ),
    .ZN(\V4/V1/V4/A1/c2 ));
 AND2_X1 \V4/V1/V4/A1/M3/M1/_0_  (.A1(\V4/V1/V4/v2 [2]),
    .A2(\V4/V1/V4/v3 [2]),
    .ZN(\V4/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M3/M1/_1_  (.A(\V4/V1/V4/v2 [2]),
    .B(\V4/V1/V4/v3 [2]),
    .Z(\V4/V1/V4/A1/M3/s1 ));
 AND2_X1 \V4/V1/V4/A1/M3/M2/_0_  (.A1(\V4/V1/V4/A1/M3/s1 ),
    .A2(\V4/V1/V4/A1/c2 ),
    .ZN(\V4/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M3/M2/_1_  (.A(\V4/V1/V4/A1/M3/s1 ),
    .B(\V4/V1/V4/A1/c2 ),
    .Z(\V4/V1/V4/s1 [2]));
 OR2_X1 \V4/V1/V4/A1/M3/_0_  (.A1(\V4/V1/V4/A1/M3/c1 ),
    .A2(\V4/V1/V4/A1/M3/c2 ),
    .ZN(\V4/V1/V4/A1/c3 ));
 AND2_X1 \V4/V1/V4/A1/M4/M1/_0_  (.A1(\V4/V1/V4/v2 [3]),
    .A2(\V4/V1/V4/v3 [3]),
    .ZN(\V4/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M4/M1/_1_  (.A(\V4/V1/V4/v2 [3]),
    .B(\V4/V1/V4/v3 [3]),
    .Z(\V4/V1/V4/A1/M4/s1 ));
 AND2_X1 \V4/V1/V4/A1/M4/M2/_0_  (.A1(\V4/V1/V4/A1/M4/s1 ),
    .A2(\V4/V1/V4/A1/c3 ),
    .ZN(\V4/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M4/M2/_1_  (.A(\V4/V1/V4/A1/M4/s1 ),
    .B(\V4/V1/V4/A1/c3 ),
    .Z(\V4/V1/V4/s1 [3]));
 OR2_X1 \V4/V1/V4/A1/M4/_0_  (.A1(\V4/V1/V4/A1/M4/c1 ),
    .A2(\V4/V1/V4/A1/M4/c2 ),
    .ZN(\V4/V1/V4/c1 ));
 AND2_X1 \V4/V1/V4/A2/M1/M1/_0_  (.A1(\V4/V1/V4/s1 [0]),
    .A2(\V4/V1/V4/v1 [2]),
    .ZN(\V4/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M1/M1/_1_  (.A(\V4/V1/V4/s1 [0]),
    .B(\V4/V1/V4/v1 [2]),
    .Z(\V4/V1/V4/A2/M1/s1 ));
 AND2_X1 \V4/V1/V4/A2/M1/M2/_0_  (.A1(\V4/V1/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M1/M2/_1_  (.A(\V4/V1/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v4 [2]));
 OR2_X1 \V4/V1/V4/A2/M1/_0_  (.A1(\V4/V1/V4/A2/M1/c1 ),
    .A2(\V4/V1/V4/A2/M1/c2 ),
    .ZN(\V4/V1/V4/A2/c1 ));
 AND2_X1 \V4/V1/V4/A2/M2/M1/_0_  (.A1(\V4/V1/V4/s1 [1]),
    .A2(\V4/V1/V4/v1 [3]),
    .ZN(\V4/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M2/M1/_1_  (.A(\V4/V1/V4/s1 [1]),
    .B(\V4/V1/V4/v1 [3]),
    .Z(\V4/V1/V4/A2/M2/s1 ));
 AND2_X1 \V4/V1/V4/A2/M2/M2/_0_  (.A1(\V4/V1/V4/A2/M2/s1 ),
    .A2(\V4/V1/V4/A2/c1 ),
    .ZN(\V4/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M2/M2/_1_  (.A(\V4/V1/V4/A2/M2/s1 ),
    .B(\V4/V1/V4/A2/c1 ),
    .Z(\V4/V1/v4 [3]));
 OR2_X1 \V4/V1/V4/A2/M2/_0_  (.A1(\V4/V1/V4/A2/M2/c1 ),
    .A2(\V4/V1/V4/A2/M2/c2 ),
    .ZN(\V4/V1/V4/A2/c2 ));
 AND2_X1 \V4/V1/V4/A2/M3/M1/_0_  (.A1(\V4/V1/V4/s1 [2]),
    .A2(ground),
    .ZN(\V4/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M3/M1/_1_  (.A(\V4/V1/V4/s1 [2]),
    .B(ground),
    .Z(\V4/V1/V4/A2/M3/s1 ));
 AND2_X1 \V4/V1/V4/A2/M3/M2/_0_  (.A1(\V4/V1/V4/A2/M3/s1 ),
    .A2(\V4/V1/V4/A2/c2 ),
    .ZN(\V4/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M3/M2/_1_  (.A(\V4/V1/V4/A2/M3/s1 ),
    .B(\V4/V1/V4/A2/c2 ),
    .Z(\V4/V1/V4/s2 [2]));
 OR2_X1 \V4/V1/V4/A2/M3/_0_  (.A1(\V4/V1/V4/A2/M3/c1 ),
    .A2(\V4/V1/V4/A2/M3/c2 ),
    .ZN(\V4/V1/V4/A2/c3 ));
 AND2_X1 \V4/V1/V4/A2/M4/M1/_0_  (.A1(\V4/V1/V4/s1 [3]),
    .A2(ground),
    .ZN(\V4/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M4/M1/_1_  (.A(\V4/V1/V4/s1 [3]),
    .B(ground),
    .Z(\V4/V1/V4/A2/M4/s1 ));
 AND2_X1 \V4/V1/V4/A2/M4/M2/_0_  (.A1(\V4/V1/V4/A2/M4/s1 ),
    .A2(\V4/V1/V4/A2/c3 ),
    .ZN(\V4/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M4/M2/_1_  (.A(\V4/V1/V4/A2/M4/s1 ),
    .B(\V4/V1/V4/A2/c3 ),
    .Z(\V4/V1/V4/s2 [3]));
 OR2_X1 \V4/V1/V4/A2/M4/_0_  (.A1(\V4/V1/V4/A2/M4/c1 ),
    .A2(\V4/V1/V4/A2/M4/c2 ),
    .ZN(\V4/V1/V4/c2 ));
 AND2_X1 \V4/V1/V4/A3/M1/M1/_0_  (.A1(\V4/V1/V4/v4 [0]),
    .A2(\V4/V1/V4/s2 [2]),
    .ZN(\V4/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M1/M1/_1_  (.A(\V4/V1/V4/v4 [0]),
    .B(\V4/V1/V4/s2 [2]),
    .Z(\V4/V1/V4/A3/M1/s1 ));
 AND2_X1 \V4/V1/V4/A3/M1/M2/_0_  (.A1(\V4/V1/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M1/M2/_1_  (.A(\V4/V1/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V1/v4 [4]));
 OR2_X1 \V4/V1/V4/A3/M1/_0_  (.A1(\V4/V1/V4/A3/M1/c1 ),
    .A2(\V4/V1/V4/A3/M1/c2 ),
    .ZN(\V4/V1/V4/A3/c1 ));
 AND2_X1 \V4/V1/V4/A3/M2/M1/_0_  (.A1(\V4/V1/V4/v4 [1]),
    .A2(\V4/V1/V4/s2 [3]),
    .ZN(\V4/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M2/M1/_1_  (.A(\V4/V1/V4/v4 [1]),
    .B(\V4/V1/V4/s2 [3]),
    .Z(\V4/V1/V4/A3/M2/s1 ));
 AND2_X1 \V4/V1/V4/A3/M2/M2/_0_  (.A1(\V4/V1/V4/A3/M2/s1 ),
    .A2(\V4/V1/V4/A3/c1 ),
    .ZN(\V4/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M2/M2/_1_  (.A(\V4/V1/V4/A3/M2/s1 ),
    .B(\V4/V1/V4/A3/c1 ),
    .Z(\V4/V1/v4 [5]));
 OR2_X1 \V4/V1/V4/A3/M2/_0_  (.A1(\V4/V1/V4/A3/M2/c1 ),
    .A2(\V4/V1/V4/A3/M2/c2 ),
    .ZN(\V4/V1/V4/A3/c2 ));
 AND2_X1 \V4/V1/V4/A3/M3/M1/_0_  (.A1(\V4/V1/V4/v4 [2]),
    .A2(\V4/V1/V4/c3 ),
    .ZN(\V4/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M3/M1/_1_  (.A(\V4/V1/V4/v4 [2]),
    .B(\V4/V1/V4/c3 ),
    .Z(\V4/V1/V4/A3/M3/s1 ));
 AND2_X1 \V4/V1/V4/A3/M3/M2/_0_  (.A1(\V4/V1/V4/A3/M3/s1 ),
    .A2(\V4/V1/V4/A3/c2 ),
    .ZN(\V4/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M3/M2/_1_  (.A(\V4/V1/V4/A3/M3/s1 ),
    .B(\V4/V1/V4/A3/c2 ),
    .Z(\V4/V1/v4 [6]));
 OR2_X1 \V4/V1/V4/A3/M3/_0_  (.A1(\V4/V1/V4/A3/M3/c1 ),
    .A2(\V4/V1/V4/A3/M3/c2 ),
    .ZN(\V4/V1/V4/A3/c3 ));
 AND2_X1 \V4/V1/V4/A3/M4/M1/_0_  (.A1(\V4/V1/V4/v4 [3]),
    .A2(ground),
    .ZN(\V4/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M4/M1/_1_  (.A(\V4/V1/V4/v4 [3]),
    .B(ground),
    .Z(\V4/V1/V4/A3/M4/s1 ));
 AND2_X1 \V4/V1/V4/A3/M4/M2/_0_  (.A1(\V4/V1/V4/A3/M4/s1 ),
    .A2(\V4/V1/V4/A3/c3 ),
    .ZN(\V4/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M4/M2/_1_  (.A(\V4/V1/V4/A3/M4/s1 ),
    .B(\V4/V1/V4/A3/c3 ),
    .Z(\V4/V1/v4 [7]));
 OR2_X1 \V4/V1/V4/A3/M4/_0_  (.A1(\V4/V1/V4/A3/M4/c1 ),
    .A2(\V4/V1/V4/A3/M4/c2 ),
    .ZN(\V4/V1/V4/overflow ));
 AND2_X1 \V4/V1/V4/V1/HA1/_0_  (.A1(\V4/V1/V4/V1/w2 ),
    .A2(\V4/V1/V4/V1/w1 ),
    .ZN(\V4/V1/V4/V1/w4 ));
 XOR2_X2 \V4/V1/V4/V1/HA1/_1_  (.A(\V4/V1/V4/V1/w2 ),
    .B(\V4/V1/V4/V1/w1 ),
    .Z(\V4/V1/v4 [1]));
 AND2_X1 \V4/V1/V4/V1/HA2/_0_  (.A1(\V4/V1/V4/V1/w4 ),
    .A2(\V4/V1/V4/V1/w3 ),
    .ZN(\V4/V1/V4/v1 [3]));
 XOR2_X2 \V4/V1/V4/V1/HA2/_1_  (.A(\V4/V1/V4/V1/w4 ),
    .B(\V4/V1/V4/V1/w3 ),
    .Z(\V4/V1/V4/v1 [2]));
 AND2_X1 \V4/V1/V4/V1/_0_  (.A1(A[20]),
    .A2(B[20]),
    .ZN(\V4/V1/v4 [0]));
 AND2_X1 \V4/V1/V4/V1/_1_  (.A1(A[20]),
    .A2(B[21]),
    .ZN(\V4/V1/V4/V1/w1 ));
 AND2_X1 \V4/V1/V4/V1/_2_  (.A1(B[20]),
    .A2(A[21]),
    .ZN(\V4/V1/V4/V1/w2 ));
 AND2_X1 \V4/V1/V4/V1/_3_  (.A1(B[21]),
    .A2(A[21]),
    .ZN(\V4/V1/V4/V1/w3 ));
 AND2_X1 \V4/V1/V4/V2/HA1/_0_  (.A1(\V4/V1/V4/V2/w2 ),
    .A2(\V4/V1/V4/V2/w1 ),
    .ZN(\V4/V1/V4/V2/w4 ));
 XOR2_X2 \V4/V1/V4/V2/HA1/_1_  (.A(\V4/V1/V4/V2/w2 ),
    .B(\V4/V1/V4/V2/w1 ),
    .Z(\V4/V1/V4/v2 [1]));
 AND2_X1 \V4/V1/V4/V2/HA2/_0_  (.A1(\V4/V1/V4/V2/w4 ),
    .A2(\V4/V1/V4/V2/w3 ),
    .ZN(\V4/V1/V4/v2 [3]));
 XOR2_X2 \V4/V1/V4/V2/HA2/_1_  (.A(\V4/V1/V4/V2/w4 ),
    .B(\V4/V1/V4/V2/w3 ),
    .Z(\V4/V1/V4/v2 [2]));
 AND2_X1 \V4/V1/V4/V2/_0_  (.A1(A[22]),
    .A2(B[20]),
    .ZN(\V4/V1/V4/v2 [0]));
 AND2_X1 \V4/V1/V4/V2/_1_  (.A1(A[22]),
    .A2(B[21]),
    .ZN(\V4/V1/V4/V2/w1 ));
 AND2_X1 \V4/V1/V4/V2/_2_  (.A1(B[20]),
    .A2(A[23]),
    .ZN(\V4/V1/V4/V2/w2 ));
 AND2_X1 \V4/V1/V4/V2/_3_  (.A1(B[21]),
    .A2(A[23]),
    .ZN(\V4/V1/V4/V2/w3 ));
 AND2_X1 \V4/V1/V4/V3/HA1/_0_  (.A1(\V4/V1/V4/V3/w2 ),
    .A2(\V4/V1/V4/V3/w1 ),
    .ZN(\V4/V1/V4/V3/w4 ));
 XOR2_X2 \V4/V1/V4/V3/HA1/_1_  (.A(\V4/V1/V4/V3/w2 ),
    .B(\V4/V1/V4/V3/w1 ),
    .Z(\V4/V1/V4/v3 [1]));
 AND2_X1 \V4/V1/V4/V3/HA2/_0_  (.A1(\V4/V1/V4/V3/w4 ),
    .A2(\V4/V1/V4/V3/w3 ),
    .ZN(\V4/V1/V4/v3 [3]));
 XOR2_X2 \V4/V1/V4/V3/HA2/_1_  (.A(\V4/V1/V4/V3/w4 ),
    .B(\V4/V1/V4/V3/w3 ),
    .Z(\V4/V1/V4/v3 [2]));
 AND2_X1 \V4/V1/V4/V3/_0_  (.A1(A[20]),
    .A2(B[22]),
    .ZN(\V4/V1/V4/v3 [0]));
 AND2_X1 \V4/V1/V4/V3/_1_  (.A1(A[20]),
    .A2(B[23]),
    .ZN(\V4/V1/V4/V3/w1 ));
 AND2_X1 \V4/V1/V4/V3/_2_  (.A1(B[22]),
    .A2(A[21]),
    .ZN(\V4/V1/V4/V3/w2 ));
 AND2_X1 \V4/V1/V4/V3/_3_  (.A1(B[23]),
    .A2(A[21]),
    .ZN(\V4/V1/V4/V3/w3 ));
 AND2_X1 \V4/V1/V4/V4/HA1/_0_  (.A1(\V4/V1/V4/V4/w2 ),
    .A2(\V4/V1/V4/V4/w1 ),
    .ZN(\V4/V1/V4/V4/w4 ));
 XOR2_X2 \V4/V1/V4/V4/HA1/_1_  (.A(\V4/V1/V4/V4/w2 ),
    .B(\V4/V1/V4/V4/w1 ),
    .Z(\V4/V1/V4/v4 [1]));
 AND2_X1 \V4/V1/V4/V4/HA2/_0_  (.A1(\V4/V1/V4/V4/w4 ),
    .A2(\V4/V1/V4/V4/w3 ),
    .ZN(\V4/V1/V4/v4 [3]));
 XOR2_X2 \V4/V1/V4/V4/HA2/_1_  (.A(\V4/V1/V4/V4/w4 ),
    .B(\V4/V1/V4/V4/w3 ),
    .Z(\V4/V1/V4/v4 [2]));
 AND2_X1 \V4/V1/V4/V4/_0_  (.A1(A[22]),
    .A2(B[22]),
    .ZN(\V4/V1/V4/v4 [0]));
 AND2_X1 \V4/V1/V4/V4/_1_  (.A1(A[22]),
    .A2(B[23]),
    .ZN(\V4/V1/V4/V4/w1 ));
 AND2_X1 \V4/V1/V4/V4/_2_  (.A1(B[22]),
    .A2(A[23]),
    .ZN(\V4/V1/V4/V4/w2 ));
 AND2_X1 \V4/V1/V4/V4/_3_  (.A1(B[23]),
    .A2(A[23]),
    .ZN(\V4/V1/V4/V4/w3 ));
 OR2_X1 \V4/V1/V4/_0_  (.A1(\V4/V1/V4/c1 ),
    .A2(\V4/V1/V4/c2 ),
    .ZN(\V4/V1/V4/c3 ));
 OR2_X1 \V4/V1/_0_  (.A1(\V4/V1/c1 ),
    .A2(\V4/V1/c2 ),
    .ZN(\V4/V1/c3 ));
 AND2_X1 \V4/V2/A1/A1/M1/M1/_0_  (.A1(\V4/V2/v2 [0]),
    .A2(\V4/V2/v3 [0]),
    .ZN(\V4/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M1/M1/_1_  (.A(\V4/V2/v2 [0]),
    .B(\V4/V2/v3 [0]),
    .Z(\V4/V2/A1/A1/M1/s1 ));
 AND2_X1 \V4/V2/A1/A1/M1/M2/_0_  (.A1(\V4/V2/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M1/M2/_1_  (.A(\V4/V2/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/s1 [0]));
 OR2_X1 \V4/V2/A1/A1/M1/_0_  (.A1(\V4/V2/A1/A1/M1/c1 ),
    .A2(\V4/V2/A1/A1/M1/c2 ),
    .ZN(\V4/V2/A1/A1/c1 ));
 AND2_X1 \V4/V2/A1/A1/M2/M1/_0_  (.A1(\V4/V2/v2 [1]),
    .A2(\V4/V2/v3 [1]),
    .ZN(\V4/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M2/M1/_1_  (.A(\V4/V2/v2 [1]),
    .B(\V4/V2/v3 [1]),
    .Z(\V4/V2/A1/A1/M2/s1 ));
 AND2_X1 \V4/V2/A1/A1/M2/M2/_0_  (.A1(\V4/V2/A1/A1/M2/s1 ),
    .A2(\V4/V2/A1/A1/c1 ),
    .ZN(\V4/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M2/M2/_1_  (.A(\V4/V2/A1/A1/M2/s1 ),
    .B(\V4/V2/A1/A1/c1 ),
    .Z(\V4/V2/s1 [1]));
 OR2_X1 \V4/V2/A1/A1/M2/_0_  (.A1(\V4/V2/A1/A1/M2/c1 ),
    .A2(\V4/V2/A1/A1/M2/c2 ),
    .ZN(\V4/V2/A1/A1/c2 ));
 AND2_X1 \V4/V2/A1/A1/M3/M1/_0_  (.A1(\V4/V2/v2 [2]),
    .A2(\V4/V2/v3 [2]),
    .ZN(\V4/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M3/M1/_1_  (.A(\V4/V2/v2 [2]),
    .B(\V4/V2/v3 [2]),
    .Z(\V4/V2/A1/A1/M3/s1 ));
 AND2_X1 \V4/V2/A1/A1/M3/M2/_0_  (.A1(\V4/V2/A1/A1/M3/s1 ),
    .A2(\V4/V2/A1/A1/c2 ),
    .ZN(\V4/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M3/M2/_1_  (.A(\V4/V2/A1/A1/M3/s1 ),
    .B(\V4/V2/A1/A1/c2 ),
    .Z(\V4/V2/s1 [2]));
 OR2_X1 \V4/V2/A1/A1/M3/_0_  (.A1(\V4/V2/A1/A1/M3/c1 ),
    .A2(\V4/V2/A1/A1/M3/c2 ),
    .ZN(\V4/V2/A1/A1/c3 ));
 AND2_X1 \V4/V2/A1/A1/M4/M1/_0_  (.A1(\V4/V2/v2 [3]),
    .A2(\V4/V2/v3 [3]),
    .ZN(\V4/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M4/M1/_1_  (.A(\V4/V2/v2 [3]),
    .B(\V4/V2/v3 [3]),
    .Z(\V4/V2/A1/A1/M4/s1 ));
 AND2_X1 \V4/V2/A1/A1/M4/M2/_0_  (.A1(\V4/V2/A1/A1/M4/s1 ),
    .A2(\V4/V2/A1/A1/c3 ),
    .ZN(\V4/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M4/M2/_1_  (.A(\V4/V2/A1/A1/M4/s1 ),
    .B(\V4/V2/A1/A1/c3 ),
    .Z(\V4/V2/s1 [3]));
 OR2_X1 \V4/V2/A1/A1/M4/_0_  (.A1(\V4/V2/A1/A1/M4/c1 ),
    .A2(\V4/V2/A1/A1/M4/c2 ),
    .ZN(\V4/V2/A1/c1 ));
 AND2_X1 \V4/V2/A1/A2/M1/M1/_0_  (.A1(\V4/V2/v2 [4]),
    .A2(\V4/V2/v3 [4]),
    .ZN(\V4/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M1/M1/_1_  (.A(\V4/V2/v2 [4]),
    .B(\V4/V2/v3 [4]),
    .Z(\V4/V2/A1/A2/M1/s1 ));
 AND2_X1 \V4/V2/A1/A2/M1/M2/_0_  (.A1(\V4/V2/A1/A2/M1/s1 ),
    .A2(\V4/V2/A1/c1 ),
    .ZN(\V4/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M1/M2/_1_  (.A(\V4/V2/A1/A2/M1/s1 ),
    .B(\V4/V2/A1/c1 ),
    .Z(\V4/V2/s1 [4]));
 OR2_X1 \V4/V2/A1/A2/M1/_0_  (.A1(\V4/V2/A1/A2/M1/c1 ),
    .A2(\V4/V2/A1/A2/M1/c2 ),
    .ZN(\V4/V2/A1/A2/c1 ));
 AND2_X1 \V4/V2/A1/A2/M2/M1/_0_  (.A1(\V4/V2/v2 [5]),
    .A2(\V4/V2/v3 [5]),
    .ZN(\V4/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M2/M1/_1_  (.A(\V4/V2/v2 [5]),
    .B(\V4/V2/v3 [5]),
    .Z(\V4/V2/A1/A2/M2/s1 ));
 AND2_X1 \V4/V2/A1/A2/M2/M2/_0_  (.A1(\V4/V2/A1/A2/M2/s1 ),
    .A2(\V4/V2/A1/A2/c1 ),
    .ZN(\V4/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M2/M2/_1_  (.A(\V4/V2/A1/A2/M2/s1 ),
    .B(\V4/V2/A1/A2/c1 ),
    .Z(\V4/V2/s1 [5]));
 OR2_X1 \V4/V2/A1/A2/M2/_0_  (.A1(\V4/V2/A1/A2/M2/c1 ),
    .A2(\V4/V2/A1/A2/M2/c2 ),
    .ZN(\V4/V2/A1/A2/c2 ));
 AND2_X1 \V4/V2/A1/A2/M3/M1/_0_  (.A1(\V4/V2/v2 [6]),
    .A2(\V4/V2/v3 [6]),
    .ZN(\V4/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M3/M1/_1_  (.A(\V4/V2/v2 [6]),
    .B(\V4/V2/v3 [6]),
    .Z(\V4/V2/A1/A2/M3/s1 ));
 AND2_X1 \V4/V2/A1/A2/M3/M2/_0_  (.A1(\V4/V2/A1/A2/M3/s1 ),
    .A2(\V4/V2/A1/A2/c2 ),
    .ZN(\V4/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M3/M2/_1_  (.A(\V4/V2/A1/A2/M3/s1 ),
    .B(\V4/V2/A1/A2/c2 ),
    .Z(\V4/V2/s1 [6]));
 OR2_X1 \V4/V2/A1/A2/M3/_0_  (.A1(\V4/V2/A1/A2/M3/c1 ),
    .A2(\V4/V2/A1/A2/M3/c2 ),
    .ZN(\V4/V2/A1/A2/c3 ));
 AND2_X1 \V4/V2/A1/A2/M4/M1/_0_  (.A1(\V4/V2/v2 [7]),
    .A2(\V4/V2/v3 [7]),
    .ZN(\V4/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M4/M1/_1_  (.A(\V4/V2/v2 [7]),
    .B(\V4/V2/v3 [7]),
    .Z(\V4/V2/A1/A2/M4/s1 ));
 AND2_X1 \V4/V2/A1/A2/M4/M2/_0_  (.A1(\V4/V2/A1/A2/M4/s1 ),
    .A2(\V4/V2/A1/A2/c3 ),
    .ZN(\V4/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M4/M2/_1_  (.A(\V4/V2/A1/A2/M4/s1 ),
    .B(\V4/V2/A1/A2/c3 ),
    .Z(\V4/V2/s1 [7]));
 OR2_X1 \V4/V2/A1/A2/M4/_0_  (.A1(\V4/V2/A1/A2/M4/c1 ),
    .A2(\V4/V2/A1/A2/M4/c2 ),
    .ZN(\V4/V2/c1 ));
 AND2_X1 \V4/V2/A2/A1/M1/M1/_0_  (.A1(\V4/V2/s1 [0]),
    .A2(\V4/V2/v1 [4]),
    .ZN(\V4/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M1/M1/_1_  (.A(\V4/V2/s1 [0]),
    .B(\V4/V2/v1 [4]),
    .Z(\V4/V2/A2/A1/M1/s1 ));
 AND2_X1 \V4/V2/A2/A1/M1/M2/_0_  (.A1(\V4/V2/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M1/M2/_1_  (.A(\V4/V2/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v2 [4]));
 OR2_X1 \V4/V2/A2/A1/M1/_0_  (.A1(\V4/V2/A2/A1/M1/c1 ),
    .A2(\V4/V2/A2/A1/M1/c2 ),
    .ZN(\V4/V2/A2/A1/c1 ));
 AND2_X1 \V4/V2/A2/A1/M2/M1/_0_  (.A1(\V4/V2/s1 [1]),
    .A2(\V4/V2/v1 [5]),
    .ZN(\V4/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M2/M1/_1_  (.A(\V4/V2/s1 [1]),
    .B(\V4/V2/v1 [5]),
    .Z(\V4/V2/A2/A1/M2/s1 ));
 AND2_X1 \V4/V2/A2/A1/M2/M2/_0_  (.A1(\V4/V2/A2/A1/M2/s1 ),
    .A2(\V4/V2/A2/A1/c1 ),
    .ZN(\V4/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M2/M2/_1_  (.A(\V4/V2/A2/A1/M2/s1 ),
    .B(\V4/V2/A2/A1/c1 ),
    .Z(\V4/v2 [5]));
 OR2_X1 \V4/V2/A2/A1/M2/_0_  (.A1(\V4/V2/A2/A1/M2/c1 ),
    .A2(\V4/V2/A2/A1/M2/c2 ),
    .ZN(\V4/V2/A2/A1/c2 ));
 AND2_X1 \V4/V2/A2/A1/M3/M1/_0_  (.A1(\V4/V2/s1 [2]),
    .A2(\V4/V2/v1 [6]),
    .ZN(\V4/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M3/M1/_1_  (.A(\V4/V2/s1 [2]),
    .B(\V4/V2/v1 [6]),
    .Z(\V4/V2/A2/A1/M3/s1 ));
 AND2_X1 \V4/V2/A2/A1/M3/M2/_0_  (.A1(\V4/V2/A2/A1/M3/s1 ),
    .A2(\V4/V2/A2/A1/c2 ),
    .ZN(\V4/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M3/M2/_1_  (.A(\V4/V2/A2/A1/M3/s1 ),
    .B(\V4/V2/A2/A1/c2 ),
    .Z(\V4/v2 [6]));
 OR2_X1 \V4/V2/A2/A1/M3/_0_  (.A1(\V4/V2/A2/A1/M3/c1 ),
    .A2(\V4/V2/A2/A1/M3/c2 ),
    .ZN(\V4/V2/A2/A1/c3 ));
 AND2_X1 \V4/V2/A2/A1/M4/M1/_0_  (.A1(\V4/V2/s1 [3]),
    .A2(\V4/V2/v1 [7]),
    .ZN(\V4/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M4/M1/_1_  (.A(\V4/V2/s1 [3]),
    .B(\V4/V2/v1 [7]),
    .Z(\V4/V2/A2/A1/M4/s1 ));
 AND2_X1 \V4/V2/A2/A1/M4/M2/_0_  (.A1(\V4/V2/A2/A1/M4/s1 ),
    .A2(\V4/V2/A2/A1/c3 ),
    .ZN(\V4/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M4/M2/_1_  (.A(\V4/V2/A2/A1/M4/s1 ),
    .B(\V4/V2/A2/A1/c3 ),
    .Z(\V4/v2 [7]));
 OR2_X1 \V4/V2/A2/A1/M4/_0_  (.A1(\V4/V2/A2/A1/M4/c1 ),
    .A2(\V4/V2/A2/A1/M4/c2 ),
    .ZN(\V4/V2/A2/c1 ));
 AND2_X1 \V4/V2/A2/A2/M1/M1/_0_  (.A1(\V4/V2/s1 [4]),
    .A2(ground),
    .ZN(\V4/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M1/M1/_1_  (.A(\V4/V2/s1 [4]),
    .B(ground),
    .Z(\V4/V2/A2/A2/M1/s1 ));
 AND2_X1 \V4/V2/A2/A2/M1/M2/_0_  (.A1(\V4/V2/A2/A2/M1/s1 ),
    .A2(\V4/V2/A2/c1 ),
    .ZN(\V4/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M1/M2/_1_  (.A(\V4/V2/A2/A2/M1/s1 ),
    .B(\V4/V2/A2/c1 ),
    .Z(\V4/V2/s2 [4]));
 OR2_X1 \V4/V2/A2/A2/M1/_0_  (.A1(\V4/V2/A2/A2/M1/c1 ),
    .A2(\V4/V2/A2/A2/M1/c2 ),
    .ZN(\V4/V2/A2/A2/c1 ));
 AND2_X1 \V4/V2/A2/A2/M2/M1/_0_  (.A1(\V4/V2/s1 [5]),
    .A2(ground),
    .ZN(\V4/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M2/M1/_1_  (.A(\V4/V2/s1 [5]),
    .B(ground),
    .Z(\V4/V2/A2/A2/M2/s1 ));
 AND2_X1 \V4/V2/A2/A2/M2/M2/_0_  (.A1(\V4/V2/A2/A2/M2/s1 ),
    .A2(\V4/V2/A2/A2/c1 ),
    .ZN(\V4/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M2/M2/_1_  (.A(\V4/V2/A2/A2/M2/s1 ),
    .B(\V4/V2/A2/A2/c1 ),
    .Z(\V4/V2/s2 [5]));
 OR2_X1 \V4/V2/A2/A2/M2/_0_  (.A1(\V4/V2/A2/A2/M2/c1 ),
    .A2(\V4/V2/A2/A2/M2/c2 ),
    .ZN(\V4/V2/A2/A2/c2 ));
 AND2_X1 \V4/V2/A2/A2/M3/M1/_0_  (.A1(\V4/V2/s1 [6]),
    .A2(ground),
    .ZN(\V4/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M3/M1/_1_  (.A(\V4/V2/s1 [6]),
    .B(ground),
    .Z(\V4/V2/A2/A2/M3/s1 ));
 AND2_X1 \V4/V2/A2/A2/M3/M2/_0_  (.A1(\V4/V2/A2/A2/M3/s1 ),
    .A2(\V4/V2/A2/A2/c2 ),
    .ZN(\V4/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M3/M2/_1_  (.A(\V4/V2/A2/A2/M3/s1 ),
    .B(\V4/V2/A2/A2/c2 ),
    .Z(\V4/V2/s2 [6]));
 OR2_X1 \V4/V2/A2/A2/M3/_0_  (.A1(\V4/V2/A2/A2/M3/c1 ),
    .A2(\V4/V2/A2/A2/M3/c2 ),
    .ZN(\V4/V2/A2/A2/c3 ));
 AND2_X1 \V4/V2/A2/A2/M4/M1/_0_  (.A1(\V4/V2/s1 [7]),
    .A2(ground),
    .ZN(\V4/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M4/M1/_1_  (.A(\V4/V2/s1 [7]),
    .B(ground),
    .Z(\V4/V2/A2/A2/M4/s1 ));
 AND2_X1 \V4/V2/A2/A2/M4/M2/_0_  (.A1(\V4/V2/A2/A2/M4/s1 ),
    .A2(\V4/V2/A2/A2/c3 ),
    .ZN(\V4/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M4/M2/_1_  (.A(\V4/V2/A2/A2/M4/s1 ),
    .B(\V4/V2/A2/A2/c3 ),
    .Z(\V4/V2/s2 [7]));
 OR2_X1 \V4/V2/A2/A2/M4/_0_  (.A1(\V4/V2/A2/A2/M4/c1 ),
    .A2(\V4/V2/A2/A2/M4/c2 ),
    .ZN(\V4/V2/c2 ));
 AND2_X1 \V4/V2/A3/A1/M1/M1/_0_  (.A1(\V4/V2/v4 [0]),
    .A2(\V4/V2/s2 [4]),
    .ZN(\V4/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M1/M1/_1_  (.A(\V4/V2/v4 [0]),
    .B(\V4/V2/s2 [4]),
    .Z(\V4/V2/A3/A1/M1/s1 ));
 AND2_X1 \V4/V2/A3/A1/M1/M2/_0_  (.A1(\V4/V2/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M1/M2/_1_  (.A(\V4/V2/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v2 [8]));
 OR2_X1 \V4/V2/A3/A1/M1/_0_  (.A1(\V4/V2/A3/A1/M1/c1 ),
    .A2(\V4/V2/A3/A1/M1/c2 ),
    .ZN(\V4/V2/A3/A1/c1 ));
 AND2_X1 \V4/V2/A3/A1/M2/M1/_0_  (.A1(\V4/V2/v4 [1]),
    .A2(\V4/V2/s2 [5]),
    .ZN(\V4/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M2/M1/_1_  (.A(\V4/V2/v4 [1]),
    .B(\V4/V2/s2 [5]),
    .Z(\V4/V2/A3/A1/M2/s1 ));
 AND2_X1 \V4/V2/A3/A1/M2/M2/_0_  (.A1(\V4/V2/A3/A1/M2/s1 ),
    .A2(\V4/V2/A3/A1/c1 ),
    .ZN(\V4/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M2/M2/_1_  (.A(\V4/V2/A3/A1/M2/s1 ),
    .B(\V4/V2/A3/A1/c1 ),
    .Z(\V4/v2 [9]));
 OR2_X1 \V4/V2/A3/A1/M2/_0_  (.A1(\V4/V2/A3/A1/M2/c1 ),
    .A2(\V4/V2/A3/A1/M2/c2 ),
    .ZN(\V4/V2/A3/A1/c2 ));
 AND2_X1 \V4/V2/A3/A1/M3/M1/_0_  (.A1(\V4/V2/v4 [2]),
    .A2(\V4/V2/s2 [6]),
    .ZN(\V4/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M3/M1/_1_  (.A(\V4/V2/v4 [2]),
    .B(\V4/V2/s2 [6]),
    .Z(\V4/V2/A3/A1/M3/s1 ));
 AND2_X1 \V4/V2/A3/A1/M3/M2/_0_  (.A1(\V4/V2/A3/A1/M3/s1 ),
    .A2(\V4/V2/A3/A1/c2 ),
    .ZN(\V4/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M3/M2/_1_  (.A(\V4/V2/A3/A1/M3/s1 ),
    .B(\V4/V2/A3/A1/c2 ),
    .Z(\V4/v2 [10]));
 OR2_X1 \V4/V2/A3/A1/M3/_0_  (.A1(\V4/V2/A3/A1/M3/c1 ),
    .A2(\V4/V2/A3/A1/M3/c2 ),
    .ZN(\V4/V2/A3/A1/c3 ));
 AND2_X1 \V4/V2/A3/A1/M4/M1/_0_  (.A1(\V4/V2/v4 [3]),
    .A2(\V4/V2/s2 [7]),
    .ZN(\V4/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M4/M1/_1_  (.A(\V4/V2/v4 [3]),
    .B(\V4/V2/s2 [7]),
    .Z(\V4/V2/A3/A1/M4/s1 ));
 AND2_X1 \V4/V2/A3/A1/M4/M2/_0_  (.A1(\V4/V2/A3/A1/M4/s1 ),
    .A2(\V4/V2/A3/A1/c3 ),
    .ZN(\V4/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M4/M2/_1_  (.A(\V4/V2/A3/A1/M4/s1 ),
    .B(\V4/V2/A3/A1/c3 ),
    .Z(\V4/v2 [11]));
 OR2_X1 \V4/V2/A3/A1/M4/_0_  (.A1(\V4/V2/A3/A1/M4/c1 ),
    .A2(\V4/V2/A3/A1/M4/c2 ),
    .ZN(\V4/V2/A3/c1 ));
 AND2_X1 \V4/V2/A3/A2/M1/M1/_0_  (.A1(\V4/V2/v4 [4]),
    .A2(\V4/V2/c3 ),
    .ZN(\V4/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M1/M1/_1_  (.A(\V4/V2/v4 [4]),
    .B(\V4/V2/c3 ),
    .Z(\V4/V2/A3/A2/M1/s1 ));
 AND2_X1 \V4/V2/A3/A2/M1/M2/_0_  (.A1(\V4/V2/A3/A2/M1/s1 ),
    .A2(\V4/V2/A3/c1 ),
    .ZN(\V4/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M1/M2/_1_  (.A(\V4/V2/A3/A2/M1/s1 ),
    .B(\V4/V2/A3/c1 ),
    .Z(\V4/v2 [12]));
 OR2_X1 \V4/V2/A3/A2/M1/_0_  (.A1(\V4/V2/A3/A2/M1/c1 ),
    .A2(\V4/V2/A3/A2/M1/c2 ),
    .ZN(\V4/V2/A3/A2/c1 ));
 AND2_X1 \V4/V2/A3/A2/M2/M1/_0_  (.A1(\V4/V2/v4 [5]),
    .A2(ground),
    .ZN(\V4/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M2/M1/_1_  (.A(\V4/V2/v4 [5]),
    .B(ground),
    .Z(\V4/V2/A3/A2/M2/s1 ));
 AND2_X1 \V4/V2/A3/A2/M2/M2/_0_  (.A1(\V4/V2/A3/A2/M2/s1 ),
    .A2(\V4/V2/A3/A2/c1 ),
    .ZN(\V4/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M2/M2/_1_  (.A(\V4/V2/A3/A2/M2/s1 ),
    .B(\V4/V2/A3/A2/c1 ),
    .Z(\V4/v2 [13]));
 OR2_X1 \V4/V2/A3/A2/M2/_0_  (.A1(\V4/V2/A3/A2/M2/c1 ),
    .A2(\V4/V2/A3/A2/M2/c2 ),
    .ZN(\V4/V2/A3/A2/c2 ));
 AND2_X1 \V4/V2/A3/A2/M3/M1/_0_  (.A1(\V4/V2/v4 [6]),
    .A2(ground),
    .ZN(\V4/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M3/M1/_1_  (.A(\V4/V2/v4 [6]),
    .B(ground),
    .Z(\V4/V2/A3/A2/M3/s1 ));
 AND2_X1 \V4/V2/A3/A2/M3/M2/_0_  (.A1(\V4/V2/A3/A2/M3/s1 ),
    .A2(\V4/V2/A3/A2/c2 ),
    .ZN(\V4/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M3/M2/_1_  (.A(\V4/V2/A3/A2/M3/s1 ),
    .B(\V4/V2/A3/A2/c2 ),
    .Z(\V4/v2 [14]));
 OR2_X1 \V4/V2/A3/A2/M3/_0_  (.A1(\V4/V2/A3/A2/M3/c1 ),
    .A2(\V4/V2/A3/A2/M3/c2 ),
    .ZN(\V4/V2/A3/A2/c3 ));
 AND2_X1 \V4/V2/A3/A2/M4/M1/_0_  (.A1(\V4/V2/v4 [7]),
    .A2(ground),
    .ZN(\V4/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M4/M1/_1_  (.A(\V4/V2/v4 [7]),
    .B(ground),
    .Z(\V4/V2/A3/A2/M4/s1 ));
 AND2_X1 \V4/V2/A3/A2/M4/M2/_0_  (.A1(\V4/V2/A3/A2/M4/s1 ),
    .A2(\V4/V2/A3/A2/c3 ),
    .ZN(\V4/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M4/M2/_1_  (.A(\V4/V2/A3/A2/M4/s1 ),
    .B(\V4/V2/A3/A2/c3 ),
    .Z(\V4/v2 [15]));
 OR2_X1 \V4/V2/A3/A2/M4/_0_  (.A1(\V4/V2/A3/A2/M4/c1 ),
    .A2(\V4/V2/A3/A2/M4/c2 ),
    .ZN(\V4/V2/overflow ));
 AND2_X1 \V4/V2/V1/A1/M1/M1/_0_  (.A1(\V4/V2/V1/v2 [0]),
    .A2(\V4/V2/V1/v3 [0]),
    .ZN(\V4/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M1/M1/_1_  (.A(\V4/V2/V1/v2 [0]),
    .B(\V4/V2/V1/v3 [0]),
    .Z(\V4/V2/V1/A1/M1/s1 ));
 AND2_X1 \V4/V2/V1/A1/M1/M2/_0_  (.A1(\V4/V2/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M1/M2/_1_  (.A(\V4/V2/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/V1/s1 [0]));
 OR2_X1 \V4/V2/V1/A1/M1/_0_  (.A1(\V4/V2/V1/A1/M1/c1 ),
    .A2(\V4/V2/V1/A1/M1/c2 ),
    .ZN(\V4/V2/V1/A1/c1 ));
 AND2_X1 \V4/V2/V1/A1/M2/M1/_0_  (.A1(\V4/V2/V1/v2 [1]),
    .A2(\V4/V2/V1/v3 [1]),
    .ZN(\V4/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M2/M1/_1_  (.A(\V4/V2/V1/v2 [1]),
    .B(\V4/V2/V1/v3 [1]),
    .Z(\V4/V2/V1/A1/M2/s1 ));
 AND2_X1 \V4/V2/V1/A1/M2/M2/_0_  (.A1(\V4/V2/V1/A1/M2/s1 ),
    .A2(\V4/V2/V1/A1/c1 ),
    .ZN(\V4/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M2/M2/_1_  (.A(\V4/V2/V1/A1/M2/s1 ),
    .B(\V4/V2/V1/A1/c1 ),
    .Z(\V4/V2/V1/s1 [1]));
 OR2_X1 \V4/V2/V1/A1/M2/_0_  (.A1(\V4/V2/V1/A1/M2/c1 ),
    .A2(\V4/V2/V1/A1/M2/c2 ),
    .ZN(\V4/V2/V1/A1/c2 ));
 AND2_X1 \V4/V2/V1/A1/M3/M1/_0_  (.A1(\V4/V2/V1/v2 [2]),
    .A2(\V4/V2/V1/v3 [2]),
    .ZN(\V4/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M3/M1/_1_  (.A(\V4/V2/V1/v2 [2]),
    .B(\V4/V2/V1/v3 [2]),
    .Z(\V4/V2/V1/A1/M3/s1 ));
 AND2_X1 \V4/V2/V1/A1/M3/M2/_0_  (.A1(\V4/V2/V1/A1/M3/s1 ),
    .A2(\V4/V2/V1/A1/c2 ),
    .ZN(\V4/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M3/M2/_1_  (.A(\V4/V2/V1/A1/M3/s1 ),
    .B(\V4/V2/V1/A1/c2 ),
    .Z(\V4/V2/V1/s1 [2]));
 OR2_X1 \V4/V2/V1/A1/M3/_0_  (.A1(\V4/V2/V1/A1/M3/c1 ),
    .A2(\V4/V2/V1/A1/M3/c2 ),
    .ZN(\V4/V2/V1/A1/c3 ));
 AND2_X1 \V4/V2/V1/A1/M4/M1/_0_  (.A1(\V4/V2/V1/v2 [3]),
    .A2(\V4/V2/V1/v3 [3]),
    .ZN(\V4/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M4/M1/_1_  (.A(\V4/V2/V1/v2 [3]),
    .B(\V4/V2/V1/v3 [3]),
    .Z(\V4/V2/V1/A1/M4/s1 ));
 AND2_X1 \V4/V2/V1/A1/M4/M2/_0_  (.A1(\V4/V2/V1/A1/M4/s1 ),
    .A2(\V4/V2/V1/A1/c3 ),
    .ZN(\V4/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M4/M2/_1_  (.A(\V4/V2/V1/A1/M4/s1 ),
    .B(\V4/V2/V1/A1/c3 ),
    .Z(\V4/V2/V1/s1 [3]));
 OR2_X1 \V4/V2/V1/A1/M4/_0_  (.A1(\V4/V2/V1/A1/M4/c1 ),
    .A2(\V4/V2/V1/A1/M4/c2 ),
    .ZN(\V4/V2/V1/c1 ));
 AND2_X1 \V4/V2/V1/A2/M1/M1/_0_  (.A1(\V4/V2/V1/s1 [0]),
    .A2(\V4/V2/V1/v1 [2]),
    .ZN(\V4/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M1/M1/_1_  (.A(\V4/V2/V1/s1 [0]),
    .B(\V4/V2/V1/v1 [2]),
    .Z(\V4/V2/V1/A2/M1/s1 ));
 AND2_X1 \V4/V2/V1/A2/M1/M2/_0_  (.A1(\V4/V2/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M1/M2/_1_  (.A(\V4/V2/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/v2 [2]));
 OR2_X1 \V4/V2/V1/A2/M1/_0_  (.A1(\V4/V2/V1/A2/M1/c1 ),
    .A2(\V4/V2/V1/A2/M1/c2 ),
    .ZN(\V4/V2/V1/A2/c1 ));
 AND2_X1 \V4/V2/V1/A2/M2/M1/_0_  (.A1(\V4/V2/V1/s1 [1]),
    .A2(\V4/V2/V1/v1 [3]),
    .ZN(\V4/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M2/M1/_1_  (.A(\V4/V2/V1/s1 [1]),
    .B(\V4/V2/V1/v1 [3]),
    .Z(\V4/V2/V1/A2/M2/s1 ));
 AND2_X1 \V4/V2/V1/A2/M2/M2/_0_  (.A1(\V4/V2/V1/A2/M2/s1 ),
    .A2(\V4/V2/V1/A2/c1 ),
    .ZN(\V4/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M2/M2/_1_  (.A(\V4/V2/V1/A2/M2/s1 ),
    .B(\V4/V2/V1/A2/c1 ),
    .Z(\V4/v2 [3]));
 OR2_X1 \V4/V2/V1/A2/M2/_0_  (.A1(\V4/V2/V1/A2/M2/c1 ),
    .A2(\V4/V2/V1/A2/M2/c2 ),
    .ZN(\V4/V2/V1/A2/c2 ));
 AND2_X1 \V4/V2/V1/A2/M3/M1/_0_  (.A1(\V4/V2/V1/s1 [2]),
    .A2(ground),
    .ZN(\V4/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M3/M1/_1_  (.A(\V4/V2/V1/s1 [2]),
    .B(ground),
    .Z(\V4/V2/V1/A2/M3/s1 ));
 AND2_X1 \V4/V2/V1/A2/M3/M2/_0_  (.A1(\V4/V2/V1/A2/M3/s1 ),
    .A2(\V4/V2/V1/A2/c2 ),
    .ZN(\V4/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M3/M2/_1_  (.A(\V4/V2/V1/A2/M3/s1 ),
    .B(\V4/V2/V1/A2/c2 ),
    .Z(\V4/V2/V1/s2 [2]));
 OR2_X1 \V4/V2/V1/A2/M3/_0_  (.A1(\V4/V2/V1/A2/M3/c1 ),
    .A2(\V4/V2/V1/A2/M3/c2 ),
    .ZN(\V4/V2/V1/A2/c3 ));
 AND2_X1 \V4/V2/V1/A2/M4/M1/_0_  (.A1(\V4/V2/V1/s1 [3]),
    .A2(ground),
    .ZN(\V4/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M4/M1/_1_  (.A(\V4/V2/V1/s1 [3]),
    .B(ground),
    .Z(\V4/V2/V1/A2/M4/s1 ));
 AND2_X1 \V4/V2/V1/A2/M4/M2/_0_  (.A1(\V4/V2/V1/A2/M4/s1 ),
    .A2(\V4/V2/V1/A2/c3 ),
    .ZN(\V4/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M4/M2/_1_  (.A(\V4/V2/V1/A2/M4/s1 ),
    .B(\V4/V2/V1/A2/c3 ),
    .Z(\V4/V2/V1/s2 [3]));
 OR2_X1 \V4/V2/V1/A2/M4/_0_  (.A1(\V4/V2/V1/A2/M4/c1 ),
    .A2(\V4/V2/V1/A2/M4/c2 ),
    .ZN(\V4/V2/V1/c2 ));
 AND2_X1 \V4/V2/V1/A3/M1/M1/_0_  (.A1(\V4/V2/V1/v4 [0]),
    .A2(\V4/V2/V1/s2 [2]),
    .ZN(\V4/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M1/M1/_1_  (.A(\V4/V2/V1/v4 [0]),
    .B(\V4/V2/V1/s2 [2]),
    .Z(\V4/V2/V1/A3/M1/s1 ));
 AND2_X1 \V4/V2/V1/A3/M1/M2/_0_  (.A1(\V4/V2/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M1/M2/_1_  (.A(\V4/V2/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v1 [4]));
 OR2_X1 \V4/V2/V1/A3/M1/_0_  (.A1(\V4/V2/V1/A3/M1/c1 ),
    .A2(\V4/V2/V1/A3/M1/c2 ),
    .ZN(\V4/V2/V1/A3/c1 ));
 AND2_X1 \V4/V2/V1/A3/M2/M1/_0_  (.A1(\V4/V2/V1/v4 [1]),
    .A2(\V4/V2/V1/s2 [3]),
    .ZN(\V4/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M2/M1/_1_  (.A(\V4/V2/V1/v4 [1]),
    .B(\V4/V2/V1/s2 [3]),
    .Z(\V4/V2/V1/A3/M2/s1 ));
 AND2_X1 \V4/V2/V1/A3/M2/M2/_0_  (.A1(\V4/V2/V1/A3/M2/s1 ),
    .A2(\V4/V2/V1/A3/c1 ),
    .ZN(\V4/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M2/M2/_1_  (.A(\V4/V2/V1/A3/M2/s1 ),
    .B(\V4/V2/V1/A3/c1 ),
    .Z(\V4/V2/v1 [5]));
 OR2_X1 \V4/V2/V1/A3/M2/_0_  (.A1(\V4/V2/V1/A3/M2/c1 ),
    .A2(\V4/V2/V1/A3/M2/c2 ),
    .ZN(\V4/V2/V1/A3/c2 ));
 AND2_X1 \V4/V2/V1/A3/M3/M1/_0_  (.A1(\V4/V2/V1/v4 [2]),
    .A2(\V4/V2/V1/c3 ),
    .ZN(\V4/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M3/M1/_1_  (.A(\V4/V2/V1/v4 [2]),
    .B(\V4/V2/V1/c3 ),
    .Z(\V4/V2/V1/A3/M3/s1 ));
 AND2_X1 \V4/V2/V1/A3/M3/M2/_0_  (.A1(\V4/V2/V1/A3/M3/s1 ),
    .A2(\V4/V2/V1/A3/c2 ),
    .ZN(\V4/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M3/M2/_1_  (.A(\V4/V2/V1/A3/M3/s1 ),
    .B(\V4/V2/V1/A3/c2 ),
    .Z(\V4/V2/v1 [6]));
 OR2_X1 \V4/V2/V1/A3/M3/_0_  (.A1(\V4/V2/V1/A3/M3/c1 ),
    .A2(\V4/V2/V1/A3/M3/c2 ),
    .ZN(\V4/V2/V1/A3/c3 ));
 AND2_X1 \V4/V2/V1/A3/M4/M1/_0_  (.A1(\V4/V2/V1/v4 [3]),
    .A2(ground),
    .ZN(\V4/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M4/M1/_1_  (.A(\V4/V2/V1/v4 [3]),
    .B(ground),
    .Z(\V4/V2/V1/A3/M4/s1 ));
 AND2_X1 \V4/V2/V1/A3/M4/M2/_0_  (.A1(\V4/V2/V1/A3/M4/s1 ),
    .A2(\V4/V2/V1/A3/c3 ),
    .ZN(\V4/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M4/M2/_1_  (.A(\V4/V2/V1/A3/M4/s1 ),
    .B(\V4/V2/V1/A3/c3 ),
    .Z(\V4/V2/v1 [7]));
 OR2_X1 \V4/V2/V1/A3/M4/_0_  (.A1(\V4/V2/V1/A3/M4/c1 ),
    .A2(\V4/V2/V1/A3/M4/c2 ),
    .ZN(\V4/V2/V1/overflow ));
 AND2_X1 \V4/V2/V1/V1/HA1/_0_  (.A1(\V4/V2/V1/V1/w2 ),
    .A2(\V4/V2/V1/V1/w1 ),
    .ZN(\V4/V2/V1/V1/w4 ));
 XOR2_X2 \V4/V2/V1/V1/HA1/_1_  (.A(\V4/V2/V1/V1/w2 ),
    .B(\V4/V2/V1/V1/w1 ),
    .Z(\V4/v2 [1]));
 AND2_X1 \V4/V2/V1/V1/HA2/_0_  (.A1(\V4/V2/V1/V1/w4 ),
    .A2(\V4/V2/V1/V1/w3 ),
    .ZN(\V4/V2/V1/v1 [3]));
 XOR2_X2 \V4/V2/V1/V1/HA2/_1_  (.A(\V4/V2/V1/V1/w4 ),
    .B(\V4/V2/V1/V1/w3 ),
    .Z(\V4/V2/V1/v1 [2]));
 AND2_X1 \V4/V2/V1/V1/_0_  (.A1(A[24]),
    .A2(B[16]),
    .ZN(\V4/v2 [0]));
 AND2_X1 \V4/V2/V1/V1/_1_  (.A1(A[24]),
    .A2(B[17]),
    .ZN(\V4/V2/V1/V1/w1 ));
 AND2_X1 \V4/V2/V1/V1/_2_  (.A1(B[16]),
    .A2(A[25]),
    .ZN(\V4/V2/V1/V1/w2 ));
 AND2_X1 \V4/V2/V1/V1/_3_  (.A1(B[17]),
    .A2(A[25]),
    .ZN(\V4/V2/V1/V1/w3 ));
 AND2_X1 \V4/V2/V1/V2/HA1/_0_  (.A1(\V4/V2/V1/V2/w2 ),
    .A2(\V4/V2/V1/V2/w1 ),
    .ZN(\V4/V2/V1/V2/w4 ));
 XOR2_X2 \V4/V2/V1/V2/HA1/_1_  (.A(\V4/V2/V1/V2/w2 ),
    .B(\V4/V2/V1/V2/w1 ),
    .Z(\V4/V2/V1/v2 [1]));
 AND2_X1 \V4/V2/V1/V2/HA2/_0_  (.A1(\V4/V2/V1/V2/w4 ),
    .A2(\V4/V2/V1/V2/w3 ),
    .ZN(\V4/V2/V1/v2 [3]));
 XOR2_X2 \V4/V2/V1/V2/HA2/_1_  (.A(\V4/V2/V1/V2/w4 ),
    .B(\V4/V2/V1/V2/w3 ),
    .Z(\V4/V2/V1/v2 [2]));
 AND2_X1 \V4/V2/V1/V2/_0_  (.A1(A[26]),
    .A2(B[16]),
    .ZN(\V4/V2/V1/v2 [0]));
 AND2_X1 \V4/V2/V1/V2/_1_  (.A1(A[26]),
    .A2(B[17]),
    .ZN(\V4/V2/V1/V2/w1 ));
 AND2_X1 \V4/V2/V1/V2/_2_  (.A1(B[16]),
    .A2(A[27]),
    .ZN(\V4/V2/V1/V2/w2 ));
 AND2_X1 \V4/V2/V1/V2/_3_  (.A1(B[17]),
    .A2(A[27]),
    .ZN(\V4/V2/V1/V2/w3 ));
 AND2_X1 \V4/V2/V1/V3/HA1/_0_  (.A1(\V4/V2/V1/V3/w2 ),
    .A2(\V4/V2/V1/V3/w1 ),
    .ZN(\V4/V2/V1/V3/w4 ));
 XOR2_X2 \V4/V2/V1/V3/HA1/_1_  (.A(\V4/V2/V1/V3/w2 ),
    .B(\V4/V2/V1/V3/w1 ),
    .Z(\V4/V2/V1/v3 [1]));
 AND2_X1 \V4/V2/V1/V3/HA2/_0_  (.A1(\V4/V2/V1/V3/w4 ),
    .A2(\V4/V2/V1/V3/w3 ),
    .ZN(\V4/V2/V1/v3 [3]));
 XOR2_X2 \V4/V2/V1/V3/HA2/_1_  (.A(\V4/V2/V1/V3/w4 ),
    .B(\V4/V2/V1/V3/w3 ),
    .Z(\V4/V2/V1/v3 [2]));
 AND2_X1 \V4/V2/V1/V3/_0_  (.A1(A[24]),
    .A2(B[18]),
    .ZN(\V4/V2/V1/v3 [0]));
 AND2_X1 \V4/V2/V1/V3/_1_  (.A1(A[24]),
    .A2(B[19]),
    .ZN(\V4/V2/V1/V3/w1 ));
 AND2_X1 \V4/V2/V1/V3/_2_  (.A1(B[18]),
    .A2(A[25]),
    .ZN(\V4/V2/V1/V3/w2 ));
 AND2_X1 \V4/V2/V1/V3/_3_  (.A1(B[19]),
    .A2(A[25]),
    .ZN(\V4/V2/V1/V3/w3 ));
 AND2_X1 \V4/V2/V1/V4/HA1/_0_  (.A1(\V4/V2/V1/V4/w2 ),
    .A2(\V4/V2/V1/V4/w1 ),
    .ZN(\V4/V2/V1/V4/w4 ));
 XOR2_X2 \V4/V2/V1/V4/HA1/_1_  (.A(\V4/V2/V1/V4/w2 ),
    .B(\V4/V2/V1/V4/w1 ),
    .Z(\V4/V2/V1/v4 [1]));
 AND2_X1 \V4/V2/V1/V4/HA2/_0_  (.A1(\V4/V2/V1/V4/w4 ),
    .A2(\V4/V2/V1/V4/w3 ),
    .ZN(\V4/V2/V1/v4 [3]));
 XOR2_X2 \V4/V2/V1/V4/HA2/_1_  (.A(\V4/V2/V1/V4/w4 ),
    .B(\V4/V2/V1/V4/w3 ),
    .Z(\V4/V2/V1/v4 [2]));
 AND2_X1 \V4/V2/V1/V4/_0_  (.A1(A[26]),
    .A2(B[18]),
    .ZN(\V4/V2/V1/v4 [0]));
 AND2_X1 \V4/V2/V1/V4/_1_  (.A1(A[26]),
    .A2(B[19]),
    .ZN(\V4/V2/V1/V4/w1 ));
 AND2_X1 \V4/V2/V1/V4/_2_  (.A1(B[18]),
    .A2(A[27]),
    .ZN(\V4/V2/V1/V4/w2 ));
 AND2_X1 \V4/V2/V1/V4/_3_  (.A1(B[19]),
    .A2(A[27]),
    .ZN(\V4/V2/V1/V4/w3 ));
 OR2_X1 \V4/V2/V1/_0_  (.A1(\V4/V2/V1/c1 ),
    .A2(\V4/V2/V1/c2 ),
    .ZN(\V4/V2/V1/c3 ));
 AND2_X1 \V4/V2/V2/A1/M1/M1/_0_  (.A1(\V4/V2/V2/v2 [0]),
    .A2(\V4/V2/V2/v3 [0]),
    .ZN(\V4/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M1/M1/_1_  (.A(\V4/V2/V2/v2 [0]),
    .B(\V4/V2/V2/v3 [0]),
    .Z(\V4/V2/V2/A1/M1/s1 ));
 AND2_X1 \V4/V2/V2/A1/M1/M2/_0_  (.A1(\V4/V2/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M1/M2/_1_  (.A(\V4/V2/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/V2/s1 [0]));
 OR2_X1 \V4/V2/V2/A1/M1/_0_  (.A1(\V4/V2/V2/A1/M1/c1 ),
    .A2(\V4/V2/V2/A1/M1/c2 ),
    .ZN(\V4/V2/V2/A1/c1 ));
 AND2_X1 \V4/V2/V2/A1/M2/M1/_0_  (.A1(\V4/V2/V2/v2 [1]),
    .A2(\V4/V2/V2/v3 [1]),
    .ZN(\V4/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M2/M1/_1_  (.A(\V4/V2/V2/v2 [1]),
    .B(\V4/V2/V2/v3 [1]),
    .Z(\V4/V2/V2/A1/M2/s1 ));
 AND2_X1 \V4/V2/V2/A1/M2/M2/_0_  (.A1(\V4/V2/V2/A1/M2/s1 ),
    .A2(\V4/V2/V2/A1/c1 ),
    .ZN(\V4/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M2/M2/_1_  (.A(\V4/V2/V2/A1/M2/s1 ),
    .B(\V4/V2/V2/A1/c1 ),
    .Z(\V4/V2/V2/s1 [1]));
 OR2_X1 \V4/V2/V2/A1/M2/_0_  (.A1(\V4/V2/V2/A1/M2/c1 ),
    .A2(\V4/V2/V2/A1/M2/c2 ),
    .ZN(\V4/V2/V2/A1/c2 ));
 AND2_X1 \V4/V2/V2/A1/M3/M1/_0_  (.A1(\V4/V2/V2/v2 [2]),
    .A2(\V4/V2/V2/v3 [2]),
    .ZN(\V4/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M3/M1/_1_  (.A(\V4/V2/V2/v2 [2]),
    .B(\V4/V2/V2/v3 [2]),
    .Z(\V4/V2/V2/A1/M3/s1 ));
 AND2_X1 \V4/V2/V2/A1/M3/M2/_0_  (.A1(\V4/V2/V2/A1/M3/s1 ),
    .A2(\V4/V2/V2/A1/c2 ),
    .ZN(\V4/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M3/M2/_1_  (.A(\V4/V2/V2/A1/M3/s1 ),
    .B(\V4/V2/V2/A1/c2 ),
    .Z(\V4/V2/V2/s1 [2]));
 OR2_X1 \V4/V2/V2/A1/M3/_0_  (.A1(\V4/V2/V2/A1/M3/c1 ),
    .A2(\V4/V2/V2/A1/M3/c2 ),
    .ZN(\V4/V2/V2/A1/c3 ));
 AND2_X1 \V4/V2/V2/A1/M4/M1/_0_  (.A1(\V4/V2/V2/v2 [3]),
    .A2(\V4/V2/V2/v3 [3]),
    .ZN(\V4/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M4/M1/_1_  (.A(\V4/V2/V2/v2 [3]),
    .B(\V4/V2/V2/v3 [3]),
    .Z(\V4/V2/V2/A1/M4/s1 ));
 AND2_X1 \V4/V2/V2/A1/M4/M2/_0_  (.A1(\V4/V2/V2/A1/M4/s1 ),
    .A2(\V4/V2/V2/A1/c3 ),
    .ZN(\V4/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M4/M2/_1_  (.A(\V4/V2/V2/A1/M4/s1 ),
    .B(\V4/V2/V2/A1/c3 ),
    .Z(\V4/V2/V2/s1 [3]));
 OR2_X1 \V4/V2/V2/A1/M4/_0_  (.A1(\V4/V2/V2/A1/M4/c1 ),
    .A2(\V4/V2/V2/A1/M4/c2 ),
    .ZN(\V4/V2/V2/c1 ));
 AND2_X1 \V4/V2/V2/A2/M1/M1/_0_  (.A1(\V4/V2/V2/s1 [0]),
    .A2(\V4/V2/V2/v1 [2]),
    .ZN(\V4/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M1/M1/_1_  (.A(\V4/V2/V2/s1 [0]),
    .B(\V4/V2/V2/v1 [2]),
    .Z(\V4/V2/V2/A2/M1/s1 ));
 AND2_X1 \V4/V2/V2/A2/M1/M2/_0_  (.A1(\V4/V2/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M1/M2/_1_  (.A(\V4/V2/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v2 [2]));
 OR2_X1 \V4/V2/V2/A2/M1/_0_  (.A1(\V4/V2/V2/A2/M1/c1 ),
    .A2(\V4/V2/V2/A2/M1/c2 ),
    .ZN(\V4/V2/V2/A2/c1 ));
 AND2_X1 \V4/V2/V2/A2/M2/M1/_0_  (.A1(\V4/V2/V2/s1 [1]),
    .A2(\V4/V2/V2/v1 [3]),
    .ZN(\V4/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M2/M1/_1_  (.A(\V4/V2/V2/s1 [1]),
    .B(\V4/V2/V2/v1 [3]),
    .Z(\V4/V2/V2/A2/M2/s1 ));
 AND2_X1 \V4/V2/V2/A2/M2/M2/_0_  (.A1(\V4/V2/V2/A2/M2/s1 ),
    .A2(\V4/V2/V2/A2/c1 ),
    .ZN(\V4/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M2/M2/_1_  (.A(\V4/V2/V2/A2/M2/s1 ),
    .B(\V4/V2/V2/A2/c1 ),
    .Z(\V4/V2/v2 [3]));
 OR2_X1 \V4/V2/V2/A2/M2/_0_  (.A1(\V4/V2/V2/A2/M2/c1 ),
    .A2(\V4/V2/V2/A2/M2/c2 ),
    .ZN(\V4/V2/V2/A2/c2 ));
 AND2_X1 \V4/V2/V2/A2/M3/M1/_0_  (.A1(\V4/V2/V2/s1 [2]),
    .A2(ground),
    .ZN(\V4/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M3/M1/_1_  (.A(\V4/V2/V2/s1 [2]),
    .B(ground),
    .Z(\V4/V2/V2/A2/M3/s1 ));
 AND2_X1 \V4/V2/V2/A2/M3/M2/_0_  (.A1(\V4/V2/V2/A2/M3/s1 ),
    .A2(\V4/V2/V2/A2/c2 ),
    .ZN(\V4/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M3/M2/_1_  (.A(\V4/V2/V2/A2/M3/s1 ),
    .B(\V4/V2/V2/A2/c2 ),
    .Z(\V4/V2/V2/s2 [2]));
 OR2_X1 \V4/V2/V2/A2/M3/_0_  (.A1(\V4/V2/V2/A2/M3/c1 ),
    .A2(\V4/V2/V2/A2/M3/c2 ),
    .ZN(\V4/V2/V2/A2/c3 ));
 AND2_X1 \V4/V2/V2/A2/M4/M1/_0_  (.A1(\V4/V2/V2/s1 [3]),
    .A2(ground),
    .ZN(\V4/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M4/M1/_1_  (.A(\V4/V2/V2/s1 [3]),
    .B(ground),
    .Z(\V4/V2/V2/A2/M4/s1 ));
 AND2_X1 \V4/V2/V2/A2/M4/M2/_0_  (.A1(\V4/V2/V2/A2/M4/s1 ),
    .A2(\V4/V2/V2/A2/c3 ),
    .ZN(\V4/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M4/M2/_1_  (.A(\V4/V2/V2/A2/M4/s1 ),
    .B(\V4/V2/V2/A2/c3 ),
    .Z(\V4/V2/V2/s2 [3]));
 OR2_X1 \V4/V2/V2/A2/M4/_0_  (.A1(\V4/V2/V2/A2/M4/c1 ),
    .A2(\V4/V2/V2/A2/M4/c2 ),
    .ZN(\V4/V2/V2/c2 ));
 AND2_X1 \V4/V2/V2/A3/M1/M1/_0_  (.A1(\V4/V2/V2/v4 [0]),
    .A2(\V4/V2/V2/s2 [2]),
    .ZN(\V4/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M1/M1/_1_  (.A(\V4/V2/V2/v4 [0]),
    .B(\V4/V2/V2/s2 [2]),
    .Z(\V4/V2/V2/A3/M1/s1 ));
 AND2_X1 \V4/V2/V2/A3/M1/M2/_0_  (.A1(\V4/V2/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M1/M2/_1_  (.A(\V4/V2/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v2 [4]));
 OR2_X1 \V4/V2/V2/A3/M1/_0_  (.A1(\V4/V2/V2/A3/M1/c1 ),
    .A2(\V4/V2/V2/A3/M1/c2 ),
    .ZN(\V4/V2/V2/A3/c1 ));
 AND2_X1 \V4/V2/V2/A3/M2/M1/_0_  (.A1(\V4/V2/V2/v4 [1]),
    .A2(\V4/V2/V2/s2 [3]),
    .ZN(\V4/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M2/M1/_1_  (.A(\V4/V2/V2/v4 [1]),
    .B(\V4/V2/V2/s2 [3]),
    .Z(\V4/V2/V2/A3/M2/s1 ));
 AND2_X1 \V4/V2/V2/A3/M2/M2/_0_  (.A1(\V4/V2/V2/A3/M2/s1 ),
    .A2(\V4/V2/V2/A3/c1 ),
    .ZN(\V4/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M2/M2/_1_  (.A(\V4/V2/V2/A3/M2/s1 ),
    .B(\V4/V2/V2/A3/c1 ),
    .Z(\V4/V2/v2 [5]));
 OR2_X1 \V4/V2/V2/A3/M2/_0_  (.A1(\V4/V2/V2/A3/M2/c1 ),
    .A2(\V4/V2/V2/A3/M2/c2 ),
    .ZN(\V4/V2/V2/A3/c2 ));
 AND2_X1 \V4/V2/V2/A3/M3/M1/_0_  (.A1(\V4/V2/V2/v4 [2]),
    .A2(\V4/V2/V2/c3 ),
    .ZN(\V4/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M3/M1/_1_  (.A(\V4/V2/V2/v4 [2]),
    .B(\V4/V2/V2/c3 ),
    .Z(\V4/V2/V2/A3/M3/s1 ));
 AND2_X1 \V4/V2/V2/A3/M3/M2/_0_  (.A1(\V4/V2/V2/A3/M3/s1 ),
    .A2(\V4/V2/V2/A3/c2 ),
    .ZN(\V4/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M3/M2/_1_  (.A(\V4/V2/V2/A3/M3/s1 ),
    .B(\V4/V2/V2/A3/c2 ),
    .Z(\V4/V2/v2 [6]));
 OR2_X1 \V4/V2/V2/A3/M3/_0_  (.A1(\V4/V2/V2/A3/M3/c1 ),
    .A2(\V4/V2/V2/A3/M3/c2 ),
    .ZN(\V4/V2/V2/A3/c3 ));
 AND2_X1 \V4/V2/V2/A3/M4/M1/_0_  (.A1(\V4/V2/V2/v4 [3]),
    .A2(ground),
    .ZN(\V4/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M4/M1/_1_  (.A(\V4/V2/V2/v4 [3]),
    .B(ground),
    .Z(\V4/V2/V2/A3/M4/s1 ));
 AND2_X1 \V4/V2/V2/A3/M4/M2/_0_  (.A1(\V4/V2/V2/A3/M4/s1 ),
    .A2(\V4/V2/V2/A3/c3 ),
    .ZN(\V4/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M4/M2/_1_  (.A(\V4/V2/V2/A3/M4/s1 ),
    .B(\V4/V2/V2/A3/c3 ),
    .Z(\V4/V2/v2 [7]));
 OR2_X1 \V4/V2/V2/A3/M4/_0_  (.A1(\V4/V2/V2/A3/M4/c1 ),
    .A2(\V4/V2/V2/A3/M4/c2 ),
    .ZN(\V4/V2/V2/overflow ));
 AND2_X1 \V4/V2/V2/V1/HA1/_0_  (.A1(\V4/V2/V2/V1/w2 ),
    .A2(\V4/V2/V2/V1/w1 ),
    .ZN(\V4/V2/V2/V1/w4 ));
 XOR2_X2 \V4/V2/V2/V1/HA1/_1_  (.A(\V4/V2/V2/V1/w2 ),
    .B(\V4/V2/V2/V1/w1 ),
    .Z(\V4/V2/v2 [1]));
 AND2_X1 \V4/V2/V2/V1/HA2/_0_  (.A1(\V4/V2/V2/V1/w4 ),
    .A2(\V4/V2/V2/V1/w3 ),
    .ZN(\V4/V2/V2/v1 [3]));
 XOR2_X2 \V4/V2/V2/V1/HA2/_1_  (.A(\V4/V2/V2/V1/w4 ),
    .B(\V4/V2/V2/V1/w3 ),
    .Z(\V4/V2/V2/v1 [2]));
 AND2_X1 \V4/V2/V2/V1/_0_  (.A1(A[28]),
    .A2(B[16]),
    .ZN(\V4/V2/v2 [0]));
 AND2_X1 \V4/V2/V2/V1/_1_  (.A1(A[28]),
    .A2(B[17]),
    .ZN(\V4/V2/V2/V1/w1 ));
 AND2_X1 \V4/V2/V2/V1/_2_  (.A1(B[16]),
    .A2(A[29]),
    .ZN(\V4/V2/V2/V1/w2 ));
 AND2_X1 \V4/V2/V2/V1/_3_  (.A1(B[17]),
    .A2(A[29]),
    .ZN(\V4/V2/V2/V1/w3 ));
 AND2_X1 \V4/V2/V2/V2/HA1/_0_  (.A1(\V4/V2/V2/V2/w2 ),
    .A2(\V4/V2/V2/V2/w1 ),
    .ZN(\V4/V2/V2/V2/w4 ));
 XOR2_X2 \V4/V2/V2/V2/HA1/_1_  (.A(\V4/V2/V2/V2/w2 ),
    .B(\V4/V2/V2/V2/w1 ),
    .Z(\V4/V2/V2/v2 [1]));
 AND2_X1 \V4/V2/V2/V2/HA2/_0_  (.A1(\V4/V2/V2/V2/w4 ),
    .A2(\V4/V2/V2/V2/w3 ),
    .ZN(\V4/V2/V2/v2 [3]));
 XOR2_X2 \V4/V2/V2/V2/HA2/_1_  (.A(\V4/V2/V2/V2/w4 ),
    .B(\V4/V2/V2/V2/w3 ),
    .Z(\V4/V2/V2/v2 [2]));
 AND2_X1 \V4/V2/V2/V2/_0_  (.A1(A[30]),
    .A2(B[16]),
    .ZN(\V4/V2/V2/v2 [0]));
 AND2_X1 \V4/V2/V2/V2/_1_  (.A1(A[30]),
    .A2(B[17]),
    .ZN(\V4/V2/V2/V2/w1 ));
 AND2_X1 \V4/V2/V2/V2/_2_  (.A1(B[16]),
    .A2(A[31]),
    .ZN(\V4/V2/V2/V2/w2 ));
 AND2_X1 \V4/V2/V2/V2/_3_  (.A1(B[17]),
    .A2(A[31]),
    .ZN(\V4/V2/V2/V2/w3 ));
 AND2_X1 \V4/V2/V2/V3/HA1/_0_  (.A1(\V4/V2/V2/V3/w2 ),
    .A2(\V4/V2/V2/V3/w1 ),
    .ZN(\V4/V2/V2/V3/w4 ));
 XOR2_X2 \V4/V2/V2/V3/HA1/_1_  (.A(\V4/V2/V2/V3/w2 ),
    .B(\V4/V2/V2/V3/w1 ),
    .Z(\V4/V2/V2/v3 [1]));
 AND2_X1 \V4/V2/V2/V3/HA2/_0_  (.A1(\V4/V2/V2/V3/w4 ),
    .A2(\V4/V2/V2/V3/w3 ),
    .ZN(\V4/V2/V2/v3 [3]));
 XOR2_X2 \V4/V2/V2/V3/HA2/_1_  (.A(\V4/V2/V2/V3/w4 ),
    .B(\V4/V2/V2/V3/w3 ),
    .Z(\V4/V2/V2/v3 [2]));
 AND2_X1 \V4/V2/V2/V3/_0_  (.A1(A[28]),
    .A2(B[18]),
    .ZN(\V4/V2/V2/v3 [0]));
 AND2_X1 \V4/V2/V2/V3/_1_  (.A1(A[28]),
    .A2(B[19]),
    .ZN(\V4/V2/V2/V3/w1 ));
 AND2_X1 \V4/V2/V2/V3/_2_  (.A1(B[18]),
    .A2(A[29]),
    .ZN(\V4/V2/V2/V3/w2 ));
 AND2_X1 \V4/V2/V2/V3/_3_  (.A1(B[19]),
    .A2(A[29]),
    .ZN(\V4/V2/V2/V3/w3 ));
 AND2_X1 \V4/V2/V2/V4/HA1/_0_  (.A1(\V4/V2/V2/V4/w2 ),
    .A2(\V4/V2/V2/V4/w1 ),
    .ZN(\V4/V2/V2/V4/w4 ));
 XOR2_X2 \V4/V2/V2/V4/HA1/_1_  (.A(\V4/V2/V2/V4/w2 ),
    .B(\V4/V2/V2/V4/w1 ),
    .Z(\V4/V2/V2/v4 [1]));
 AND2_X1 \V4/V2/V2/V4/HA2/_0_  (.A1(\V4/V2/V2/V4/w4 ),
    .A2(\V4/V2/V2/V4/w3 ),
    .ZN(\V4/V2/V2/v4 [3]));
 XOR2_X2 \V4/V2/V2/V4/HA2/_1_  (.A(\V4/V2/V2/V4/w4 ),
    .B(\V4/V2/V2/V4/w3 ),
    .Z(\V4/V2/V2/v4 [2]));
 AND2_X1 \V4/V2/V2/V4/_0_  (.A1(A[30]),
    .A2(B[18]),
    .ZN(\V4/V2/V2/v4 [0]));
 AND2_X1 \V4/V2/V2/V4/_1_  (.A1(A[30]),
    .A2(B[19]),
    .ZN(\V4/V2/V2/V4/w1 ));
 AND2_X1 \V4/V2/V2/V4/_2_  (.A1(B[18]),
    .A2(A[31]),
    .ZN(\V4/V2/V2/V4/w2 ));
 AND2_X1 \V4/V2/V2/V4/_3_  (.A1(B[19]),
    .A2(A[31]),
    .ZN(\V4/V2/V2/V4/w3 ));
 OR2_X1 \V4/V2/V2/_0_  (.A1(\V4/V2/V2/c1 ),
    .A2(\V4/V2/V2/c2 ),
    .ZN(\V4/V2/V2/c3 ));
 AND2_X1 \V4/V2/V3/A1/M1/M1/_0_  (.A1(\V4/V2/V3/v2 [0]),
    .A2(\V4/V2/V3/v3 [0]),
    .ZN(\V4/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M1/M1/_1_  (.A(\V4/V2/V3/v2 [0]),
    .B(\V4/V2/V3/v3 [0]),
    .Z(\V4/V2/V3/A1/M1/s1 ));
 AND2_X1 \V4/V2/V3/A1/M1/M2/_0_  (.A1(\V4/V2/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M1/M2/_1_  (.A(\V4/V2/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/V3/s1 [0]));
 OR2_X1 \V4/V2/V3/A1/M1/_0_  (.A1(\V4/V2/V3/A1/M1/c1 ),
    .A2(\V4/V2/V3/A1/M1/c2 ),
    .ZN(\V4/V2/V3/A1/c1 ));
 AND2_X1 \V4/V2/V3/A1/M2/M1/_0_  (.A1(\V4/V2/V3/v2 [1]),
    .A2(\V4/V2/V3/v3 [1]),
    .ZN(\V4/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M2/M1/_1_  (.A(\V4/V2/V3/v2 [1]),
    .B(\V4/V2/V3/v3 [1]),
    .Z(\V4/V2/V3/A1/M2/s1 ));
 AND2_X1 \V4/V2/V3/A1/M2/M2/_0_  (.A1(\V4/V2/V3/A1/M2/s1 ),
    .A2(\V4/V2/V3/A1/c1 ),
    .ZN(\V4/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M2/M2/_1_  (.A(\V4/V2/V3/A1/M2/s1 ),
    .B(\V4/V2/V3/A1/c1 ),
    .Z(\V4/V2/V3/s1 [1]));
 OR2_X1 \V4/V2/V3/A1/M2/_0_  (.A1(\V4/V2/V3/A1/M2/c1 ),
    .A2(\V4/V2/V3/A1/M2/c2 ),
    .ZN(\V4/V2/V3/A1/c2 ));
 AND2_X1 \V4/V2/V3/A1/M3/M1/_0_  (.A1(\V4/V2/V3/v2 [2]),
    .A2(\V4/V2/V3/v3 [2]),
    .ZN(\V4/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M3/M1/_1_  (.A(\V4/V2/V3/v2 [2]),
    .B(\V4/V2/V3/v3 [2]),
    .Z(\V4/V2/V3/A1/M3/s1 ));
 AND2_X1 \V4/V2/V3/A1/M3/M2/_0_  (.A1(\V4/V2/V3/A1/M3/s1 ),
    .A2(\V4/V2/V3/A1/c2 ),
    .ZN(\V4/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M3/M2/_1_  (.A(\V4/V2/V3/A1/M3/s1 ),
    .B(\V4/V2/V3/A1/c2 ),
    .Z(\V4/V2/V3/s1 [2]));
 OR2_X1 \V4/V2/V3/A1/M3/_0_  (.A1(\V4/V2/V3/A1/M3/c1 ),
    .A2(\V4/V2/V3/A1/M3/c2 ),
    .ZN(\V4/V2/V3/A1/c3 ));
 AND2_X1 \V4/V2/V3/A1/M4/M1/_0_  (.A1(\V4/V2/V3/v2 [3]),
    .A2(\V4/V2/V3/v3 [3]),
    .ZN(\V4/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M4/M1/_1_  (.A(\V4/V2/V3/v2 [3]),
    .B(\V4/V2/V3/v3 [3]),
    .Z(\V4/V2/V3/A1/M4/s1 ));
 AND2_X1 \V4/V2/V3/A1/M4/M2/_0_  (.A1(\V4/V2/V3/A1/M4/s1 ),
    .A2(\V4/V2/V3/A1/c3 ),
    .ZN(\V4/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M4/M2/_1_  (.A(\V4/V2/V3/A1/M4/s1 ),
    .B(\V4/V2/V3/A1/c3 ),
    .Z(\V4/V2/V3/s1 [3]));
 OR2_X1 \V4/V2/V3/A1/M4/_0_  (.A1(\V4/V2/V3/A1/M4/c1 ),
    .A2(\V4/V2/V3/A1/M4/c2 ),
    .ZN(\V4/V2/V3/c1 ));
 AND2_X1 \V4/V2/V3/A2/M1/M1/_0_  (.A1(\V4/V2/V3/s1 [0]),
    .A2(\V4/V2/V3/v1 [2]),
    .ZN(\V4/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M1/M1/_1_  (.A(\V4/V2/V3/s1 [0]),
    .B(\V4/V2/V3/v1 [2]),
    .Z(\V4/V2/V3/A2/M1/s1 ));
 AND2_X1 \V4/V2/V3/A2/M1/M2/_0_  (.A1(\V4/V2/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M1/M2/_1_  (.A(\V4/V2/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v3 [2]));
 OR2_X1 \V4/V2/V3/A2/M1/_0_  (.A1(\V4/V2/V3/A2/M1/c1 ),
    .A2(\V4/V2/V3/A2/M1/c2 ),
    .ZN(\V4/V2/V3/A2/c1 ));
 AND2_X1 \V4/V2/V3/A2/M2/M1/_0_  (.A1(\V4/V2/V3/s1 [1]),
    .A2(\V4/V2/V3/v1 [3]),
    .ZN(\V4/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M2/M1/_1_  (.A(\V4/V2/V3/s1 [1]),
    .B(\V4/V2/V3/v1 [3]),
    .Z(\V4/V2/V3/A2/M2/s1 ));
 AND2_X1 \V4/V2/V3/A2/M2/M2/_0_  (.A1(\V4/V2/V3/A2/M2/s1 ),
    .A2(\V4/V2/V3/A2/c1 ),
    .ZN(\V4/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M2/M2/_1_  (.A(\V4/V2/V3/A2/M2/s1 ),
    .B(\V4/V2/V3/A2/c1 ),
    .Z(\V4/V2/v3 [3]));
 OR2_X1 \V4/V2/V3/A2/M2/_0_  (.A1(\V4/V2/V3/A2/M2/c1 ),
    .A2(\V4/V2/V3/A2/M2/c2 ),
    .ZN(\V4/V2/V3/A2/c2 ));
 AND2_X1 \V4/V2/V3/A2/M3/M1/_0_  (.A1(\V4/V2/V3/s1 [2]),
    .A2(ground),
    .ZN(\V4/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M3/M1/_1_  (.A(\V4/V2/V3/s1 [2]),
    .B(ground),
    .Z(\V4/V2/V3/A2/M3/s1 ));
 AND2_X1 \V4/V2/V3/A2/M3/M2/_0_  (.A1(\V4/V2/V3/A2/M3/s1 ),
    .A2(\V4/V2/V3/A2/c2 ),
    .ZN(\V4/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M3/M2/_1_  (.A(\V4/V2/V3/A2/M3/s1 ),
    .B(\V4/V2/V3/A2/c2 ),
    .Z(\V4/V2/V3/s2 [2]));
 OR2_X1 \V4/V2/V3/A2/M3/_0_  (.A1(\V4/V2/V3/A2/M3/c1 ),
    .A2(\V4/V2/V3/A2/M3/c2 ),
    .ZN(\V4/V2/V3/A2/c3 ));
 AND2_X1 \V4/V2/V3/A2/M4/M1/_0_  (.A1(\V4/V2/V3/s1 [3]),
    .A2(ground),
    .ZN(\V4/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M4/M1/_1_  (.A(\V4/V2/V3/s1 [3]),
    .B(ground),
    .Z(\V4/V2/V3/A2/M4/s1 ));
 AND2_X1 \V4/V2/V3/A2/M4/M2/_0_  (.A1(\V4/V2/V3/A2/M4/s1 ),
    .A2(\V4/V2/V3/A2/c3 ),
    .ZN(\V4/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M4/M2/_1_  (.A(\V4/V2/V3/A2/M4/s1 ),
    .B(\V4/V2/V3/A2/c3 ),
    .Z(\V4/V2/V3/s2 [3]));
 OR2_X1 \V4/V2/V3/A2/M4/_0_  (.A1(\V4/V2/V3/A2/M4/c1 ),
    .A2(\V4/V2/V3/A2/M4/c2 ),
    .ZN(\V4/V2/V3/c2 ));
 AND2_X1 \V4/V2/V3/A3/M1/M1/_0_  (.A1(\V4/V2/V3/v4 [0]),
    .A2(\V4/V2/V3/s2 [2]),
    .ZN(\V4/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M1/M1/_1_  (.A(\V4/V2/V3/v4 [0]),
    .B(\V4/V2/V3/s2 [2]),
    .Z(\V4/V2/V3/A3/M1/s1 ));
 AND2_X1 \V4/V2/V3/A3/M1/M2/_0_  (.A1(\V4/V2/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M1/M2/_1_  (.A(\V4/V2/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v3 [4]));
 OR2_X1 \V4/V2/V3/A3/M1/_0_  (.A1(\V4/V2/V3/A3/M1/c1 ),
    .A2(\V4/V2/V3/A3/M1/c2 ),
    .ZN(\V4/V2/V3/A3/c1 ));
 AND2_X1 \V4/V2/V3/A3/M2/M1/_0_  (.A1(\V4/V2/V3/v4 [1]),
    .A2(\V4/V2/V3/s2 [3]),
    .ZN(\V4/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M2/M1/_1_  (.A(\V4/V2/V3/v4 [1]),
    .B(\V4/V2/V3/s2 [3]),
    .Z(\V4/V2/V3/A3/M2/s1 ));
 AND2_X1 \V4/V2/V3/A3/M2/M2/_0_  (.A1(\V4/V2/V3/A3/M2/s1 ),
    .A2(\V4/V2/V3/A3/c1 ),
    .ZN(\V4/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M2/M2/_1_  (.A(\V4/V2/V3/A3/M2/s1 ),
    .B(\V4/V2/V3/A3/c1 ),
    .Z(\V4/V2/v3 [5]));
 OR2_X1 \V4/V2/V3/A3/M2/_0_  (.A1(\V4/V2/V3/A3/M2/c1 ),
    .A2(\V4/V2/V3/A3/M2/c2 ),
    .ZN(\V4/V2/V3/A3/c2 ));
 AND2_X1 \V4/V2/V3/A3/M3/M1/_0_  (.A1(\V4/V2/V3/v4 [2]),
    .A2(\V4/V2/V3/c3 ),
    .ZN(\V4/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M3/M1/_1_  (.A(\V4/V2/V3/v4 [2]),
    .B(\V4/V2/V3/c3 ),
    .Z(\V4/V2/V3/A3/M3/s1 ));
 AND2_X1 \V4/V2/V3/A3/M3/M2/_0_  (.A1(\V4/V2/V3/A3/M3/s1 ),
    .A2(\V4/V2/V3/A3/c2 ),
    .ZN(\V4/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M3/M2/_1_  (.A(\V4/V2/V3/A3/M3/s1 ),
    .B(\V4/V2/V3/A3/c2 ),
    .Z(\V4/V2/v3 [6]));
 OR2_X1 \V4/V2/V3/A3/M3/_0_  (.A1(\V4/V2/V3/A3/M3/c1 ),
    .A2(\V4/V2/V3/A3/M3/c2 ),
    .ZN(\V4/V2/V3/A3/c3 ));
 AND2_X1 \V4/V2/V3/A3/M4/M1/_0_  (.A1(\V4/V2/V3/v4 [3]),
    .A2(ground),
    .ZN(\V4/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M4/M1/_1_  (.A(\V4/V2/V3/v4 [3]),
    .B(ground),
    .Z(\V4/V2/V3/A3/M4/s1 ));
 AND2_X1 \V4/V2/V3/A3/M4/M2/_0_  (.A1(\V4/V2/V3/A3/M4/s1 ),
    .A2(\V4/V2/V3/A3/c3 ),
    .ZN(\V4/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M4/M2/_1_  (.A(\V4/V2/V3/A3/M4/s1 ),
    .B(\V4/V2/V3/A3/c3 ),
    .Z(\V4/V2/v3 [7]));
 OR2_X1 \V4/V2/V3/A3/M4/_0_  (.A1(\V4/V2/V3/A3/M4/c1 ),
    .A2(\V4/V2/V3/A3/M4/c2 ),
    .ZN(\V4/V2/V3/overflow ));
 AND2_X1 \V4/V2/V3/V1/HA1/_0_  (.A1(\V4/V2/V3/V1/w2 ),
    .A2(\V4/V2/V3/V1/w1 ),
    .ZN(\V4/V2/V3/V1/w4 ));
 XOR2_X2 \V4/V2/V3/V1/HA1/_1_  (.A(\V4/V2/V3/V1/w2 ),
    .B(\V4/V2/V3/V1/w1 ),
    .Z(\V4/V2/v3 [1]));
 AND2_X1 \V4/V2/V3/V1/HA2/_0_  (.A1(\V4/V2/V3/V1/w4 ),
    .A2(\V4/V2/V3/V1/w3 ),
    .ZN(\V4/V2/V3/v1 [3]));
 XOR2_X2 \V4/V2/V3/V1/HA2/_1_  (.A(\V4/V2/V3/V1/w4 ),
    .B(\V4/V2/V3/V1/w3 ),
    .Z(\V4/V2/V3/v1 [2]));
 AND2_X1 \V4/V2/V3/V1/_0_  (.A1(A[24]),
    .A2(B[20]),
    .ZN(\V4/V2/v3 [0]));
 AND2_X1 \V4/V2/V3/V1/_1_  (.A1(A[24]),
    .A2(B[21]),
    .ZN(\V4/V2/V3/V1/w1 ));
 AND2_X1 \V4/V2/V3/V1/_2_  (.A1(B[20]),
    .A2(A[25]),
    .ZN(\V4/V2/V3/V1/w2 ));
 AND2_X1 \V4/V2/V3/V1/_3_  (.A1(B[21]),
    .A2(A[25]),
    .ZN(\V4/V2/V3/V1/w3 ));
 AND2_X1 \V4/V2/V3/V2/HA1/_0_  (.A1(\V4/V2/V3/V2/w2 ),
    .A2(\V4/V2/V3/V2/w1 ),
    .ZN(\V4/V2/V3/V2/w4 ));
 XOR2_X2 \V4/V2/V3/V2/HA1/_1_  (.A(\V4/V2/V3/V2/w2 ),
    .B(\V4/V2/V3/V2/w1 ),
    .Z(\V4/V2/V3/v2 [1]));
 AND2_X1 \V4/V2/V3/V2/HA2/_0_  (.A1(\V4/V2/V3/V2/w4 ),
    .A2(\V4/V2/V3/V2/w3 ),
    .ZN(\V4/V2/V3/v2 [3]));
 XOR2_X2 \V4/V2/V3/V2/HA2/_1_  (.A(\V4/V2/V3/V2/w4 ),
    .B(\V4/V2/V3/V2/w3 ),
    .Z(\V4/V2/V3/v2 [2]));
 AND2_X1 \V4/V2/V3/V2/_0_  (.A1(A[26]),
    .A2(B[20]),
    .ZN(\V4/V2/V3/v2 [0]));
 AND2_X1 \V4/V2/V3/V2/_1_  (.A1(A[26]),
    .A2(B[21]),
    .ZN(\V4/V2/V3/V2/w1 ));
 AND2_X1 \V4/V2/V3/V2/_2_  (.A1(B[20]),
    .A2(A[27]),
    .ZN(\V4/V2/V3/V2/w2 ));
 AND2_X1 \V4/V2/V3/V2/_3_  (.A1(B[21]),
    .A2(A[27]),
    .ZN(\V4/V2/V3/V2/w3 ));
 AND2_X1 \V4/V2/V3/V3/HA1/_0_  (.A1(\V4/V2/V3/V3/w2 ),
    .A2(\V4/V2/V3/V3/w1 ),
    .ZN(\V4/V2/V3/V3/w4 ));
 XOR2_X2 \V4/V2/V3/V3/HA1/_1_  (.A(\V4/V2/V3/V3/w2 ),
    .B(\V4/V2/V3/V3/w1 ),
    .Z(\V4/V2/V3/v3 [1]));
 AND2_X1 \V4/V2/V3/V3/HA2/_0_  (.A1(\V4/V2/V3/V3/w4 ),
    .A2(\V4/V2/V3/V3/w3 ),
    .ZN(\V4/V2/V3/v3 [3]));
 XOR2_X2 \V4/V2/V3/V3/HA2/_1_  (.A(\V4/V2/V3/V3/w4 ),
    .B(\V4/V2/V3/V3/w3 ),
    .Z(\V4/V2/V3/v3 [2]));
 AND2_X1 \V4/V2/V3/V3/_0_  (.A1(A[24]),
    .A2(B[22]),
    .ZN(\V4/V2/V3/v3 [0]));
 AND2_X1 \V4/V2/V3/V3/_1_  (.A1(A[24]),
    .A2(B[23]),
    .ZN(\V4/V2/V3/V3/w1 ));
 AND2_X1 \V4/V2/V3/V3/_2_  (.A1(B[22]),
    .A2(A[25]),
    .ZN(\V4/V2/V3/V3/w2 ));
 AND2_X1 \V4/V2/V3/V3/_3_  (.A1(B[23]),
    .A2(A[25]),
    .ZN(\V4/V2/V3/V3/w3 ));
 AND2_X1 \V4/V2/V3/V4/HA1/_0_  (.A1(\V4/V2/V3/V4/w2 ),
    .A2(\V4/V2/V3/V4/w1 ),
    .ZN(\V4/V2/V3/V4/w4 ));
 XOR2_X2 \V4/V2/V3/V4/HA1/_1_  (.A(\V4/V2/V3/V4/w2 ),
    .B(\V4/V2/V3/V4/w1 ),
    .Z(\V4/V2/V3/v4 [1]));
 AND2_X1 \V4/V2/V3/V4/HA2/_0_  (.A1(\V4/V2/V3/V4/w4 ),
    .A2(\V4/V2/V3/V4/w3 ),
    .ZN(\V4/V2/V3/v4 [3]));
 XOR2_X2 \V4/V2/V3/V4/HA2/_1_  (.A(\V4/V2/V3/V4/w4 ),
    .B(\V4/V2/V3/V4/w3 ),
    .Z(\V4/V2/V3/v4 [2]));
 AND2_X1 \V4/V2/V3/V4/_0_  (.A1(A[26]),
    .A2(B[22]),
    .ZN(\V4/V2/V3/v4 [0]));
 AND2_X1 \V4/V2/V3/V4/_1_  (.A1(A[26]),
    .A2(B[23]),
    .ZN(\V4/V2/V3/V4/w1 ));
 AND2_X1 \V4/V2/V3/V4/_2_  (.A1(B[22]),
    .A2(A[27]),
    .ZN(\V4/V2/V3/V4/w2 ));
 AND2_X1 \V4/V2/V3/V4/_3_  (.A1(B[23]),
    .A2(A[27]),
    .ZN(\V4/V2/V3/V4/w3 ));
 OR2_X1 \V4/V2/V3/_0_  (.A1(\V4/V2/V3/c1 ),
    .A2(\V4/V2/V3/c2 ),
    .ZN(\V4/V2/V3/c3 ));
 AND2_X1 \V4/V2/V4/A1/M1/M1/_0_  (.A1(\V4/V2/V4/v2 [0]),
    .A2(\V4/V2/V4/v3 [0]),
    .ZN(\V4/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M1/M1/_1_  (.A(\V4/V2/V4/v2 [0]),
    .B(\V4/V2/V4/v3 [0]),
    .Z(\V4/V2/V4/A1/M1/s1 ));
 AND2_X1 \V4/V2/V4/A1/M1/M2/_0_  (.A1(\V4/V2/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M1/M2/_1_  (.A(\V4/V2/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/V4/s1 [0]));
 OR2_X1 \V4/V2/V4/A1/M1/_0_  (.A1(\V4/V2/V4/A1/M1/c1 ),
    .A2(\V4/V2/V4/A1/M1/c2 ),
    .ZN(\V4/V2/V4/A1/c1 ));
 AND2_X1 \V4/V2/V4/A1/M2/M1/_0_  (.A1(\V4/V2/V4/v2 [1]),
    .A2(\V4/V2/V4/v3 [1]),
    .ZN(\V4/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M2/M1/_1_  (.A(\V4/V2/V4/v2 [1]),
    .B(\V4/V2/V4/v3 [1]),
    .Z(\V4/V2/V4/A1/M2/s1 ));
 AND2_X1 \V4/V2/V4/A1/M2/M2/_0_  (.A1(\V4/V2/V4/A1/M2/s1 ),
    .A2(\V4/V2/V4/A1/c1 ),
    .ZN(\V4/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M2/M2/_1_  (.A(\V4/V2/V4/A1/M2/s1 ),
    .B(\V4/V2/V4/A1/c1 ),
    .Z(\V4/V2/V4/s1 [1]));
 OR2_X1 \V4/V2/V4/A1/M2/_0_  (.A1(\V4/V2/V4/A1/M2/c1 ),
    .A2(\V4/V2/V4/A1/M2/c2 ),
    .ZN(\V4/V2/V4/A1/c2 ));
 AND2_X1 \V4/V2/V4/A1/M3/M1/_0_  (.A1(\V4/V2/V4/v2 [2]),
    .A2(\V4/V2/V4/v3 [2]),
    .ZN(\V4/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M3/M1/_1_  (.A(\V4/V2/V4/v2 [2]),
    .B(\V4/V2/V4/v3 [2]),
    .Z(\V4/V2/V4/A1/M3/s1 ));
 AND2_X1 \V4/V2/V4/A1/M3/M2/_0_  (.A1(\V4/V2/V4/A1/M3/s1 ),
    .A2(\V4/V2/V4/A1/c2 ),
    .ZN(\V4/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M3/M2/_1_  (.A(\V4/V2/V4/A1/M3/s1 ),
    .B(\V4/V2/V4/A1/c2 ),
    .Z(\V4/V2/V4/s1 [2]));
 OR2_X1 \V4/V2/V4/A1/M3/_0_  (.A1(\V4/V2/V4/A1/M3/c1 ),
    .A2(\V4/V2/V4/A1/M3/c2 ),
    .ZN(\V4/V2/V4/A1/c3 ));
 AND2_X1 \V4/V2/V4/A1/M4/M1/_0_  (.A1(\V4/V2/V4/v2 [3]),
    .A2(\V4/V2/V4/v3 [3]),
    .ZN(\V4/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M4/M1/_1_  (.A(\V4/V2/V4/v2 [3]),
    .B(\V4/V2/V4/v3 [3]),
    .Z(\V4/V2/V4/A1/M4/s1 ));
 AND2_X1 \V4/V2/V4/A1/M4/M2/_0_  (.A1(\V4/V2/V4/A1/M4/s1 ),
    .A2(\V4/V2/V4/A1/c3 ),
    .ZN(\V4/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M4/M2/_1_  (.A(\V4/V2/V4/A1/M4/s1 ),
    .B(\V4/V2/V4/A1/c3 ),
    .Z(\V4/V2/V4/s1 [3]));
 OR2_X1 \V4/V2/V4/A1/M4/_0_  (.A1(\V4/V2/V4/A1/M4/c1 ),
    .A2(\V4/V2/V4/A1/M4/c2 ),
    .ZN(\V4/V2/V4/c1 ));
 AND2_X1 \V4/V2/V4/A2/M1/M1/_0_  (.A1(\V4/V2/V4/s1 [0]),
    .A2(\V4/V2/V4/v1 [2]),
    .ZN(\V4/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M1/M1/_1_  (.A(\V4/V2/V4/s1 [0]),
    .B(\V4/V2/V4/v1 [2]),
    .Z(\V4/V2/V4/A2/M1/s1 ));
 AND2_X1 \V4/V2/V4/A2/M1/M2/_0_  (.A1(\V4/V2/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M1/M2/_1_  (.A(\V4/V2/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v4 [2]));
 OR2_X1 \V4/V2/V4/A2/M1/_0_  (.A1(\V4/V2/V4/A2/M1/c1 ),
    .A2(\V4/V2/V4/A2/M1/c2 ),
    .ZN(\V4/V2/V4/A2/c1 ));
 AND2_X1 \V4/V2/V4/A2/M2/M1/_0_  (.A1(\V4/V2/V4/s1 [1]),
    .A2(\V4/V2/V4/v1 [3]),
    .ZN(\V4/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M2/M1/_1_  (.A(\V4/V2/V4/s1 [1]),
    .B(\V4/V2/V4/v1 [3]),
    .Z(\V4/V2/V4/A2/M2/s1 ));
 AND2_X1 \V4/V2/V4/A2/M2/M2/_0_  (.A1(\V4/V2/V4/A2/M2/s1 ),
    .A2(\V4/V2/V4/A2/c1 ),
    .ZN(\V4/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M2/M2/_1_  (.A(\V4/V2/V4/A2/M2/s1 ),
    .B(\V4/V2/V4/A2/c1 ),
    .Z(\V4/V2/v4 [3]));
 OR2_X1 \V4/V2/V4/A2/M2/_0_  (.A1(\V4/V2/V4/A2/M2/c1 ),
    .A2(\V4/V2/V4/A2/M2/c2 ),
    .ZN(\V4/V2/V4/A2/c2 ));
 AND2_X1 \V4/V2/V4/A2/M3/M1/_0_  (.A1(\V4/V2/V4/s1 [2]),
    .A2(ground),
    .ZN(\V4/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M3/M1/_1_  (.A(\V4/V2/V4/s1 [2]),
    .B(ground),
    .Z(\V4/V2/V4/A2/M3/s1 ));
 AND2_X1 \V4/V2/V4/A2/M3/M2/_0_  (.A1(\V4/V2/V4/A2/M3/s1 ),
    .A2(\V4/V2/V4/A2/c2 ),
    .ZN(\V4/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M3/M2/_1_  (.A(\V4/V2/V4/A2/M3/s1 ),
    .B(\V4/V2/V4/A2/c2 ),
    .Z(\V4/V2/V4/s2 [2]));
 OR2_X1 \V4/V2/V4/A2/M3/_0_  (.A1(\V4/V2/V4/A2/M3/c1 ),
    .A2(\V4/V2/V4/A2/M3/c2 ),
    .ZN(\V4/V2/V4/A2/c3 ));
 AND2_X1 \V4/V2/V4/A2/M4/M1/_0_  (.A1(\V4/V2/V4/s1 [3]),
    .A2(ground),
    .ZN(\V4/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M4/M1/_1_  (.A(\V4/V2/V4/s1 [3]),
    .B(ground),
    .Z(\V4/V2/V4/A2/M4/s1 ));
 AND2_X1 \V4/V2/V4/A2/M4/M2/_0_  (.A1(\V4/V2/V4/A2/M4/s1 ),
    .A2(\V4/V2/V4/A2/c3 ),
    .ZN(\V4/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M4/M2/_1_  (.A(\V4/V2/V4/A2/M4/s1 ),
    .B(\V4/V2/V4/A2/c3 ),
    .Z(\V4/V2/V4/s2 [3]));
 OR2_X1 \V4/V2/V4/A2/M4/_0_  (.A1(\V4/V2/V4/A2/M4/c1 ),
    .A2(\V4/V2/V4/A2/M4/c2 ),
    .ZN(\V4/V2/V4/c2 ));
 AND2_X1 \V4/V2/V4/A3/M1/M1/_0_  (.A1(\V4/V2/V4/v4 [0]),
    .A2(\V4/V2/V4/s2 [2]),
    .ZN(\V4/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M1/M1/_1_  (.A(\V4/V2/V4/v4 [0]),
    .B(\V4/V2/V4/s2 [2]),
    .Z(\V4/V2/V4/A3/M1/s1 ));
 AND2_X1 \V4/V2/V4/A3/M1/M2/_0_  (.A1(\V4/V2/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M1/M2/_1_  (.A(\V4/V2/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V2/v4 [4]));
 OR2_X1 \V4/V2/V4/A3/M1/_0_  (.A1(\V4/V2/V4/A3/M1/c1 ),
    .A2(\V4/V2/V4/A3/M1/c2 ),
    .ZN(\V4/V2/V4/A3/c1 ));
 AND2_X1 \V4/V2/V4/A3/M2/M1/_0_  (.A1(\V4/V2/V4/v4 [1]),
    .A2(\V4/V2/V4/s2 [3]),
    .ZN(\V4/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M2/M1/_1_  (.A(\V4/V2/V4/v4 [1]),
    .B(\V4/V2/V4/s2 [3]),
    .Z(\V4/V2/V4/A3/M2/s1 ));
 AND2_X1 \V4/V2/V4/A3/M2/M2/_0_  (.A1(\V4/V2/V4/A3/M2/s1 ),
    .A2(\V4/V2/V4/A3/c1 ),
    .ZN(\V4/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M2/M2/_1_  (.A(\V4/V2/V4/A3/M2/s1 ),
    .B(\V4/V2/V4/A3/c1 ),
    .Z(\V4/V2/v4 [5]));
 OR2_X1 \V4/V2/V4/A3/M2/_0_  (.A1(\V4/V2/V4/A3/M2/c1 ),
    .A2(\V4/V2/V4/A3/M2/c2 ),
    .ZN(\V4/V2/V4/A3/c2 ));
 AND2_X1 \V4/V2/V4/A3/M3/M1/_0_  (.A1(\V4/V2/V4/v4 [2]),
    .A2(\V4/V2/V4/c3 ),
    .ZN(\V4/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M3/M1/_1_  (.A(\V4/V2/V4/v4 [2]),
    .B(\V4/V2/V4/c3 ),
    .Z(\V4/V2/V4/A3/M3/s1 ));
 AND2_X1 \V4/V2/V4/A3/M3/M2/_0_  (.A1(\V4/V2/V4/A3/M3/s1 ),
    .A2(\V4/V2/V4/A3/c2 ),
    .ZN(\V4/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M3/M2/_1_  (.A(\V4/V2/V4/A3/M3/s1 ),
    .B(\V4/V2/V4/A3/c2 ),
    .Z(\V4/V2/v4 [6]));
 OR2_X1 \V4/V2/V4/A3/M3/_0_  (.A1(\V4/V2/V4/A3/M3/c1 ),
    .A2(\V4/V2/V4/A3/M3/c2 ),
    .ZN(\V4/V2/V4/A3/c3 ));
 AND2_X1 \V4/V2/V4/A3/M4/M1/_0_  (.A1(\V4/V2/V4/v4 [3]),
    .A2(ground),
    .ZN(\V4/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M4/M1/_1_  (.A(\V4/V2/V4/v4 [3]),
    .B(ground),
    .Z(\V4/V2/V4/A3/M4/s1 ));
 AND2_X1 \V4/V2/V4/A3/M4/M2/_0_  (.A1(\V4/V2/V4/A3/M4/s1 ),
    .A2(\V4/V2/V4/A3/c3 ),
    .ZN(\V4/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M4/M2/_1_  (.A(\V4/V2/V4/A3/M4/s1 ),
    .B(\V4/V2/V4/A3/c3 ),
    .Z(\V4/V2/v4 [7]));
 OR2_X1 \V4/V2/V4/A3/M4/_0_  (.A1(\V4/V2/V4/A3/M4/c1 ),
    .A2(\V4/V2/V4/A3/M4/c2 ),
    .ZN(\V4/V2/V4/overflow ));
 AND2_X1 \V4/V2/V4/V1/HA1/_0_  (.A1(\V4/V2/V4/V1/w2 ),
    .A2(\V4/V2/V4/V1/w1 ),
    .ZN(\V4/V2/V4/V1/w4 ));
 XOR2_X2 \V4/V2/V4/V1/HA1/_1_  (.A(\V4/V2/V4/V1/w2 ),
    .B(\V4/V2/V4/V1/w1 ),
    .Z(\V4/V2/v4 [1]));
 AND2_X1 \V4/V2/V4/V1/HA2/_0_  (.A1(\V4/V2/V4/V1/w4 ),
    .A2(\V4/V2/V4/V1/w3 ),
    .ZN(\V4/V2/V4/v1 [3]));
 XOR2_X2 \V4/V2/V4/V1/HA2/_1_  (.A(\V4/V2/V4/V1/w4 ),
    .B(\V4/V2/V4/V1/w3 ),
    .Z(\V4/V2/V4/v1 [2]));
 AND2_X1 \V4/V2/V4/V1/_0_  (.A1(A[28]),
    .A2(B[20]),
    .ZN(\V4/V2/v4 [0]));
 AND2_X1 \V4/V2/V4/V1/_1_  (.A1(A[28]),
    .A2(B[21]),
    .ZN(\V4/V2/V4/V1/w1 ));
 AND2_X1 \V4/V2/V4/V1/_2_  (.A1(B[20]),
    .A2(A[29]),
    .ZN(\V4/V2/V4/V1/w2 ));
 AND2_X1 \V4/V2/V4/V1/_3_  (.A1(B[21]),
    .A2(A[29]),
    .ZN(\V4/V2/V4/V1/w3 ));
 AND2_X1 \V4/V2/V4/V2/HA1/_0_  (.A1(\V4/V2/V4/V2/w2 ),
    .A2(\V4/V2/V4/V2/w1 ),
    .ZN(\V4/V2/V4/V2/w4 ));
 XOR2_X2 \V4/V2/V4/V2/HA1/_1_  (.A(\V4/V2/V4/V2/w2 ),
    .B(\V4/V2/V4/V2/w1 ),
    .Z(\V4/V2/V4/v2 [1]));
 AND2_X1 \V4/V2/V4/V2/HA2/_0_  (.A1(\V4/V2/V4/V2/w4 ),
    .A2(\V4/V2/V4/V2/w3 ),
    .ZN(\V4/V2/V4/v2 [3]));
 XOR2_X2 \V4/V2/V4/V2/HA2/_1_  (.A(\V4/V2/V4/V2/w4 ),
    .B(\V4/V2/V4/V2/w3 ),
    .Z(\V4/V2/V4/v2 [2]));
 AND2_X1 \V4/V2/V4/V2/_0_  (.A1(A[30]),
    .A2(B[20]),
    .ZN(\V4/V2/V4/v2 [0]));
 AND2_X1 \V4/V2/V4/V2/_1_  (.A1(A[30]),
    .A2(B[21]),
    .ZN(\V4/V2/V4/V2/w1 ));
 AND2_X1 \V4/V2/V4/V2/_2_  (.A1(B[20]),
    .A2(A[31]),
    .ZN(\V4/V2/V4/V2/w2 ));
 AND2_X1 \V4/V2/V4/V2/_3_  (.A1(B[21]),
    .A2(A[31]),
    .ZN(\V4/V2/V4/V2/w3 ));
 AND2_X1 \V4/V2/V4/V3/HA1/_0_  (.A1(\V4/V2/V4/V3/w2 ),
    .A2(\V4/V2/V4/V3/w1 ),
    .ZN(\V4/V2/V4/V3/w4 ));
 XOR2_X2 \V4/V2/V4/V3/HA1/_1_  (.A(\V4/V2/V4/V3/w2 ),
    .B(\V4/V2/V4/V3/w1 ),
    .Z(\V4/V2/V4/v3 [1]));
 AND2_X1 \V4/V2/V4/V3/HA2/_0_  (.A1(\V4/V2/V4/V3/w4 ),
    .A2(\V4/V2/V4/V3/w3 ),
    .ZN(\V4/V2/V4/v3 [3]));
 XOR2_X2 \V4/V2/V4/V3/HA2/_1_  (.A(\V4/V2/V4/V3/w4 ),
    .B(\V4/V2/V4/V3/w3 ),
    .Z(\V4/V2/V4/v3 [2]));
 AND2_X1 \V4/V2/V4/V3/_0_  (.A1(A[28]),
    .A2(B[22]),
    .ZN(\V4/V2/V4/v3 [0]));
 AND2_X1 \V4/V2/V4/V3/_1_  (.A1(A[28]),
    .A2(B[23]),
    .ZN(\V4/V2/V4/V3/w1 ));
 AND2_X1 \V4/V2/V4/V3/_2_  (.A1(B[22]),
    .A2(A[29]),
    .ZN(\V4/V2/V4/V3/w2 ));
 AND2_X1 \V4/V2/V4/V3/_3_  (.A1(B[23]),
    .A2(A[29]),
    .ZN(\V4/V2/V4/V3/w3 ));
 AND2_X1 \V4/V2/V4/V4/HA1/_0_  (.A1(\V4/V2/V4/V4/w2 ),
    .A2(\V4/V2/V4/V4/w1 ),
    .ZN(\V4/V2/V4/V4/w4 ));
 XOR2_X2 \V4/V2/V4/V4/HA1/_1_  (.A(\V4/V2/V4/V4/w2 ),
    .B(\V4/V2/V4/V4/w1 ),
    .Z(\V4/V2/V4/v4 [1]));
 AND2_X1 \V4/V2/V4/V4/HA2/_0_  (.A1(\V4/V2/V4/V4/w4 ),
    .A2(\V4/V2/V4/V4/w3 ),
    .ZN(\V4/V2/V4/v4 [3]));
 XOR2_X2 \V4/V2/V4/V4/HA2/_1_  (.A(\V4/V2/V4/V4/w4 ),
    .B(\V4/V2/V4/V4/w3 ),
    .Z(\V4/V2/V4/v4 [2]));
 AND2_X1 \V4/V2/V4/V4/_0_  (.A1(A[30]),
    .A2(B[22]),
    .ZN(\V4/V2/V4/v4 [0]));
 AND2_X1 \V4/V2/V4/V4/_1_  (.A1(A[30]),
    .A2(B[23]),
    .ZN(\V4/V2/V4/V4/w1 ));
 AND2_X1 \V4/V2/V4/V4/_2_  (.A1(B[22]),
    .A2(A[31]),
    .ZN(\V4/V2/V4/V4/w2 ));
 AND2_X1 \V4/V2/V4/V4/_3_  (.A1(B[23]),
    .A2(A[31]),
    .ZN(\V4/V2/V4/V4/w3 ));
 OR2_X1 \V4/V2/V4/_0_  (.A1(\V4/V2/V4/c1 ),
    .A2(\V4/V2/V4/c2 ),
    .ZN(\V4/V2/V4/c3 ));
 OR2_X1 \V4/V2/_0_  (.A1(\V4/V2/c1 ),
    .A2(\V4/V2/c2 ),
    .ZN(\V4/V2/c3 ));
 AND2_X1 \V4/V3/A1/A1/M1/M1/_0_  (.A1(\V4/V3/v2 [0]),
    .A2(\V4/V3/v3 [0]),
    .ZN(\V4/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M1/M1/_1_  (.A(\V4/V3/v2 [0]),
    .B(\V4/V3/v3 [0]),
    .Z(\V4/V3/A1/A1/M1/s1 ));
 AND2_X1 \V4/V3/A1/A1/M1/M2/_0_  (.A1(\V4/V3/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M1/M2/_1_  (.A(\V4/V3/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/s1 [0]));
 OR2_X1 \V4/V3/A1/A1/M1/_0_  (.A1(\V4/V3/A1/A1/M1/c1 ),
    .A2(\V4/V3/A1/A1/M1/c2 ),
    .ZN(\V4/V3/A1/A1/c1 ));
 AND2_X1 \V4/V3/A1/A1/M2/M1/_0_  (.A1(\V4/V3/v2 [1]),
    .A2(\V4/V3/v3 [1]),
    .ZN(\V4/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M2/M1/_1_  (.A(\V4/V3/v2 [1]),
    .B(\V4/V3/v3 [1]),
    .Z(\V4/V3/A1/A1/M2/s1 ));
 AND2_X1 \V4/V3/A1/A1/M2/M2/_0_  (.A1(\V4/V3/A1/A1/M2/s1 ),
    .A2(\V4/V3/A1/A1/c1 ),
    .ZN(\V4/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M2/M2/_1_  (.A(\V4/V3/A1/A1/M2/s1 ),
    .B(\V4/V3/A1/A1/c1 ),
    .Z(\V4/V3/s1 [1]));
 OR2_X1 \V4/V3/A1/A1/M2/_0_  (.A1(\V4/V3/A1/A1/M2/c1 ),
    .A2(\V4/V3/A1/A1/M2/c2 ),
    .ZN(\V4/V3/A1/A1/c2 ));
 AND2_X1 \V4/V3/A1/A1/M3/M1/_0_  (.A1(\V4/V3/v2 [2]),
    .A2(\V4/V3/v3 [2]),
    .ZN(\V4/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M3/M1/_1_  (.A(\V4/V3/v2 [2]),
    .B(\V4/V3/v3 [2]),
    .Z(\V4/V3/A1/A1/M3/s1 ));
 AND2_X1 \V4/V3/A1/A1/M3/M2/_0_  (.A1(\V4/V3/A1/A1/M3/s1 ),
    .A2(\V4/V3/A1/A1/c2 ),
    .ZN(\V4/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M3/M2/_1_  (.A(\V4/V3/A1/A1/M3/s1 ),
    .B(\V4/V3/A1/A1/c2 ),
    .Z(\V4/V3/s1 [2]));
 OR2_X1 \V4/V3/A1/A1/M3/_0_  (.A1(\V4/V3/A1/A1/M3/c1 ),
    .A2(\V4/V3/A1/A1/M3/c2 ),
    .ZN(\V4/V3/A1/A1/c3 ));
 AND2_X1 \V4/V3/A1/A1/M4/M1/_0_  (.A1(\V4/V3/v2 [3]),
    .A2(\V4/V3/v3 [3]),
    .ZN(\V4/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M4/M1/_1_  (.A(\V4/V3/v2 [3]),
    .B(\V4/V3/v3 [3]),
    .Z(\V4/V3/A1/A1/M4/s1 ));
 AND2_X1 \V4/V3/A1/A1/M4/M2/_0_  (.A1(\V4/V3/A1/A1/M4/s1 ),
    .A2(\V4/V3/A1/A1/c3 ),
    .ZN(\V4/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M4/M2/_1_  (.A(\V4/V3/A1/A1/M4/s1 ),
    .B(\V4/V3/A1/A1/c3 ),
    .Z(\V4/V3/s1 [3]));
 OR2_X1 \V4/V3/A1/A1/M4/_0_  (.A1(\V4/V3/A1/A1/M4/c1 ),
    .A2(\V4/V3/A1/A1/M4/c2 ),
    .ZN(\V4/V3/A1/c1 ));
 AND2_X1 \V4/V3/A1/A2/M1/M1/_0_  (.A1(\V4/V3/v2 [4]),
    .A2(\V4/V3/v3 [4]),
    .ZN(\V4/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M1/M1/_1_  (.A(\V4/V3/v2 [4]),
    .B(\V4/V3/v3 [4]),
    .Z(\V4/V3/A1/A2/M1/s1 ));
 AND2_X1 \V4/V3/A1/A2/M1/M2/_0_  (.A1(\V4/V3/A1/A2/M1/s1 ),
    .A2(\V4/V3/A1/c1 ),
    .ZN(\V4/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M1/M2/_1_  (.A(\V4/V3/A1/A2/M1/s1 ),
    .B(\V4/V3/A1/c1 ),
    .Z(\V4/V3/s1 [4]));
 OR2_X1 \V4/V3/A1/A2/M1/_0_  (.A1(\V4/V3/A1/A2/M1/c1 ),
    .A2(\V4/V3/A1/A2/M1/c2 ),
    .ZN(\V4/V3/A1/A2/c1 ));
 AND2_X1 \V4/V3/A1/A2/M2/M1/_0_  (.A1(\V4/V3/v2 [5]),
    .A2(\V4/V3/v3 [5]),
    .ZN(\V4/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M2/M1/_1_  (.A(\V4/V3/v2 [5]),
    .B(\V4/V3/v3 [5]),
    .Z(\V4/V3/A1/A2/M2/s1 ));
 AND2_X1 \V4/V3/A1/A2/M2/M2/_0_  (.A1(\V4/V3/A1/A2/M2/s1 ),
    .A2(\V4/V3/A1/A2/c1 ),
    .ZN(\V4/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M2/M2/_1_  (.A(\V4/V3/A1/A2/M2/s1 ),
    .B(\V4/V3/A1/A2/c1 ),
    .Z(\V4/V3/s1 [5]));
 OR2_X1 \V4/V3/A1/A2/M2/_0_  (.A1(\V4/V3/A1/A2/M2/c1 ),
    .A2(\V4/V3/A1/A2/M2/c2 ),
    .ZN(\V4/V3/A1/A2/c2 ));
 AND2_X1 \V4/V3/A1/A2/M3/M1/_0_  (.A1(\V4/V3/v2 [6]),
    .A2(\V4/V3/v3 [6]),
    .ZN(\V4/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M3/M1/_1_  (.A(\V4/V3/v2 [6]),
    .B(\V4/V3/v3 [6]),
    .Z(\V4/V3/A1/A2/M3/s1 ));
 AND2_X1 \V4/V3/A1/A2/M3/M2/_0_  (.A1(\V4/V3/A1/A2/M3/s1 ),
    .A2(\V4/V3/A1/A2/c2 ),
    .ZN(\V4/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M3/M2/_1_  (.A(\V4/V3/A1/A2/M3/s1 ),
    .B(\V4/V3/A1/A2/c2 ),
    .Z(\V4/V3/s1 [6]));
 OR2_X1 \V4/V3/A1/A2/M3/_0_  (.A1(\V4/V3/A1/A2/M3/c1 ),
    .A2(\V4/V3/A1/A2/M3/c2 ),
    .ZN(\V4/V3/A1/A2/c3 ));
 AND2_X1 \V4/V3/A1/A2/M4/M1/_0_  (.A1(\V4/V3/v2 [7]),
    .A2(\V4/V3/v3 [7]),
    .ZN(\V4/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M4/M1/_1_  (.A(\V4/V3/v2 [7]),
    .B(\V4/V3/v3 [7]),
    .Z(\V4/V3/A1/A2/M4/s1 ));
 AND2_X1 \V4/V3/A1/A2/M4/M2/_0_  (.A1(\V4/V3/A1/A2/M4/s1 ),
    .A2(\V4/V3/A1/A2/c3 ),
    .ZN(\V4/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M4/M2/_1_  (.A(\V4/V3/A1/A2/M4/s1 ),
    .B(\V4/V3/A1/A2/c3 ),
    .Z(\V4/V3/s1 [7]));
 OR2_X1 \V4/V3/A1/A2/M4/_0_  (.A1(\V4/V3/A1/A2/M4/c1 ),
    .A2(\V4/V3/A1/A2/M4/c2 ),
    .ZN(\V4/V3/c1 ));
 AND2_X1 \V4/V3/A2/A1/M1/M1/_0_  (.A1(\V4/V3/s1 [0]),
    .A2(\V4/V3/v1 [4]),
    .ZN(\V4/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M1/M1/_1_  (.A(\V4/V3/s1 [0]),
    .B(\V4/V3/v1 [4]),
    .Z(\V4/V3/A2/A1/M1/s1 ));
 AND2_X1 \V4/V3/A2/A1/M1/M2/_0_  (.A1(\V4/V3/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M1/M2/_1_  (.A(\V4/V3/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v3 [4]));
 OR2_X1 \V4/V3/A2/A1/M1/_0_  (.A1(\V4/V3/A2/A1/M1/c1 ),
    .A2(\V4/V3/A2/A1/M1/c2 ),
    .ZN(\V4/V3/A2/A1/c1 ));
 AND2_X1 \V4/V3/A2/A1/M2/M1/_0_  (.A1(\V4/V3/s1 [1]),
    .A2(\V4/V3/v1 [5]),
    .ZN(\V4/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M2/M1/_1_  (.A(\V4/V3/s1 [1]),
    .B(\V4/V3/v1 [5]),
    .Z(\V4/V3/A2/A1/M2/s1 ));
 AND2_X1 \V4/V3/A2/A1/M2/M2/_0_  (.A1(\V4/V3/A2/A1/M2/s1 ),
    .A2(\V4/V3/A2/A1/c1 ),
    .ZN(\V4/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M2/M2/_1_  (.A(\V4/V3/A2/A1/M2/s1 ),
    .B(\V4/V3/A2/A1/c1 ),
    .Z(\V4/v3 [5]));
 OR2_X1 \V4/V3/A2/A1/M2/_0_  (.A1(\V4/V3/A2/A1/M2/c1 ),
    .A2(\V4/V3/A2/A1/M2/c2 ),
    .ZN(\V4/V3/A2/A1/c2 ));
 AND2_X1 \V4/V3/A2/A1/M3/M1/_0_  (.A1(\V4/V3/s1 [2]),
    .A2(\V4/V3/v1 [6]),
    .ZN(\V4/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M3/M1/_1_  (.A(\V4/V3/s1 [2]),
    .B(\V4/V3/v1 [6]),
    .Z(\V4/V3/A2/A1/M3/s1 ));
 AND2_X1 \V4/V3/A2/A1/M3/M2/_0_  (.A1(\V4/V3/A2/A1/M3/s1 ),
    .A2(\V4/V3/A2/A1/c2 ),
    .ZN(\V4/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M3/M2/_1_  (.A(\V4/V3/A2/A1/M3/s1 ),
    .B(\V4/V3/A2/A1/c2 ),
    .Z(\V4/v3 [6]));
 OR2_X1 \V4/V3/A2/A1/M3/_0_  (.A1(\V4/V3/A2/A1/M3/c1 ),
    .A2(\V4/V3/A2/A1/M3/c2 ),
    .ZN(\V4/V3/A2/A1/c3 ));
 AND2_X1 \V4/V3/A2/A1/M4/M1/_0_  (.A1(\V4/V3/s1 [3]),
    .A2(\V4/V3/v1 [7]),
    .ZN(\V4/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M4/M1/_1_  (.A(\V4/V3/s1 [3]),
    .B(\V4/V3/v1 [7]),
    .Z(\V4/V3/A2/A1/M4/s1 ));
 AND2_X1 \V4/V3/A2/A1/M4/M2/_0_  (.A1(\V4/V3/A2/A1/M4/s1 ),
    .A2(\V4/V3/A2/A1/c3 ),
    .ZN(\V4/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M4/M2/_1_  (.A(\V4/V3/A2/A1/M4/s1 ),
    .B(\V4/V3/A2/A1/c3 ),
    .Z(\V4/v3 [7]));
 OR2_X1 \V4/V3/A2/A1/M4/_0_  (.A1(\V4/V3/A2/A1/M4/c1 ),
    .A2(\V4/V3/A2/A1/M4/c2 ),
    .ZN(\V4/V3/A2/c1 ));
 AND2_X1 \V4/V3/A2/A2/M1/M1/_0_  (.A1(\V4/V3/s1 [4]),
    .A2(ground),
    .ZN(\V4/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M1/M1/_1_  (.A(\V4/V3/s1 [4]),
    .B(ground),
    .Z(\V4/V3/A2/A2/M1/s1 ));
 AND2_X1 \V4/V3/A2/A2/M1/M2/_0_  (.A1(\V4/V3/A2/A2/M1/s1 ),
    .A2(\V4/V3/A2/c1 ),
    .ZN(\V4/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M1/M2/_1_  (.A(\V4/V3/A2/A2/M1/s1 ),
    .B(\V4/V3/A2/c1 ),
    .Z(\V4/V3/s2 [4]));
 OR2_X1 \V4/V3/A2/A2/M1/_0_  (.A1(\V4/V3/A2/A2/M1/c1 ),
    .A2(\V4/V3/A2/A2/M1/c2 ),
    .ZN(\V4/V3/A2/A2/c1 ));
 AND2_X1 \V4/V3/A2/A2/M2/M1/_0_  (.A1(\V4/V3/s1 [5]),
    .A2(ground),
    .ZN(\V4/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M2/M1/_1_  (.A(\V4/V3/s1 [5]),
    .B(ground),
    .Z(\V4/V3/A2/A2/M2/s1 ));
 AND2_X1 \V4/V3/A2/A2/M2/M2/_0_  (.A1(\V4/V3/A2/A2/M2/s1 ),
    .A2(\V4/V3/A2/A2/c1 ),
    .ZN(\V4/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M2/M2/_1_  (.A(\V4/V3/A2/A2/M2/s1 ),
    .B(\V4/V3/A2/A2/c1 ),
    .Z(\V4/V3/s2 [5]));
 OR2_X1 \V4/V3/A2/A2/M2/_0_  (.A1(\V4/V3/A2/A2/M2/c1 ),
    .A2(\V4/V3/A2/A2/M2/c2 ),
    .ZN(\V4/V3/A2/A2/c2 ));
 AND2_X1 \V4/V3/A2/A2/M3/M1/_0_  (.A1(\V4/V3/s1 [6]),
    .A2(ground),
    .ZN(\V4/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M3/M1/_1_  (.A(\V4/V3/s1 [6]),
    .B(ground),
    .Z(\V4/V3/A2/A2/M3/s1 ));
 AND2_X1 \V4/V3/A2/A2/M3/M2/_0_  (.A1(\V4/V3/A2/A2/M3/s1 ),
    .A2(\V4/V3/A2/A2/c2 ),
    .ZN(\V4/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M3/M2/_1_  (.A(\V4/V3/A2/A2/M3/s1 ),
    .B(\V4/V3/A2/A2/c2 ),
    .Z(\V4/V3/s2 [6]));
 OR2_X1 \V4/V3/A2/A2/M3/_0_  (.A1(\V4/V3/A2/A2/M3/c1 ),
    .A2(\V4/V3/A2/A2/M3/c2 ),
    .ZN(\V4/V3/A2/A2/c3 ));
 AND2_X1 \V4/V3/A2/A2/M4/M1/_0_  (.A1(\V4/V3/s1 [7]),
    .A2(ground),
    .ZN(\V4/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M4/M1/_1_  (.A(\V4/V3/s1 [7]),
    .B(ground),
    .Z(\V4/V3/A2/A2/M4/s1 ));
 AND2_X1 \V4/V3/A2/A2/M4/M2/_0_  (.A1(\V4/V3/A2/A2/M4/s1 ),
    .A2(\V4/V3/A2/A2/c3 ),
    .ZN(\V4/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M4/M2/_1_  (.A(\V4/V3/A2/A2/M4/s1 ),
    .B(\V4/V3/A2/A2/c3 ),
    .Z(\V4/V3/s2 [7]));
 OR2_X1 \V4/V3/A2/A2/M4/_0_  (.A1(\V4/V3/A2/A2/M4/c1 ),
    .A2(\V4/V3/A2/A2/M4/c2 ),
    .ZN(\V4/V3/c2 ));
 AND2_X1 \V4/V3/A3/A1/M1/M1/_0_  (.A1(\V4/V3/v4 [0]),
    .A2(\V4/V3/s2 [4]),
    .ZN(\V4/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M1/M1/_1_  (.A(\V4/V3/v4 [0]),
    .B(\V4/V3/s2 [4]),
    .Z(\V4/V3/A3/A1/M1/s1 ));
 AND2_X1 \V4/V3/A3/A1/M1/M2/_0_  (.A1(\V4/V3/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M1/M2/_1_  (.A(\V4/V3/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v3 [8]));
 OR2_X1 \V4/V3/A3/A1/M1/_0_  (.A1(\V4/V3/A3/A1/M1/c1 ),
    .A2(\V4/V3/A3/A1/M1/c2 ),
    .ZN(\V4/V3/A3/A1/c1 ));
 AND2_X1 \V4/V3/A3/A1/M2/M1/_0_  (.A1(\V4/V3/v4 [1]),
    .A2(\V4/V3/s2 [5]),
    .ZN(\V4/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M2/M1/_1_  (.A(\V4/V3/v4 [1]),
    .B(\V4/V3/s2 [5]),
    .Z(\V4/V3/A3/A1/M2/s1 ));
 AND2_X1 \V4/V3/A3/A1/M2/M2/_0_  (.A1(\V4/V3/A3/A1/M2/s1 ),
    .A2(\V4/V3/A3/A1/c1 ),
    .ZN(\V4/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M2/M2/_1_  (.A(\V4/V3/A3/A1/M2/s1 ),
    .B(\V4/V3/A3/A1/c1 ),
    .Z(\V4/v3 [9]));
 OR2_X1 \V4/V3/A3/A1/M2/_0_  (.A1(\V4/V3/A3/A1/M2/c1 ),
    .A2(\V4/V3/A3/A1/M2/c2 ),
    .ZN(\V4/V3/A3/A1/c2 ));
 AND2_X1 \V4/V3/A3/A1/M3/M1/_0_  (.A1(\V4/V3/v4 [2]),
    .A2(\V4/V3/s2 [6]),
    .ZN(\V4/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M3/M1/_1_  (.A(\V4/V3/v4 [2]),
    .B(\V4/V3/s2 [6]),
    .Z(\V4/V3/A3/A1/M3/s1 ));
 AND2_X1 \V4/V3/A3/A1/M3/M2/_0_  (.A1(\V4/V3/A3/A1/M3/s1 ),
    .A2(\V4/V3/A3/A1/c2 ),
    .ZN(\V4/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M3/M2/_1_  (.A(\V4/V3/A3/A1/M3/s1 ),
    .B(\V4/V3/A3/A1/c2 ),
    .Z(\V4/v3 [10]));
 OR2_X1 \V4/V3/A3/A1/M3/_0_  (.A1(\V4/V3/A3/A1/M3/c1 ),
    .A2(\V4/V3/A3/A1/M3/c2 ),
    .ZN(\V4/V3/A3/A1/c3 ));
 AND2_X1 \V4/V3/A3/A1/M4/M1/_0_  (.A1(\V4/V3/v4 [3]),
    .A2(\V4/V3/s2 [7]),
    .ZN(\V4/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M4/M1/_1_  (.A(\V4/V3/v4 [3]),
    .B(\V4/V3/s2 [7]),
    .Z(\V4/V3/A3/A1/M4/s1 ));
 AND2_X1 \V4/V3/A3/A1/M4/M2/_0_  (.A1(\V4/V3/A3/A1/M4/s1 ),
    .A2(\V4/V3/A3/A1/c3 ),
    .ZN(\V4/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M4/M2/_1_  (.A(\V4/V3/A3/A1/M4/s1 ),
    .B(\V4/V3/A3/A1/c3 ),
    .Z(\V4/v3 [11]));
 OR2_X1 \V4/V3/A3/A1/M4/_0_  (.A1(\V4/V3/A3/A1/M4/c1 ),
    .A2(\V4/V3/A3/A1/M4/c2 ),
    .ZN(\V4/V3/A3/c1 ));
 AND2_X1 \V4/V3/A3/A2/M1/M1/_0_  (.A1(\V4/V3/v4 [4]),
    .A2(\V4/V3/c3 ),
    .ZN(\V4/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M1/M1/_1_  (.A(\V4/V3/v4 [4]),
    .B(\V4/V3/c3 ),
    .Z(\V4/V3/A3/A2/M1/s1 ));
 AND2_X1 \V4/V3/A3/A2/M1/M2/_0_  (.A1(\V4/V3/A3/A2/M1/s1 ),
    .A2(\V4/V3/A3/c1 ),
    .ZN(\V4/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M1/M2/_1_  (.A(\V4/V3/A3/A2/M1/s1 ),
    .B(\V4/V3/A3/c1 ),
    .Z(\V4/v3 [12]));
 OR2_X1 \V4/V3/A3/A2/M1/_0_  (.A1(\V4/V3/A3/A2/M1/c1 ),
    .A2(\V4/V3/A3/A2/M1/c2 ),
    .ZN(\V4/V3/A3/A2/c1 ));
 AND2_X1 \V4/V3/A3/A2/M2/M1/_0_  (.A1(\V4/V3/v4 [5]),
    .A2(ground),
    .ZN(\V4/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M2/M1/_1_  (.A(\V4/V3/v4 [5]),
    .B(ground),
    .Z(\V4/V3/A3/A2/M2/s1 ));
 AND2_X1 \V4/V3/A3/A2/M2/M2/_0_  (.A1(\V4/V3/A3/A2/M2/s1 ),
    .A2(\V4/V3/A3/A2/c1 ),
    .ZN(\V4/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M2/M2/_1_  (.A(\V4/V3/A3/A2/M2/s1 ),
    .B(\V4/V3/A3/A2/c1 ),
    .Z(\V4/v3 [13]));
 OR2_X1 \V4/V3/A3/A2/M2/_0_  (.A1(\V4/V3/A3/A2/M2/c1 ),
    .A2(\V4/V3/A3/A2/M2/c2 ),
    .ZN(\V4/V3/A3/A2/c2 ));
 AND2_X1 \V4/V3/A3/A2/M3/M1/_0_  (.A1(\V4/V3/v4 [6]),
    .A2(ground),
    .ZN(\V4/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M3/M1/_1_  (.A(\V4/V3/v4 [6]),
    .B(ground),
    .Z(\V4/V3/A3/A2/M3/s1 ));
 AND2_X1 \V4/V3/A3/A2/M3/M2/_0_  (.A1(\V4/V3/A3/A2/M3/s1 ),
    .A2(\V4/V3/A3/A2/c2 ),
    .ZN(\V4/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M3/M2/_1_  (.A(\V4/V3/A3/A2/M3/s1 ),
    .B(\V4/V3/A3/A2/c2 ),
    .Z(\V4/v3 [14]));
 OR2_X1 \V4/V3/A3/A2/M3/_0_  (.A1(\V4/V3/A3/A2/M3/c1 ),
    .A2(\V4/V3/A3/A2/M3/c2 ),
    .ZN(\V4/V3/A3/A2/c3 ));
 AND2_X1 \V4/V3/A3/A2/M4/M1/_0_  (.A1(\V4/V3/v4 [7]),
    .A2(ground),
    .ZN(\V4/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M4/M1/_1_  (.A(\V4/V3/v4 [7]),
    .B(ground),
    .Z(\V4/V3/A3/A2/M4/s1 ));
 AND2_X1 \V4/V3/A3/A2/M4/M2/_0_  (.A1(\V4/V3/A3/A2/M4/s1 ),
    .A2(\V4/V3/A3/A2/c3 ),
    .ZN(\V4/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M4/M2/_1_  (.A(\V4/V3/A3/A2/M4/s1 ),
    .B(\V4/V3/A3/A2/c3 ),
    .Z(\V4/v3 [15]));
 OR2_X1 \V4/V3/A3/A2/M4/_0_  (.A1(\V4/V3/A3/A2/M4/c1 ),
    .A2(\V4/V3/A3/A2/M4/c2 ),
    .ZN(\V4/V3/overflow ));
 AND2_X1 \V4/V3/V1/A1/M1/M1/_0_  (.A1(\V4/V3/V1/v2 [0]),
    .A2(\V4/V3/V1/v3 [0]),
    .ZN(\V4/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M1/M1/_1_  (.A(\V4/V3/V1/v2 [0]),
    .B(\V4/V3/V1/v3 [0]),
    .Z(\V4/V3/V1/A1/M1/s1 ));
 AND2_X1 \V4/V3/V1/A1/M1/M2/_0_  (.A1(\V4/V3/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M1/M2/_1_  (.A(\V4/V3/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/V1/s1 [0]));
 OR2_X1 \V4/V3/V1/A1/M1/_0_  (.A1(\V4/V3/V1/A1/M1/c1 ),
    .A2(\V4/V3/V1/A1/M1/c2 ),
    .ZN(\V4/V3/V1/A1/c1 ));
 AND2_X1 \V4/V3/V1/A1/M2/M1/_0_  (.A1(\V4/V3/V1/v2 [1]),
    .A2(\V4/V3/V1/v3 [1]),
    .ZN(\V4/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M2/M1/_1_  (.A(\V4/V3/V1/v2 [1]),
    .B(\V4/V3/V1/v3 [1]),
    .Z(\V4/V3/V1/A1/M2/s1 ));
 AND2_X1 \V4/V3/V1/A1/M2/M2/_0_  (.A1(\V4/V3/V1/A1/M2/s1 ),
    .A2(\V4/V3/V1/A1/c1 ),
    .ZN(\V4/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M2/M2/_1_  (.A(\V4/V3/V1/A1/M2/s1 ),
    .B(\V4/V3/V1/A1/c1 ),
    .Z(\V4/V3/V1/s1 [1]));
 OR2_X1 \V4/V3/V1/A1/M2/_0_  (.A1(\V4/V3/V1/A1/M2/c1 ),
    .A2(\V4/V3/V1/A1/M2/c2 ),
    .ZN(\V4/V3/V1/A1/c2 ));
 AND2_X1 \V4/V3/V1/A1/M3/M1/_0_  (.A1(\V4/V3/V1/v2 [2]),
    .A2(\V4/V3/V1/v3 [2]),
    .ZN(\V4/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M3/M1/_1_  (.A(\V4/V3/V1/v2 [2]),
    .B(\V4/V3/V1/v3 [2]),
    .Z(\V4/V3/V1/A1/M3/s1 ));
 AND2_X1 \V4/V3/V1/A1/M3/M2/_0_  (.A1(\V4/V3/V1/A1/M3/s1 ),
    .A2(\V4/V3/V1/A1/c2 ),
    .ZN(\V4/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M3/M2/_1_  (.A(\V4/V3/V1/A1/M3/s1 ),
    .B(\V4/V3/V1/A1/c2 ),
    .Z(\V4/V3/V1/s1 [2]));
 OR2_X1 \V4/V3/V1/A1/M3/_0_  (.A1(\V4/V3/V1/A1/M3/c1 ),
    .A2(\V4/V3/V1/A1/M3/c2 ),
    .ZN(\V4/V3/V1/A1/c3 ));
 AND2_X1 \V4/V3/V1/A1/M4/M1/_0_  (.A1(\V4/V3/V1/v2 [3]),
    .A2(\V4/V3/V1/v3 [3]),
    .ZN(\V4/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M4/M1/_1_  (.A(\V4/V3/V1/v2 [3]),
    .B(\V4/V3/V1/v3 [3]),
    .Z(\V4/V3/V1/A1/M4/s1 ));
 AND2_X1 \V4/V3/V1/A1/M4/M2/_0_  (.A1(\V4/V3/V1/A1/M4/s1 ),
    .A2(\V4/V3/V1/A1/c3 ),
    .ZN(\V4/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M4/M2/_1_  (.A(\V4/V3/V1/A1/M4/s1 ),
    .B(\V4/V3/V1/A1/c3 ),
    .Z(\V4/V3/V1/s1 [3]));
 OR2_X1 \V4/V3/V1/A1/M4/_0_  (.A1(\V4/V3/V1/A1/M4/c1 ),
    .A2(\V4/V3/V1/A1/M4/c2 ),
    .ZN(\V4/V3/V1/c1 ));
 AND2_X1 \V4/V3/V1/A2/M1/M1/_0_  (.A1(\V4/V3/V1/s1 [0]),
    .A2(\V4/V3/V1/v1 [2]),
    .ZN(\V4/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M1/M1/_1_  (.A(\V4/V3/V1/s1 [0]),
    .B(\V4/V3/V1/v1 [2]),
    .Z(\V4/V3/V1/A2/M1/s1 ));
 AND2_X1 \V4/V3/V1/A2/M1/M2/_0_  (.A1(\V4/V3/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M1/M2/_1_  (.A(\V4/V3/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/v3 [2]));
 OR2_X1 \V4/V3/V1/A2/M1/_0_  (.A1(\V4/V3/V1/A2/M1/c1 ),
    .A2(\V4/V3/V1/A2/M1/c2 ),
    .ZN(\V4/V3/V1/A2/c1 ));
 AND2_X1 \V4/V3/V1/A2/M2/M1/_0_  (.A1(\V4/V3/V1/s1 [1]),
    .A2(\V4/V3/V1/v1 [3]),
    .ZN(\V4/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M2/M1/_1_  (.A(\V4/V3/V1/s1 [1]),
    .B(\V4/V3/V1/v1 [3]),
    .Z(\V4/V3/V1/A2/M2/s1 ));
 AND2_X1 \V4/V3/V1/A2/M2/M2/_0_  (.A1(\V4/V3/V1/A2/M2/s1 ),
    .A2(\V4/V3/V1/A2/c1 ),
    .ZN(\V4/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M2/M2/_1_  (.A(\V4/V3/V1/A2/M2/s1 ),
    .B(\V4/V3/V1/A2/c1 ),
    .Z(\V4/v3 [3]));
 OR2_X1 \V4/V3/V1/A2/M2/_0_  (.A1(\V4/V3/V1/A2/M2/c1 ),
    .A2(\V4/V3/V1/A2/M2/c2 ),
    .ZN(\V4/V3/V1/A2/c2 ));
 AND2_X1 \V4/V3/V1/A2/M3/M1/_0_  (.A1(\V4/V3/V1/s1 [2]),
    .A2(ground),
    .ZN(\V4/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M3/M1/_1_  (.A(\V4/V3/V1/s1 [2]),
    .B(ground),
    .Z(\V4/V3/V1/A2/M3/s1 ));
 AND2_X1 \V4/V3/V1/A2/M3/M2/_0_  (.A1(\V4/V3/V1/A2/M3/s1 ),
    .A2(\V4/V3/V1/A2/c2 ),
    .ZN(\V4/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M3/M2/_1_  (.A(\V4/V3/V1/A2/M3/s1 ),
    .B(\V4/V3/V1/A2/c2 ),
    .Z(\V4/V3/V1/s2 [2]));
 OR2_X1 \V4/V3/V1/A2/M3/_0_  (.A1(\V4/V3/V1/A2/M3/c1 ),
    .A2(\V4/V3/V1/A2/M3/c2 ),
    .ZN(\V4/V3/V1/A2/c3 ));
 AND2_X1 \V4/V3/V1/A2/M4/M1/_0_  (.A1(\V4/V3/V1/s1 [3]),
    .A2(ground),
    .ZN(\V4/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M4/M1/_1_  (.A(\V4/V3/V1/s1 [3]),
    .B(ground),
    .Z(\V4/V3/V1/A2/M4/s1 ));
 AND2_X1 \V4/V3/V1/A2/M4/M2/_0_  (.A1(\V4/V3/V1/A2/M4/s1 ),
    .A2(\V4/V3/V1/A2/c3 ),
    .ZN(\V4/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M4/M2/_1_  (.A(\V4/V3/V1/A2/M4/s1 ),
    .B(\V4/V3/V1/A2/c3 ),
    .Z(\V4/V3/V1/s2 [3]));
 OR2_X1 \V4/V3/V1/A2/M4/_0_  (.A1(\V4/V3/V1/A2/M4/c1 ),
    .A2(\V4/V3/V1/A2/M4/c2 ),
    .ZN(\V4/V3/V1/c2 ));
 AND2_X1 \V4/V3/V1/A3/M1/M1/_0_  (.A1(\V4/V3/V1/v4 [0]),
    .A2(\V4/V3/V1/s2 [2]),
    .ZN(\V4/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M1/M1/_1_  (.A(\V4/V3/V1/v4 [0]),
    .B(\V4/V3/V1/s2 [2]),
    .Z(\V4/V3/V1/A3/M1/s1 ));
 AND2_X1 \V4/V3/V1/A3/M1/M2/_0_  (.A1(\V4/V3/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M1/M2/_1_  (.A(\V4/V3/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v1 [4]));
 OR2_X1 \V4/V3/V1/A3/M1/_0_  (.A1(\V4/V3/V1/A3/M1/c1 ),
    .A2(\V4/V3/V1/A3/M1/c2 ),
    .ZN(\V4/V3/V1/A3/c1 ));
 AND2_X1 \V4/V3/V1/A3/M2/M1/_0_  (.A1(\V4/V3/V1/v4 [1]),
    .A2(\V4/V3/V1/s2 [3]),
    .ZN(\V4/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M2/M1/_1_  (.A(\V4/V3/V1/v4 [1]),
    .B(\V4/V3/V1/s2 [3]),
    .Z(\V4/V3/V1/A3/M2/s1 ));
 AND2_X1 \V4/V3/V1/A3/M2/M2/_0_  (.A1(\V4/V3/V1/A3/M2/s1 ),
    .A2(\V4/V3/V1/A3/c1 ),
    .ZN(\V4/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M2/M2/_1_  (.A(\V4/V3/V1/A3/M2/s1 ),
    .B(\V4/V3/V1/A3/c1 ),
    .Z(\V4/V3/v1 [5]));
 OR2_X1 \V4/V3/V1/A3/M2/_0_  (.A1(\V4/V3/V1/A3/M2/c1 ),
    .A2(\V4/V3/V1/A3/M2/c2 ),
    .ZN(\V4/V3/V1/A3/c2 ));
 AND2_X1 \V4/V3/V1/A3/M3/M1/_0_  (.A1(\V4/V3/V1/v4 [2]),
    .A2(\V4/V3/V1/c3 ),
    .ZN(\V4/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M3/M1/_1_  (.A(\V4/V3/V1/v4 [2]),
    .B(\V4/V3/V1/c3 ),
    .Z(\V4/V3/V1/A3/M3/s1 ));
 AND2_X1 \V4/V3/V1/A3/M3/M2/_0_  (.A1(\V4/V3/V1/A3/M3/s1 ),
    .A2(\V4/V3/V1/A3/c2 ),
    .ZN(\V4/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M3/M2/_1_  (.A(\V4/V3/V1/A3/M3/s1 ),
    .B(\V4/V3/V1/A3/c2 ),
    .Z(\V4/V3/v1 [6]));
 OR2_X1 \V4/V3/V1/A3/M3/_0_  (.A1(\V4/V3/V1/A3/M3/c1 ),
    .A2(\V4/V3/V1/A3/M3/c2 ),
    .ZN(\V4/V3/V1/A3/c3 ));
 AND2_X1 \V4/V3/V1/A3/M4/M1/_0_  (.A1(\V4/V3/V1/v4 [3]),
    .A2(ground),
    .ZN(\V4/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M4/M1/_1_  (.A(\V4/V3/V1/v4 [3]),
    .B(ground),
    .Z(\V4/V3/V1/A3/M4/s1 ));
 AND2_X1 \V4/V3/V1/A3/M4/M2/_0_  (.A1(\V4/V3/V1/A3/M4/s1 ),
    .A2(\V4/V3/V1/A3/c3 ),
    .ZN(\V4/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M4/M2/_1_  (.A(\V4/V3/V1/A3/M4/s1 ),
    .B(\V4/V3/V1/A3/c3 ),
    .Z(\V4/V3/v1 [7]));
 OR2_X1 \V4/V3/V1/A3/M4/_0_  (.A1(\V4/V3/V1/A3/M4/c1 ),
    .A2(\V4/V3/V1/A3/M4/c2 ),
    .ZN(\V4/V3/V1/overflow ));
 AND2_X1 \V4/V3/V1/V1/HA1/_0_  (.A1(\V4/V3/V1/V1/w2 ),
    .A2(\V4/V3/V1/V1/w1 ),
    .ZN(\V4/V3/V1/V1/w4 ));
 XOR2_X2 \V4/V3/V1/V1/HA1/_1_  (.A(\V4/V3/V1/V1/w2 ),
    .B(\V4/V3/V1/V1/w1 ),
    .Z(\V4/v3 [1]));
 AND2_X1 \V4/V3/V1/V1/HA2/_0_  (.A1(\V4/V3/V1/V1/w4 ),
    .A2(\V4/V3/V1/V1/w3 ),
    .ZN(\V4/V3/V1/v1 [3]));
 XOR2_X2 \V4/V3/V1/V1/HA2/_1_  (.A(\V4/V3/V1/V1/w4 ),
    .B(\V4/V3/V1/V1/w3 ),
    .Z(\V4/V3/V1/v1 [2]));
 AND2_X1 \V4/V3/V1/V1/_0_  (.A1(A[16]),
    .A2(B[24]),
    .ZN(\V4/v3 [0]));
 AND2_X1 \V4/V3/V1/V1/_1_  (.A1(A[16]),
    .A2(B[25]),
    .ZN(\V4/V3/V1/V1/w1 ));
 AND2_X1 \V4/V3/V1/V1/_2_  (.A1(B[24]),
    .A2(A[17]),
    .ZN(\V4/V3/V1/V1/w2 ));
 AND2_X1 \V4/V3/V1/V1/_3_  (.A1(B[25]),
    .A2(A[17]),
    .ZN(\V4/V3/V1/V1/w3 ));
 AND2_X1 \V4/V3/V1/V2/HA1/_0_  (.A1(\V4/V3/V1/V2/w2 ),
    .A2(\V4/V3/V1/V2/w1 ),
    .ZN(\V4/V3/V1/V2/w4 ));
 XOR2_X2 \V4/V3/V1/V2/HA1/_1_  (.A(\V4/V3/V1/V2/w2 ),
    .B(\V4/V3/V1/V2/w1 ),
    .Z(\V4/V3/V1/v2 [1]));
 AND2_X1 \V4/V3/V1/V2/HA2/_0_  (.A1(\V4/V3/V1/V2/w4 ),
    .A2(\V4/V3/V1/V2/w3 ),
    .ZN(\V4/V3/V1/v2 [3]));
 XOR2_X2 \V4/V3/V1/V2/HA2/_1_  (.A(\V4/V3/V1/V2/w4 ),
    .B(\V4/V3/V1/V2/w3 ),
    .Z(\V4/V3/V1/v2 [2]));
 AND2_X1 \V4/V3/V1/V2/_0_  (.A1(A[18]),
    .A2(B[24]),
    .ZN(\V4/V3/V1/v2 [0]));
 AND2_X1 \V4/V3/V1/V2/_1_  (.A1(A[18]),
    .A2(B[25]),
    .ZN(\V4/V3/V1/V2/w1 ));
 AND2_X1 \V4/V3/V1/V2/_2_  (.A1(B[24]),
    .A2(A[19]),
    .ZN(\V4/V3/V1/V2/w2 ));
 AND2_X1 \V4/V3/V1/V2/_3_  (.A1(B[25]),
    .A2(A[19]),
    .ZN(\V4/V3/V1/V2/w3 ));
 AND2_X1 \V4/V3/V1/V3/HA1/_0_  (.A1(\V4/V3/V1/V3/w2 ),
    .A2(\V4/V3/V1/V3/w1 ),
    .ZN(\V4/V3/V1/V3/w4 ));
 XOR2_X2 \V4/V3/V1/V3/HA1/_1_  (.A(\V4/V3/V1/V3/w2 ),
    .B(\V4/V3/V1/V3/w1 ),
    .Z(\V4/V3/V1/v3 [1]));
 AND2_X1 \V4/V3/V1/V3/HA2/_0_  (.A1(\V4/V3/V1/V3/w4 ),
    .A2(\V4/V3/V1/V3/w3 ),
    .ZN(\V4/V3/V1/v3 [3]));
 XOR2_X2 \V4/V3/V1/V3/HA2/_1_  (.A(\V4/V3/V1/V3/w4 ),
    .B(\V4/V3/V1/V3/w3 ),
    .Z(\V4/V3/V1/v3 [2]));
 AND2_X1 \V4/V3/V1/V3/_0_  (.A1(A[16]),
    .A2(B[26]),
    .ZN(\V4/V3/V1/v3 [0]));
 AND2_X1 \V4/V3/V1/V3/_1_  (.A1(A[16]),
    .A2(B[27]),
    .ZN(\V4/V3/V1/V3/w1 ));
 AND2_X1 \V4/V3/V1/V3/_2_  (.A1(B[26]),
    .A2(A[17]),
    .ZN(\V4/V3/V1/V3/w2 ));
 AND2_X1 \V4/V3/V1/V3/_3_  (.A1(B[27]),
    .A2(A[17]),
    .ZN(\V4/V3/V1/V3/w3 ));
 AND2_X1 \V4/V3/V1/V4/HA1/_0_  (.A1(\V4/V3/V1/V4/w2 ),
    .A2(\V4/V3/V1/V4/w1 ),
    .ZN(\V4/V3/V1/V4/w4 ));
 XOR2_X2 \V4/V3/V1/V4/HA1/_1_  (.A(\V4/V3/V1/V4/w2 ),
    .B(\V4/V3/V1/V4/w1 ),
    .Z(\V4/V3/V1/v4 [1]));
 AND2_X1 \V4/V3/V1/V4/HA2/_0_  (.A1(\V4/V3/V1/V4/w4 ),
    .A2(\V4/V3/V1/V4/w3 ),
    .ZN(\V4/V3/V1/v4 [3]));
 XOR2_X2 \V4/V3/V1/V4/HA2/_1_  (.A(\V4/V3/V1/V4/w4 ),
    .B(\V4/V3/V1/V4/w3 ),
    .Z(\V4/V3/V1/v4 [2]));
 AND2_X1 \V4/V3/V1/V4/_0_  (.A1(A[18]),
    .A2(B[26]),
    .ZN(\V4/V3/V1/v4 [0]));
 AND2_X1 \V4/V3/V1/V4/_1_  (.A1(A[18]),
    .A2(B[27]),
    .ZN(\V4/V3/V1/V4/w1 ));
 AND2_X1 \V4/V3/V1/V4/_2_  (.A1(B[26]),
    .A2(A[19]),
    .ZN(\V4/V3/V1/V4/w2 ));
 AND2_X1 \V4/V3/V1/V4/_3_  (.A1(B[27]),
    .A2(A[19]),
    .ZN(\V4/V3/V1/V4/w3 ));
 OR2_X1 \V4/V3/V1/_0_  (.A1(\V4/V3/V1/c1 ),
    .A2(\V4/V3/V1/c2 ),
    .ZN(\V4/V3/V1/c3 ));
 AND2_X1 \V4/V3/V2/A1/M1/M1/_0_  (.A1(\V4/V3/V2/v2 [0]),
    .A2(\V4/V3/V2/v3 [0]),
    .ZN(\V4/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M1/M1/_1_  (.A(\V4/V3/V2/v2 [0]),
    .B(\V4/V3/V2/v3 [0]),
    .Z(\V4/V3/V2/A1/M1/s1 ));
 AND2_X1 \V4/V3/V2/A1/M1/M2/_0_  (.A1(\V4/V3/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M1/M2/_1_  (.A(\V4/V3/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/V2/s1 [0]));
 OR2_X1 \V4/V3/V2/A1/M1/_0_  (.A1(\V4/V3/V2/A1/M1/c1 ),
    .A2(\V4/V3/V2/A1/M1/c2 ),
    .ZN(\V4/V3/V2/A1/c1 ));
 AND2_X1 \V4/V3/V2/A1/M2/M1/_0_  (.A1(\V4/V3/V2/v2 [1]),
    .A2(\V4/V3/V2/v3 [1]),
    .ZN(\V4/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M2/M1/_1_  (.A(\V4/V3/V2/v2 [1]),
    .B(\V4/V3/V2/v3 [1]),
    .Z(\V4/V3/V2/A1/M2/s1 ));
 AND2_X1 \V4/V3/V2/A1/M2/M2/_0_  (.A1(\V4/V3/V2/A1/M2/s1 ),
    .A2(\V4/V3/V2/A1/c1 ),
    .ZN(\V4/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M2/M2/_1_  (.A(\V4/V3/V2/A1/M2/s1 ),
    .B(\V4/V3/V2/A1/c1 ),
    .Z(\V4/V3/V2/s1 [1]));
 OR2_X1 \V4/V3/V2/A1/M2/_0_  (.A1(\V4/V3/V2/A1/M2/c1 ),
    .A2(\V4/V3/V2/A1/M2/c2 ),
    .ZN(\V4/V3/V2/A1/c2 ));
 AND2_X1 \V4/V3/V2/A1/M3/M1/_0_  (.A1(\V4/V3/V2/v2 [2]),
    .A2(\V4/V3/V2/v3 [2]),
    .ZN(\V4/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M3/M1/_1_  (.A(\V4/V3/V2/v2 [2]),
    .B(\V4/V3/V2/v3 [2]),
    .Z(\V4/V3/V2/A1/M3/s1 ));
 AND2_X1 \V4/V3/V2/A1/M3/M2/_0_  (.A1(\V4/V3/V2/A1/M3/s1 ),
    .A2(\V4/V3/V2/A1/c2 ),
    .ZN(\V4/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M3/M2/_1_  (.A(\V4/V3/V2/A1/M3/s1 ),
    .B(\V4/V3/V2/A1/c2 ),
    .Z(\V4/V3/V2/s1 [2]));
 OR2_X1 \V4/V3/V2/A1/M3/_0_  (.A1(\V4/V3/V2/A1/M3/c1 ),
    .A2(\V4/V3/V2/A1/M3/c2 ),
    .ZN(\V4/V3/V2/A1/c3 ));
 AND2_X1 \V4/V3/V2/A1/M4/M1/_0_  (.A1(\V4/V3/V2/v2 [3]),
    .A2(\V4/V3/V2/v3 [3]),
    .ZN(\V4/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M4/M1/_1_  (.A(\V4/V3/V2/v2 [3]),
    .B(\V4/V3/V2/v3 [3]),
    .Z(\V4/V3/V2/A1/M4/s1 ));
 AND2_X1 \V4/V3/V2/A1/M4/M2/_0_  (.A1(\V4/V3/V2/A1/M4/s1 ),
    .A2(\V4/V3/V2/A1/c3 ),
    .ZN(\V4/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M4/M2/_1_  (.A(\V4/V3/V2/A1/M4/s1 ),
    .B(\V4/V3/V2/A1/c3 ),
    .Z(\V4/V3/V2/s1 [3]));
 OR2_X1 \V4/V3/V2/A1/M4/_0_  (.A1(\V4/V3/V2/A1/M4/c1 ),
    .A2(\V4/V3/V2/A1/M4/c2 ),
    .ZN(\V4/V3/V2/c1 ));
 AND2_X1 \V4/V3/V2/A2/M1/M1/_0_  (.A1(\V4/V3/V2/s1 [0]),
    .A2(\V4/V3/V2/v1 [2]),
    .ZN(\V4/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M1/M1/_1_  (.A(\V4/V3/V2/s1 [0]),
    .B(\V4/V3/V2/v1 [2]),
    .Z(\V4/V3/V2/A2/M1/s1 ));
 AND2_X1 \V4/V3/V2/A2/M1/M2/_0_  (.A1(\V4/V3/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M1/M2/_1_  (.A(\V4/V3/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v2 [2]));
 OR2_X1 \V4/V3/V2/A2/M1/_0_  (.A1(\V4/V3/V2/A2/M1/c1 ),
    .A2(\V4/V3/V2/A2/M1/c2 ),
    .ZN(\V4/V3/V2/A2/c1 ));
 AND2_X1 \V4/V3/V2/A2/M2/M1/_0_  (.A1(\V4/V3/V2/s1 [1]),
    .A2(\V4/V3/V2/v1 [3]),
    .ZN(\V4/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M2/M1/_1_  (.A(\V4/V3/V2/s1 [1]),
    .B(\V4/V3/V2/v1 [3]),
    .Z(\V4/V3/V2/A2/M2/s1 ));
 AND2_X1 \V4/V3/V2/A2/M2/M2/_0_  (.A1(\V4/V3/V2/A2/M2/s1 ),
    .A2(\V4/V3/V2/A2/c1 ),
    .ZN(\V4/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M2/M2/_1_  (.A(\V4/V3/V2/A2/M2/s1 ),
    .B(\V4/V3/V2/A2/c1 ),
    .Z(\V4/V3/v2 [3]));
 OR2_X1 \V4/V3/V2/A2/M2/_0_  (.A1(\V4/V3/V2/A2/M2/c1 ),
    .A2(\V4/V3/V2/A2/M2/c2 ),
    .ZN(\V4/V3/V2/A2/c2 ));
 AND2_X1 \V4/V3/V2/A2/M3/M1/_0_  (.A1(\V4/V3/V2/s1 [2]),
    .A2(ground),
    .ZN(\V4/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M3/M1/_1_  (.A(\V4/V3/V2/s1 [2]),
    .B(ground),
    .Z(\V4/V3/V2/A2/M3/s1 ));
 AND2_X1 \V4/V3/V2/A2/M3/M2/_0_  (.A1(\V4/V3/V2/A2/M3/s1 ),
    .A2(\V4/V3/V2/A2/c2 ),
    .ZN(\V4/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M3/M2/_1_  (.A(\V4/V3/V2/A2/M3/s1 ),
    .B(\V4/V3/V2/A2/c2 ),
    .Z(\V4/V3/V2/s2 [2]));
 OR2_X1 \V4/V3/V2/A2/M3/_0_  (.A1(\V4/V3/V2/A2/M3/c1 ),
    .A2(\V4/V3/V2/A2/M3/c2 ),
    .ZN(\V4/V3/V2/A2/c3 ));
 AND2_X1 \V4/V3/V2/A2/M4/M1/_0_  (.A1(\V4/V3/V2/s1 [3]),
    .A2(ground),
    .ZN(\V4/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M4/M1/_1_  (.A(\V4/V3/V2/s1 [3]),
    .B(ground),
    .Z(\V4/V3/V2/A2/M4/s1 ));
 AND2_X1 \V4/V3/V2/A2/M4/M2/_0_  (.A1(\V4/V3/V2/A2/M4/s1 ),
    .A2(\V4/V3/V2/A2/c3 ),
    .ZN(\V4/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M4/M2/_1_  (.A(\V4/V3/V2/A2/M4/s1 ),
    .B(\V4/V3/V2/A2/c3 ),
    .Z(\V4/V3/V2/s2 [3]));
 OR2_X1 \V4/V3/V2/A2/M4/_0_  (.A1(\V4/V3/V2/A2/M4/c1 ),
    .A2(\V4/V3/V2/A2/M4/c2 ),
    .ZN(\V4/V3/V2/c2 ));
 AND2_X1 \V4/V3/V2/A3/M1/M1/_0_  (.A1(\V4/V3/V2/v4 [0]),
    .A2(\V4/V3/V2/s2 [2]),
    .ZN(\V4/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M1/M1/_1_  (.A(\V4/V3/V2/v4 [0]),
    .B(\V4/V3/V2/s2 [2]),
    .Z(\V4/V3/V2/A3/M1/s1 ));
 AND2_X1 \V4/V3/V2/A3/M1/M2/_0_  (.A1(\V4/V3/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M1/M2/_1_  (.A(\V4/V3/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v2 [4]));
 OR2_X1 \V4/V3/V2/A3/M1/_0_  (.A1(\V4/V3/V2/A3/M1/c1 ),
    .A2(\V4/V3/V2/A3/M1/c2 ),
    .ZN(\V4/V3/V2/A3/c1 ));
 AND2_X1 \V4/V3/V2/A3/M2/M1/_0_  (.A1(\V4/V3/V2/v4 [1]),
    .A2(\V4/V3/V2/s2 [3]),
    .ZN(\V4/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M2/M1/_1_  (.A(\V4/V3/V2/v4 [1]),
    .B(\V4/V3/V2/s2 [3]),
    .Z(\V4/V3/V2/A3/M2/s1 ));
 AND2_X1 \V4/V3/V2/A3/M2/M2/_0_  (.A1(\V4/V3/V2/A3/M2/s1 ),
    .A2(\V4/V3/V2/A3/c1 ),
    .ZN(\V4/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M2/M2/_1_  (.A(\V4/V3/V2/A3/M2/s1 ),
    .B(\V4/V3/V2/A3/c1 ),
    .Z(\V4/V3/v2 [5]));
 OR2_X1 \V4/V3/V2/A3/M2/_0_  (.A1(\V4/V3/V2/A3/M2/c1 ),
    .A2(\V4/V3/V2/A3/M2/c2 ),
    .ZN(\V4/V3/V2/A3/c2 ));
 AND2_X1 \V4/V3/V2/A3/M3/M1/_0_  (.A1(\V4/V3/V2/v4 [2]),
    .A2(\V4/V3/V2/c3 ),
    .ZN(\V4/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M3/M1/_1_  (.A(\V4/V3/V2/v4 [2]),
    .B(\V4/V3/V2/c3 ),
    .Z(\V4/V3/V2/A3/M3/s1 ));
 AND2_X1 \V4/V3/V2/A3/M3/M2/_0_  (.A1(\V4/V3/V2/A3/M3/s1 ),
    .A2(\V4/V3/V2/A3/c2 ),
    .ZN(\V4/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M3/M2/_1_  (.A(\V4/V3/V2/A3/M3/s1 ),
    .B(\V4/V3/V2/A3/c2 ),
    .Z(\V4/V3/v2 [6]));
 OR2_X1 \V4/V3/V2/A3/M3/_0_  (.A1(\V4/V3/V2/A3/M3/c1 ),
    .A2(\V4/V3/V2/A3/M3/c2 ),
    .ZN(\V4/V3/V2/A3/c3 ));
 AND2_X1 \V4/V3/V2/A3/M4/M1/_0_  (.A1(\V4/V3/V2/v4 [3]),
    .A2(ground),
    .ZN(\V4/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M4/M1/_1_  (.A(\V4/V3/V2/v4 [3]),
    .B(ground),
    .Z(\V4/V3/V2/A3/M4/s1 ));
 AND2_X1 \V4/V3/V2/A3/M4/M2/_0_  (.A1(\V4/V3/V2/A3/M4/s1 ),
    .A2(\V4/V3/V2/A3/c3 ),
    .ZN(\V4/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M4/M2/_1_  (.A(\V4/V3/V2/A3/M4/s1 ),
    .B(\V4/V3/V2/A3/c3 ),
    .Z(\V4/V3/v2 [7]));
 OR2_X1 \V4/V3/V2/A3/M4/_0_  (.A1(\V4/V3/V2/A3/M4/c1 ),
    .A2(\V4/V3/V2/A3/M4/c2 ),
    .ZN(\V4/V3/V2/overflow ));
 AND2_X1 \V4/V3/V2/V1/HA1/_0_  (.A1(\V4/V3/V2/V1/w2 ),
    .A2(\V4/V3/V2/V1/w1 ),
    .ZN(\V4/V3/V2/V1/w4 ));
 XOR2_X2 \V4/V3/V2/V1/HA1/_1_  (.A(\V4/V3/V2/V1/w2 ),
    .B(\V4/V3/V2/V1/w1 ),
    .Z(\V4/V3/v2 [1]));
 AND2_X1 \V4/V3/V2/V1/HA2/_0_  (.A1(\V4/V3/V2/V1/w4 ),
    .A2(\V4/V3/V2/V1/w3 ),
    .ZN(\V4/V3/V2/v1 [3]));
 XOR2_X2 \V4/V3/V2/V1/HA2/_1_  (.A(\V4/V3/V2/V1/w4 ),
    .B(\V4/V3/V2/V1/w3 ),
    .Z(\V4/V3/V2/v1 [2]));
 AND2_X1 \V4/V3/V2/V1/_0_  (.A1(A[20]),
    .A2(B[24]),
    .ZN(\V4/V3/v2 [0]));
 AND2_X1 \V4/V3/V2/V1/_1_  (.A1(A[20]),
    .A2(B[25]),
    .ZN(\V4/V3/V2/V1/w1 ));
 AND2_X1 \V4/V3/V2/V1/_2_  (.A1(B[24]),
    .A2(A[21]),
    .ZN(\V4/V3/V2/V1/w2 ));
 AND2_X1 \V4/V3/V2/V1/_3_  (.A1(B[25]),
    .A2(A[21]),
    .ZN(\V4/V3/V2/V1/w3 ));
 AND2_X1 \V4/V3/V2/V2/HA1/_0_  (.A1(\V4/V3/V2/V2/w2 ),
    .A2(\V4/V3/V2/V2/w1 ),
    .ZN(\V4/V3/V2/V2/w4 ));
 XOR2_X2 \V4/V3/V2/V2/HA1/_1_  (.A(\V4/V3/V2/V2/w2 ),
    .B(\V4/V3/V2/V2/w1 ),
    .Z(\V4/V3/V2/v2 [1]));
 AND2_X1 \V4/V3/V2/V2/HA2/_0_  (.A1(\V4/V3/V2/V2/w4 ),
    .A2(\V4/V3/V2/V2/w3 ),
    .ZN(\V4/V3/V2/v2 [3]));
 XOR2_X2 \V4/V3/V2/V2/HA2/_1_  (.A(\V4/V3/V2/V2/w4 ),
    .B(\V4/V3/V2/V2/w3 ),
    .Z(\V4/V3/V2/v2 [2]));
 AND2_X1 \V4/V3/V2/V2/_0_  (.A1(A[22]),
    .A2(B[24]),
    .ZN(\V4/V3/V2/v2 [0]));
 AND2_X1 \V4/V3/V2/V2/_1_  (.A1(A[22]),
    .A2(B[25]),
    .ZN(\V4/V3/V2/V2/w1 ));
 AND2_X1 \V4/V3/V2/V2/_2_  (.A1(B[24]),
    .A2(A[23]),
    .ZN(\V4/V3/V2/V2/w2 ));
 AND2_X1 \V4/V3/V2/V2/_3_  (.A1(B[25]),
    .A2(A[23]),
    .ZN(\V4/V3/V2/V2/w3 ));
 AND2_X1 \V4/V3/V2/V3/HA1/_0_  (.A1(\V4/V3/V2/V3/w2 ),
    .A2(\V4/V3/V2/V3/w1 ),
    .ZN(\V4/V3/V2/V3/w4 ));
 XOR2_X2 \V4/V3/V2/V3/HA1/_1_  (.A(\V4/V3/V2/V3/w2 ),
    .B(\V4/V3/V2/V3/w1 ),
    .Z(\V4/V3/V2/v3 [1]));
 AND2_X1 \V4/V3/V2/V3/HA2/_0_  (.A1(\V4/V3/V2/V3/w4 ),
    .A2(\V4/V3/V2/V3/w3 ),
    .ZN(\V4/V3/V2/v3 [3]));
 XOR2_X2 \V4/V3/V2/V3/HA2/_1_  (.A(\V4/V3/V2/V3/w4 ),
    .B(\V4/V3/V2/V3/w3 ),
    .Z(\V4/V3/V2/v3 [2]));
 AND2_X1 \V4/V3/V2/V3/_0_  (.A1(A[20]),
    .A2(B[26]),
    .ZN(\V4/V3/V2/v3 [0]));
 AND2_X1 \V4/V3/V2/V3/_1_  (.A1(A[20]),
    .A2(B[27]),
    .ZN(\V4/V3/V2/V3/w1 ));
 AND2_X1 \V4/V3/V2/V3/_2_  (.A1(B[26]),
    .A2(A[21]),
    .ZN(\V4/V3/V2/V3/w2 ));
 AND2_X1 \V4/V3/V2/V3/_3_  (.A1(B[27]),
    .A2(A[21]),
    .ZN(\V4/V3/V2/V3/w3 ));
 AND2_X1 \V4/V3/V2/V4/HA1/_0_  (.A1(\V4/V3/V2/V4/w2 ),
    .A2(\V4/V3/V2/V4/w1 ),
    .ZN(\V4/V3/V2/V4/w4 ));
 XOR2_X2 \V4/V3/V2/V4/HA1/_1_  (.A(\V4/V3/V2/V4/w2 ),
    .B(\V4/V3/V2/V4/w1 ),
    .Z(\V4/V3/V2/v4 [1]));
 AND2_X1 \V4/V3/V2/V4/HA2/_0_  (.A1(\V4/V3/V2/V4/w4 ),
    .A2(\V4/V3/V2/V4/w3 ),
    .ZN(\V4/V3/V2/v4 [3]));
 XOR2_X2 \V4/V3/V2/V4/HA2/_1_  (.A(\V4/V3/V2/V4/w4 ),
    .B(\V4/V3/V2/V4/w3 ),
    .Z(\V4/V3/V2/v4 [2]));
 AND2_X1 \V4/V3/V2/V4/_0_  (.A1(A[22]),
    .A2(B[26]),
    .ZN(\V4/V3/V2/v4 [0]));
 AND2_X1 \V4/V3/V2/V4/_1_  (.A1(A[22]),
    .A2(B[27]),
    .ZN(\V4/V3/V2/V4/w1 ));
 AND2_X1 \V4/V3/V2/V4/_2_  (.A1(B[26]),
    .A2(A[23]),
    .ZN(\V4/V3/V2/V4/w2 ));
 AND2_X1 \V4/V3/V2/V4/_3_  (.A1(B[27]),
    .A2(A[23]),
    .ZN(\V4/V3/V2/V4/w3 ));
 OR2_X1 \V4/V3/V2/_0_  (.A1(\V4/V3/V2/c1 ),
    .A2(\V4/V3/V2/c2 ),
    .ZN(\V4/V3/V2/c3 ));
 AND2_X1 \V4/V3/V3/A1/M1/M1/_0_  (.A1(\V4/V3/V3/v2 [0]),
    .A2(\V4/V3/V3/v3 [0]),
    .ZN(\V4/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M1/M1/_1_  (.A(\V4/V3/V3/v2 [0]),
    .B(\V4/V3/V3/v3 [0]),
    .Z(\V4/V3/V3/A1/M1/s1 ));
 AND2_X1 \V4/V3/V3/A1/M1/M2/_0_  (.A1(\V4/V3/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M1/M2/_1_  (.A(\V4/V3/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/V3/s1 [0]));
 OR2_X1 \V4/V3/V3/A1/M1/_0_  (.A1(\V4/V3/V3/A1/M1/c1 ),
    .A2(\V4/V3/V3/A1/M1/c2 ),
    .ZN(\V4/V3/V3/A1/c1 ));
 AND2_X1 \V4/V3/V3/A1/M2/M1/_0_  (.A1(\V4/V3/V3/v2 [1]),
    .A2(\V4/V3/V3/v3 [1]),
    .ZN(\V4/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M2/M1/_1_  (.A(\V4/V3/V3/v2 [1]),
    .B(\V4/V3/V3/v3 [1]),
    .Z(\V4/V3/V3/A1/M2/s1 ));
 AND2_X1 \V4/V3/V3/A1/M2/M2/_0_  (.A1(\V4/V3/V3/A1/M2/s1 ),
    .A2(\V4/V3/V3/A1/c1 ),
    .ZN(\V4/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M2/M2/_1_  (.A(\V4/V3/V3/A1/M2/s1 ),
    .B(\V4/V3/V3/A1/c1 ),
    .Z(\V4/V3/V3/s1 [1]));
 OR2_X1 \V4/V3/V3/A1/M2/_0_  (.A1(\V4/V3/V3/A1/M2/c1 ),
    .A2(\V4/V3/V3/A1/M2/c2 ),
    .ZN(\V4/V3/V3/A1/c2 ));
 AND2_X1 \V4/V3/V3/A1/M3/M1/_0_  (.A1(\V4/V3/V3/v2 [2]),
    .A2(\V4/V3/V3/v3 [2]),
    .ZN(\V4/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M3/M1/_1_  (.A(\V4/V3/V3/v2 [2]),
    .B(\V4/V3/V3/v3 [2]),
    .Z(\V4/V3/V3/A1/M3/s1 ));
 AND2_X1 \V4/V3/V3/A1/M3/M2/_0_  (.A1(\V4/V3/V3/A1/M3/s1 ),
    .A2(\V4/V3/V3/A1/c2 ),
    .ZN(\V4/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M3/M2/_1_  (.A(\V4/V3/V3/A1/M3/s1 ),
    .B(\V4/V3/V3/A1/c2 ),
    .Z(\V4/V3/V3/s1 [2]));
 OR2_X1 \V4/V3/V3/A1/M3/_0_  (.A1(\V4/V3/V3/A1/M3/c1 ),
    .A2(\V4/V3/V3/A1/M3/c2 ),
    .ZN(\V4/V3/V3/A1/c3 ));
 AND2_X1 \V4/V3/V3/A1/M4/M1/_0_  (.A1(\V4/V3/V3/v2 [3]),
    .A2(\V4/V3/V3/v3 [3]),
    .ZN(\V4/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M4/M1/_1_  (.A(\V4/V3/V3/v2 [3]),
    .B(\V4/V3/V3/v3 [3]),
    .Z(\V4/V3/V3/A1/M4/s1 ));
 AND2_X1 \V4/V3/V3/A1/M4/M2/_0_  (.A1(\V4/V3/V3/A1/M4/s1 ),
    .A2(\V4/V3/V3/A1/c3 ),
    .ZN(\V4/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M4/M2/_1_  (.A(\V4/V3/V3/A1/M4/s1 ),
    .B(\V4/V3/V3/A1/c3 ),
    .Z(\V4/V3/V3/s1 [3]));
 OR2_X1 \V4/V3/V3/A1/M4/_0_  (.A1(\V4/V3/V3/A1/M4/c1 ),
    .A2(\V4/V3/V3/A1/M4/c2 ),
    .ZN(\V4/V3/V3/c1 ));
 AND2_X1 \V4/V3/V3/A2/M1/M1/_0_  (.A1(\V4/V3/V3/s1 [0]),
    .A2(\V4/V3/V3/v1 [2]),
    .ZN(\V4/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M1/M1/_1_  (.A(\V4/V3/V3/s1 [0]),
    .B(\V4/V3/V3/v1 [2]),
    .Z(\V4/V3/V3/A2/M1/s1 ));
 AND2_X1 \V4/V3/V3/A2/M1/M2/_0_  (.A1(\V4/V3/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M1/M2/_1_  (.A(\V4/V3/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v3 [2]));
 OR2_X1 \V4/V3/V3/A2/M1/_0_  (.A1(\V4/V3/V3/A2/M1/c1 ),
    .A2(\V4/V3/V3/A2/M1/c2 ),
    .ZN(\V4/V3/V3/A2/c1 ));
 AND2_X1 \V4/V3/V3/A2/M2/M1/_0_  (.A1(\V4/V3/V3/s1 [1]),
    .A2(\V4/V3/V3/v1 [3]),
    .ZN(\V4/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M2/M1/_1_  (.A(\V4/V3/V3/s1 [1]),
    .B(\V4/V3/V3/v1 [3]),
    .Z(\V4/V3/V3/A2/M2/s1 ));
 AND2_X1 \V4/V3/V3/A2/M2/M2/_0_  (.A1(\V4/V3/V3/A2/M2/s1 ),
    .A2(\V4/V3/V3/A2/c1 ),
    .ZN(\V4/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M2/M2/_1_  (.A(\V4/V3/V3/A2/M2/s1 ),
    .B(\V4/V3/V3/A2/c1 ),
    .Z(\V4/V3/v3 [3]));
 OR2_X1 \V4/V3/V3/A2/M2/_0_  (.A1(\V4/V3/V3/A2/M2/c1 ),
    .A2(\V4/V3/V3/A2/M2/c2 ),
    .ZN(\V4/V3/V3/A2/c2 ));
 AND2_X1 \V4/V3/V3/A2/M3/M1/_0_  (.A1(\V4/V3/V3/s1 [2]),
    .A2(ground),
    .ZN(\V4/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M3/M1/_1_  (.A(\V4/V3/V3/s1 [2]),
    .B(ground),
    .Z(\V4/V3/V3/A2/M3/s1 ));
 AND2_X1 \V4/V3/V3/A2/M3/M2/_0_  (.A1(\V4/V3/V3/A2/M3/s1 ),
    .A2(\V4/V3/V3/A2/c2 ),
    .ZN(\V4/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M3/M2/_1_  (.A(\V4/V3/V3/A2/M3/s1 ),
    .B(\V4/V3/V3/A2/c2 ),
    .Z(\V4/V3/V3/s2 [2]));
 OR2_X1 \V4/V3/V3/A2/M3/_0_  (.A1(\V4/V3/V3/A2/M3/c1 ),
    .A2(\V4/V3/V3/A2/M3/c2 ),
    .ZN(\V4/V3/V3/A2/c3 ));
 AND2_X1 \V4/V3/V3/A2/M4/M1/_0_  (.A1(\V4/V3/V3/s1 [3]),
    .A2(ground),
    .ZN(\V4/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M4/M1/_1_  (.A(\V4/V3/V3/s1 [3]),
    .B(ground),
    .Z(\V4/V3/V3/A2/M4/s1 ));
 AND2_X1 \V4/V3/V3/A2/M4/M2/_0_  (.A1(\V4/V3/V3/A2/M4/s1 ),
    .A2(\V4/V3/V3/A2/c3 ),
    .ZN(\V4/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M4/M2/_1_  (.A(\V4/V3/V3/A2/M4/s1 ),
    .B(\V4/V3/V3/A2/c3 ),
    .Z(\V4/V3/V3/s2 [3]));
 OR2_X1 \V4/V3/V3/A2/M4/_0_  (.A1(\V4/V3/V3/A2/M4/c1 ),
    .A2(\V4/V3/V3/A2/M4/c2 ),
    .ZN(\V4/V3/V3/c2 ));
 AND2_X1 \V4/V3/V3/A3/M1/M1/_0_  (.A1(\V4/V3/V3/v4 [0]),
    .A2(\V4/V3/V3/s2 [2]),
    .ZN(\V4/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M1/M1/_1_  (.A(\V4/V3/V3/v4 [0]),
    .B(\V4/V3/V3/s2 [2]),
    .Z(\V4/V3/V3/A3/M1/s1 ));
 AND2_X1 \V4/V3/V3/A3/M1/M2/_0_  (.A1(\V4/V3/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M1/M2/_1_  (.A(\V4/V3/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v3 [4]));
 OR2_X1 \V4/V3/V3/A3/M1/_0_  (.A1(\V4/V3/V3/A3/M1/c1 ),
    .A2(\V4/V3/V3/A3/M1/c2 ),
    .ZN(\V4/V3/V3/A3/c1 ));
 AND2_X1 \V4/V3/V3/A3/M2/M1/_0_  (.A1(\V4/V3/V3/v4 [1]),
    .A2(\V4/V3/V3/s2 [3]),
    .ZN(\V4/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M2/M1/_1_  (.A(\V4/V3/V3/v4 [1]),
    .B(\V4/V3/V3/s2 [3]),
    .Z(\V4/V3/V3/A3/M2/s1 ));
 AND2_X1 \V4/V3/V3/A3/M2/M2/_0_  (.A1(\V4/V3/V3/A3/M2/s1 ),
    .A2(\V4/V3/V3/A3/c1 ),
    .ZN(\V4/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M2/M2/_1_  (.A(\V4/V3/V3/A3/M2/s1 ),
    .B(\V4/V3/V3/A3/c1 ),
    .Z(\V4/V3/v3 [5]));
 OR2_X1 \V4/V3/V3/A3/M2/_0_  (.A1(\V4/V3/V3/A3/M2/c1 ),
    .A2(\V4/V3/V3/A3/M2/c2 ),
    .ZN(\V4/V3/V3/A3/c2 ));
 AND2_X1 \V4/V3/V3/A3/M3/M1/_0_  (.A1(\V4/V3/V3/v4 [2]),
    .A2(\V4/V3/V3/c3 ),
    .ZN(\V4/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M3/M1/_1_  (.A(\V4/V3/V3/v4 [2]),
    .B(\V4/V3/V3/c3 ),
    .Z(\V4/V3/V3/A3/M3/s1 ));
 AND2_X1 \V4/V3/V3/A3/M3/M2/_0_  (.A1(\V4/V3/V3/A3/M3/s1 ),
    .A2(\V4/V3/V3/A3/c2 ),
    .ZN(\V4/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M3/M2/_1_  (.A(\V4/V3/V3/A3/M3/s1 ),
    .B(\V4/V3/V3/A3/c2 ),
    .Z(\V4/V3/v3 [6]));
 OR2_X1 \V4/V3/V3/A3/M3/_0_  (.A1(\V4/V3/V3/A3/M3/c1 ),
    .A2(\V4/V3/V3/A3/M3/c2 ),
    .ZN(\V4/V3/V3/A3/c3 ));
 AND2_X1 \V4/V3/V3/A3/M4/M1/_0_  (.A1(\V4/V3/V3/v4 [3]),
    .A2(ground),
    .ZN(\V4/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M4/M1/_1_  (.A(\V4/V3/V3/v4 [3]),
    .B(ground),
    .Z(\V4/V3/V3/A3/M4/s1 ));
 AND2_X1 \V4/V3/V3/A3/M4/M2/_0_  (.A1(\V4/V3/V3/A3/M4/s1 ),
    .A2(\V4/V3/V3/A3/c3 ),
    .ZN(\V4/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M4/M2/_1_  (.A(\V4/V3/V3/A3/M4/s1 ),
    .B(\V4/V3/V3/A3/c3 ),
    .Z(\V4/V3/v3 [7]));
 OR2_X1 \V4/V3/V3/A3/M4/_0_  (.A1(\V4/V3/V3/A3/M4/c1 ),
    .A2(\V4/V3/V3/A3/M4/c2 ),
    .ZN(\V4/V3/V3/overflow ));
 AND2_X1 \V4/V3/V3/V1/HA1/_0_  (.A1(\V4/V3/V3/V1/w2 ),
    .A2(\V4/V3/V3/V1/w1 ),
    .ZN(\V4/V3/V3/V1/w4 ));
 XOR2_X2 \V4/V3/V3/V1/HA1/_1_  (.A(\V4/V3/V3/V1/w2 ),
    .B(\V4/V3/V3/V1/w1 ),
    .Z(\V4/V3/v3 [1]));
 AND2_X1 \V4/V3/V3/V1/HA2/_0_  (.A1(\V4/V3/V3/V1/w4 ),
    .A2(\V4/V3/V3/V1/w3 ),
    .ZN(\V4/V3/V3/v1 [3]));
 XOR2_X2 \V4/V3/V3/V1/HA2/_1_  (.A(\V4/V3/V3/V1/w4 ),
    .B(\V4/V3/V3/V1/w3 ),
    .Z(\V4/V3/V3/v1 [2]));
 AND2_X1 \V4/V3/V3/V1/_0_  (.A1(A[16]),
    .A2(B[28]),
    .ZN(\V4/V3/v3 [0]));
 AND2_X1 \V4/V3/V3/V1/_1_  (.A1(A[16]),
    .A2(B[29]),
    .ZN(\V4/V3/V3/V1/w1 ));
 AND2_X1 \V4/V3/V3/V1/_2_  (.A1(B[28]),
    .A2(A[17]),
    .ZN(\V4/V3/V3/V1/w2 ));
 AND2_X1 \V4/V3/V3/V1/_3_  (.A1(B[29]),
    .A2(A[17]),
    .ZN(\V4/V3/V3/V1/w3 ));
 AND2_X1 \V4/V3/V3/V2/HA1/_0_  (.A1(\V4/V3/V3/V2/w2 ),
    .A2(\V4/V3/V3/V2/w1 ),
    .ZN(\V4/V3/V3/V2/w4 ));
 XOR2_X2 \V4/V3/V3/V2/HA1/_1_  (.A(\V4/V3/V3/V2/w2 ),
    .B(\V4/V3/V3/V2/w1 ),
    .Z(\V4/V3/V3/v2 [1]));
 AND2_X1 \V4/V3/V3/V2/HA2/_0_  (.A1(\V4/V3/V3/V2/w4 ),
    .A2(\V4/V3/V3/V2/w3 ),
    .ZN(\V4/V3/V3/v2 [3]));
 XOR2_X2 \V4/V3/V3/V2/HA2/_1_  (.A(\V4/V3/V3/V2/w4 ),
    .B(\V4/V3/V3/V2/w3 ),
    .Z(\V4/V3/V3/v2 [2]));
 AND2_X1 \V4/V3/V3/V2/_0_  (.A1(A[18]),
    .A2(B[28]),
    .ZN(\V4/V3/V3/v2 [0]));
 AND2_X1 \V4/V3/V3/V2/_1_  (.A1(A[18]),
    .A2(B[29]),
    .ZN(\V4/V3/V3/V2/w1 ));
 AND2_X1 \V4/V3/V3/V2/_2_  (.A1(B[28]),
    .A2(A[19]),
    .ZN(\V4/V3/V3/V2/w2 ));
 AND2_X1 \V4/V3/V3/V2/_3_  (.A1(B[29]),
    .A2(A[19]),
    .ZN(\V4/V3/V3/V2/w3 ));
 AND2_X1 \V4/V3/V3/V3/HA1/_0_  (.A1(\V4/V3/V3/V3/w2 ),
    .A2(\V4/V3/V3/V3/w1 ),
    .ZN(\V4/V3/V3/V3/w4 ));
 XOR2_X2 \V4/V3/V3/V3/HA1/_1_  (.A(\V4/V3/V3/V3/w2 ),
    .B(\V4/V3/V3/V3/w1 ),
    .Z(\V4/V3/V3/v3 [1]));
 AND2_X1 \V4/V3/V3/V3/HA2/_0_  (.A1(\V4/V3/V3/V3/w4 ),
    .A2(\V4/V3/V3/V3/w3 ),
    .ZN(\V4/V3/V3/v3 [3]));
 XOR2_X2 \V4/V3/V3/V3/HA2/_1_  (.A(\V4/V3/V3/V3/w4 ),
    .B(\V4/V3/V3/V3/w3 ),
    .Z(\V4/V3/V3/v3 [2]));
 AND2_X1 \V4/V3/V3/V3/_0_  (.A1(A[16]),
    .A2(B[30]),
    .ZN(\V4/V3/V3/v3 [0]));
 AND2_X1 \V4/V3/V3/V3/_1_  (.A1(A[16]),
    .A2(B[31]),
    .ZN(\V4/V3/V3/V3/w1 ));
 AND2_X1 \V4/V3/V3/V3/_2_  (.A1(B[30]),
    .A2(A[17]),
    .ZN(\V4/V3/V3/V3/w2 ));
 AND2_X1 \V4/V3/V3/V3/_3_  (.A1(B[31]),
    .A2(A[17]),
    .ZN(\V4/V3/V3/V3/w3 ));
 AND2_X1 \V4/V3/V3/V4/HA1/_0_  (.A1(\V4/V3/V3/V4/w2 ),
    .A2(\V4/V3/V3/V4/w1 ),
    .ZN(\V4/V3/V3/V4/w4 ));
 XOR2_X2 \V4/V3/V3/V4/HA1/_1_  (.A(\V4/V3/V3/V4/w2 ),
    .B(\V4/V3/V3/V4/w1 ),
    .Z(\V4/V3/V3/v4 [1]));
 AND2_X1 \V4/V3/V3/V4/HA2/_0_  (.A1(\V4/V3/V3/V4/w4 ),
    .A2(\V4/V3/V3/V4/w3 ),
    .ZN(\V4/V3/V3/v4 [3]));
 XOR2_X2 \V4/V3/V3/V4/HA2/_1_  (.A(\V4/V3/V3/V4/w4 ),
    .B(\V4/V3/V3/V4/w3 ),
    .Z(\V4/V3/V3/v4 [2]));
 AND2_X1 \V4/V3/V3/V4/_0_  (.A1(A[18]),
    .A2(B[30]),
    .ZN(\V4/V3/V3/v4 [0]));
 AND2_X1 \V4/V3/V3/V4/_1_  (.A1(A[18]),
    .A2(B[31]),
    .ZN(\V4/V3/V3/V4/w1 ));
 AND2_X1 \V4/V3/V3/V4/_2_  (.A1(B[30]),
    .A2(A[19]),
    .ZN(\V4/V3/V3/V4/w2 ));
 AND2_X1 \V4/V3/V3/V4/_3_  (.A1(B[31]),
    .A2(A[19]),
    .ZN(\V4/V3/V3/V4/w3 ));
 OR2_X1 \V4/V3/V3/_0_  (.A1(\V4/V3/V3/c1 ),
    .A2(\V4/V3/V3/c2 ),
    .ZN(\V4/V3/V3/c3 ));
 AND2_X1 \V4/V3/V4/A1/M1/M1/_0_  (.A1(\V4/V3/V4/v2 [0]),
    .A2(\V4/V3/V4/v3 [0]),
    .ZN(\V4/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M1/M1/_1_  (.A(\V4/V3/V4/v2 [0]),
    .B(\V4/V3/V4/v3 [0]),
    .Z(\V4/V3/V4/A1/M1/s1 ));
 AND2_X1 \V4/V3/V4/A1/M1/M2/_0_  (.A1(\V4/V3/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M1/M2/_1_  (.A(\V4/V3/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/V4/s1 [0]));
 OR2_X1 \V4/V3/V4/A1/M1/_0_  (.A1(\V4/V3/V4/A1/M1/c1 ),
    .A2(\V4/V3/V4/A1/M1/c2 ),
    .ZN(\V4/V3/V4/A1/c1 ));
 AND2_X1 \V4/V3/V4/A1/M2/M1/_0_  (.A1(\V4/V3/V4/v2 [1]),
    .A2(\V4/V3/V4/v3 [1]),
    .ZN(\V4/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M2/M1/_1_  (.A(\V4/V3/V4/v2 [1]),
    .B(\V4/V3/V4/v3 [1]),
    .Z(\V4/V3/V4/A1/M2/s1 ));
 AND2_X1 \V4/V3/V4/A1/M2/M2/_0_  (.A1(\V4/V3/V4/A1/M2/s1 ),
    .A2(\V4/V3/V4/A1/c1 ),
    .ZN(\V4/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M2/M2/_1_  (.A(\V4/V3/V4/A1/M2/s1 ),
    .B(\V4/V3/V4/A1/c1 ),
    .Z(\V4/V3/V4/s1 [1]));
 OR2_X1 \V4/V3/V4/A1/M2/_0_  (.A1(\V4/V3/V4/A1/M2/c1 ),
    .A2(\V4/V3/V4/A1/M2/c2 ),
    .ZN(\V4/V3/V4/A1/c2 ));
 AND2_X1 \V4/V3/V4/A1/M3/M1/_0_  (.A1(\V4/V3/V4/v2 [2]),
    .A2(\V4/V3/V4/v3 [2]),
    .ZN(\V4/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M3/M1/_1_  (.A(\V4/V3/V4/v2 [2]),
    .B(\V4/V3/V4/v3 [2]),
    .Z(\V4/V3/V4/A1/M3/s1 ));
 AND2_X1 \V4/V3/V4/A1/M3/M2/_0_  (.A1(\V4/V3/V4/A1/M3/s1 ),
    .A2(\V4/V3/V4/A1/c2 ),
    .ZN(\V4/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M3/M2/_1_  (.A(\V4/V3/V4/A1/M3/s1 ),
    .B(\V4/V3/V4/A1/c2 ),
    .Z(\V4/V3/V4/s1 [2]));
 OR2_X1 \V4/V3/V4/A1/M3/_0_  (.A1(\V4/V3/V4/A1/M3/c1 ),
    .A2(\V4/V3/V4/A1/M3/c2 ),
    .ZN(\V4/V3/V4/A1/c3 ));
 AND2_X1 \V4/V3/V4/A1/M4/M1/_0_  (.A1(\V4/V3/V4/v2 [3]),
    .A2(\V4/V3/V4/v3 [3]),
    .ZN(\V4/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M4/M1/_1_  (.A(\V4/V3/V4/v2 [3]),
    .B(\V4/V3/V4/v3 [3]),
    .Z(\V4/V3/V4/A1/M4/s1 ));
 AND2_X1 \V4/V3/V4/A1/M4/M2/_0_  (.A1(\V4/V3/V4/A1/M4/s1 ),
    .A2(\V4/V3/V4/A1/c3 ),
    .ZN(\V4/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M4/M2/_1_  (.A(\V4/V3/V4/A1/M4/s1 ),
    .B(\V4/V3/V4/A1/c3 ),
    .Z(\V4/V3/V4/s1 [3]));
 OR2_X1 \V4/V3/V4/A1/M4/_0_  (.A1(\V4/V3/V4/A1/M4/c1 ),
    .A2(\V4/V3/V4/A1/M4/c2 ),
    .ZN(\V4/V3/V4/c1 ));
 AND2_X1 \V4/V3/V4/A2/M1/M1/_0_  (.A1(\V4/V3/V4/s1 [0]),
    .A2(\V4/V3/V4/v1 [2]),
    .ZN(\V4/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M1/M1/_1_  (.A(\V4/V3/V4/s1 [0]),
    .B(\V4/V3/V4/v1 [2]),
    .Z(\V4/V3/V4/A2/M1/s1 ));
 AND2_X1 \V4/V3/V4/A2/M1/M2/_0_  (.A1(\V4/V3/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M1/M2/_1_  (.A(\V4/V3/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v4 [2]));
 OR2_X1 \V4/V3/V4/A2/M1/_0_  (.A1(\V4/V3/V4/A2/M1/c1 ),
    .A2(\V4/V3/V4/A2/M1/c2 ),
    .ZN(\V4/V3/V4/A2/c1 ));
 AND2_X1 \V4/V3/V4/A2/M2/M1/_0_  (.A1(\V4/V3/V4/s1 [1]),
    .A2(\V4/V3/V4/v1 [3]),
    .ZN(\V4/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M2/M1/_1_  (.A(\V4/V3/V4/s1 [1]),
    .B(\V4/V3/V4/v1 [3]),
    .Z(\V4/V3/V4/A2/M2/s1 ));
 AND2_X1 \V4/V3/V4/A2/M2/M2/_0_  (.A1(\V4/V3/V4/A2/M2/s1 ),
    .A2(\V4/V3/V4/A2/c1 ),
    .ZN(\V4/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M2/M2/_1_  (.A(\V4/V3/V4/A2/M2/s1 ),
    .B(\V4/V3/V4/A2/c1 ),
    .Z(\V4/V3/v4 [3]));
 OR2_X1 \V4/V3/V4/A2/M2/_0_  (.A1(\V4/V3/V4/A2/M2/c1 ),
    .A2(\V4/V3/V4/A2/M2/c2 ),
    .ZN(\V4/V3/V4/A2/c2 ));
 AND2_X1 \V4/V3/V4/A2/M3/M1/_0_  (.A1(\V4/V3/V4/s1 [2]),
    .A2(ground),
    .ZN(\V4/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M3/M1/_1_  (.A(\V4/V3/V4/s1 [2]),
    .B(ground),
    .Z(\V4/V3/V4/A2/M3/s1 ));
 AND2_X1 \V4/V3/V4/A2/M3/M2/_0_  (.A1(\V4/V3/V4/A2/M3/s1 ),
    .A2(\V4/V3/V4/A2/c2 ),
    .ZN(\V4/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M3/M2/_1_  (.A(\V4/V3/V4/A2/M3/s1 ),
    .B(\V4/V3/V4/A2/c2 ),
    .Z(\V4/V3/V4/s2 [2]));
 OR2_X1 \V4/V3/V4/A2/M3/_0_  (.A1(\V4/V3/V4/A2/M3/c1 ),
    .A2(\V4/V3/V4/A2/M3/c2 ),
    .ZN(\V4/V3/V4/A2/c3 ));
 AND2_X1 \V4/V3/V4/A2/M4/M1/_0_  (.A1(\V4/V3/V4/s1 [3]),
    .A2(ground),
    .ZN(\V4/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M4/M1/_1_  (.A(\V4/V3/V4/s1 [3]),
    .B(ground),
    .Z(\V4/V3/V4/A2/M4/s1 ));
 AND2_X1 \V4/V3/V4/A2/M4/M2/_0_  (.A1(\V4/V3/V4/A2/M4/s1 ),
    .A2(\V4/V3/V4/A2/c3 ),
    .ZN(\V4/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M4/M2/_1_  (.A(\V4/V3/V4/A2/M4/s1 ),
    .B(\V4/V3/V4/A2/c3 ),
    .Z(\V4/V3/V4/s2 [3]));
 OR2_X1 \V4/V3/V4/A2/M4/_0_  (.A1(\V4/V3/V4/A2/M4/c1 ),
    .A2(\V4/V3/V4/A2/M4/c2 ),
    .ZN(\V4/V3/V4/c2 ));
 AND2_X1 \V4/V3/V4/A3/M1/M1/_0_  (.A1(\V4/V3/V4/v4 [0]),
    .A2(\V4/V3/V4/s2 [2]),
    .ZN(\V4/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M1/M1/_1_  (.A(\V4/V3/V4/v4 [0]),
    .B(\V4/V3/V4/s2 [2]),
    .Z(\V4/V3/V4/A3/M1/s1 ));
 AND2_X1 \V4/V3/V4/A3/M1/M2/_0_  (.A1(\V4/V3/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M1/M2/_1_  (.A(\V4/V3/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V3/v4 [4]));
 OR2_X1 \V4/V3/V4/A3/M1/_0_  (.A1(\V4/V3/V4/A3/M1/c1 ),
    .A2(\V4/V3/V4/A3/M1/c2 ),
    .ZN(\V4/V3/V4/A3/c1 ));
 AND2_X1 \V4/V3/V4/A3/M2/M1/_0_  (.A1(\V4/V3/V4/v4 [1]),
    .A2(\V4/V3/V4/s2 [3]),
    .ZN(\V4/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M2/M1/_1_  (.A(\V4/V3/V4/v4 [1]),
    .B(\V4/V3/V4/s2 [3]),
    .Z(\V4/V3/V4/A3/M2/s1 ));
 AND2_X1 \V4/V3/V4/A3/M2/M2/_0_  (.A1(\V4/V3/V4/A3/M2/s1 ),
    .A2(\V4/V3/V4/A3/c1 ),
    .ZN(\V4/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M2/M2/_1_  (.A(\V4/V3/V4/A3/M2/s1 ),
    .B(\V4/V3/V4/A3/c1 ),
    .Z(\V4/V3/v4 [5]));
 OR2_X1 \V4/V3/V4/A3/M2/_0_  (.A1(\V4/V3/V4/A3/M2/c1 ),
    .A2(\V4/V3/V4/A3/M2/c2 ),
    .ZN(\V4/V3/V4/A3/c2 ));
 AND2_X1 \V4/V3/V4/A3/M3/M1/_0_  (.A1(\V4/V3/V4/v4 [2]),
    .A2(\V4/V3/V4/c3 ),
    .ZN(\V4/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M3/M1/_1_  (.A(\V4/V3/V4/v4 [2]),
    .B(\V4/V3/V4/c3 ),
    .Z(\V4/V3/V4/A3/M3/s1 ));
 AND2_X1 \V4/V3/V4/A3/M3/M2/_0_  (.A1(\V4/V3/V4/A3/M3/s1 ),
    .A2(\V4/V3/V4/A3/c2 ),
    .ZN(\V4/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M3/M2/_1_  (.A(\V4/V3/V4/A3/M3/s1 ),
    .B(\V4/V3/V4/A3/c2 ),
    .Z(\V4/V3/v4 [6]));
 OR2_X1 \V4/V3/V4/A3/M3/_0_  (.A1(\V4/V3/V4/A3/M3/c1 ),
    .A2(\V4/V3/V4/A3/M3/c2 ),
    .ZN(\V4/V3/V4/A3/c3 ));
 AND2_X1 \V4/V3/V4/A3/M4/M1/_0_  (.A1(\V4/V3/V4/v4 [3]),
    .A2(ground),
    .ZN(\V4/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M4/M1/_1_  (.A(\V4/V3/V4/v4 [3]),
    .B(ground),
    .Z(\V4/V3/V4/A3/M4/s1 ));
 AND2_X1 \V4/V3/V4/A3/M4/M2/_0_  (.A1(\V4/V3/V4/A3/M4/s1 ),
    .A2(\V4/V3/V4/A3/c3 ),
    .ZN(\V4/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M4/M2/_1_  (.A(\V4/V3/V4/A3/M4/s1 ),
    .B(\V4/V3/V4/A3/c3 ),
    .Z(\V4/V3/v4 [7]));
 OR2_X1 \V4/V3/V4/A3/M4/_0_  (.A1(\V4/V3/V4/A3/M4/c1 ),
    .A2(\V4/V3/V4/A3/M4/c2 ),
    .ZN(\V4/V3/V4/overflow ));
 AND2_X1 \V4/V3/V4/V1/HA1/_0_  (.A1(\V4/V3/V4/V1/w2 ),
    .A2(\V4/V3/V4/V1/w1 ),
    .ZN(\V4/V3/V4/V1/w4 ));
 XOR2_X2 \V4/V3/V4/V1/HA1/_1_  (.A(\V4/V3/V4/V1/w2 ),
    .B(\V4/V3/V4/V1/w1 ),
    .Z(\V4/V3/v4 [1]));
 AND2_X1 \V4/V3/V4/V1/HA2/_0_  (.A1(\V4/V3/V4/V1/w4 ),
    .A2(\V4/V3/V4/V1/w3 ),
    .ZN(\V4/V3/V4/v1 [3]));
 XOR2_X2 \V4/V3/V4/V1/HA2/_1_  (.A(\V4/V3/V4/V1/w4 ),
    .B(\V4/V3/V4/V1/w3 ),
    .Z(\V4/V3/V4/v1 [2]));
 AND2_X1 \V4/V3/V4/V1/_0_  (.A1(A[20]),
    .A2(B[28]),
    .ZN(\V4/V3/v4 [0]));
 AND2_X1 \V4/V3/V4/V1/_1_  (.A1(A[20]),
    .A2(B[29]),
    .ZN(\V4/V3/V4/V1/w1 ));
 AND2_X1 \V4/V3/V4/V1/_2_  (.A1(B[28]),
    .A2(A[21]),
    .ZN(\V4/V3/V4/V1/w2 ));
 AND2_X1 \V4/V3/V4/V1/_3_  (.A1(B[29]),
    .A2(A[21]),
    .ZN(\V4/V3/V4/V1/w3 ));
 AND2_X1 \V4/V3/V4/V2/HA1/_0_  (.A1(\V4/V3/V4/V2/w2 ),
    .A2(\V4/V3/V4/V2/w1 ),
    .ZN(\V4/V3/V4/V2/w4 ));
 XOR2_X2 \V4/V3/V4/V2/HA1/_1_  (.A(\V4/V3/V4/V2/w2 ),
    .B(\V4/V3/V4/V2/w1 ),
    .Z(\V4/V3/V4/v2 [1]));
 AND2_X1 \V4/V3/V4/V2/HA2/_0_  (.A1(\V4/V3/V4/V2/w4 ),
    .A2(\V4/V3/V4/V2/w3 ),
    .ZN(\V4/V3/V4/v2 [3]));
 XOR2_X2 \V4/V3/V4/V2/HA2/_1_  (.A(\V4/V3/V4/V2/w4 ),
    .B(\V4/V3/V4/V2/w3 ),
    .Z(\V4/V3/V4/v2 [2]));
 AND2_X1 \V4/V3/V4/V2/_0_  (.A1(A[22]),
    .A2(B[28]),
    .ZN(\V4/V3/V4/v2 [0]));
 AND2_X1 \V4/V3/V4/V2/_1_  (.A1(A[22]),
    .A2(B[29]),
    .ZN(\V4/V3/V4/V2/w1 ));
 AND2_X1 \V4/V3/V4/V2/_2_  (.A1(B[28]),
    .A2(A[23]),
    .ZN(\V4/V3/V4/V2/w2 ));
 AND2_X1 \V4/V3/V4/V2/_3_  (.A1(B[29]),
    .A2(A[23]),
    .ZN(\V4/V3/V4/V2/w3 ));
 AND2_X1 \V4/V3/V4/V3/HA1/_0_  (.A1(\V4/V3/V4/V3/w2 ),
    .A2(\V4/V3/V4/V3/w1 ),
    .ZN(\V4/V3/V4/V3/w4 ));
 XOR2_X2 \V4/V3/V4/V3/HA1/_1_  (.A(\V4/V3/V4/V3/w2 ),
    .B(\V4/V3/V4/V3/w1 ),
    .Z(\V4/V3/V4/v3 [1]));
 AND2_X1 \V4/V3/V4/V3/HA2/_0_  (.A1(\V4/V3/V4/V3/w4 ),
    .A2(\V4/V3/V4/V3/w3 ),
    .ZN(\V4/V3/V4/v3 [3]));
 XOR2_X2 \V4/V3/V4/V3/HA2/_1_  (.A(\V4/V3/V4/V3/w4 ),
    .B(\V4/V3/V4/V3/w3 ),
    .Z(\V4/V3/V4/v3 [2]));
 AND2_X1 \V4/V3/V4/V3/_0_  (.A1(A[20]),
    .A2(B[30]),
    .ZN(\V4/V3/V4/v3 [0]));
 AND2_X1 \V4/V3/V4/V3/_1_  (.A1(A[20]),
    .A2(B[31]),
    .ZN(\V4/V3/V4/V3/w1 ));
 AND2_X1 \V4/V3/V4/V3/_2_  (.A1(B[30]),
    .A2(A[21]),
    .ZN(\V4/V3/V4/V3/w2 ));
 AND2_X1 \V4/V3/V4/V3/_3_  (.A1(B[31]),
    .A2(A[21]),
    .ZN(\V4/V3/V4/V3/w3 ));
 AND2_X1 \V4/V3/V4/V4/HA1/_0_  (.A1(\V4/V3/V4/V4/w2 ),
    .A2(\V4/V3/V4/V4/w1 ),
    .ZN(\V4/V3/V4/V4/w4 ));
 XOR2_X2 \V4/V3/V4/V4/HA1/_1_  (.A(\V4/V3/V4/V4/w2 ),
    .B(\V4/V3/V4/V4/w1 ),
    .Z(\V4/V3/V4/v4 [1]));
 AND2_X1 \V4/V3/V4/V4/HA2/_0_  (.A1(\V4/V3/V4/V4/w4 ),
    .A2(\V4/V3/V4/V4/w3 ),
    .ZN(\V4/V3/V4/v4 [3]));
 XOR2_X2 \V4/V3/V4/V4/HA2/_1_  (.A(\V4/V3/V4/V4/w4 ),
    .B(\V4/V3/V4/V4/w3 ),
    .Z(\V4/V3/V4/v4 [2]));
 AND2_X1 \V4/V3/V4/V4/_0_  (.A1(A[22]),
    .A2(B[30]),
    .ZN(\V4/V3/V4/v4 [0]));
 AND2_X1 \V4/V3/V4/V4/_1_  (.A1(A[22]),
    .A2(B[31]),
    .ZN(\V4/V3/V4/V4/w1 ));
 AND2_X1 \V4/V3/V4/V4/_2_  (.A1(B[30]),
    .A2(A[23]),
    .ZN(\V4/V3/V4/V4/w2 ));
 AND2_X1 \V4/V3/V4/V4/_3_  (.A1(B[31]),
    .A2(A[23]),
    .ZN(\V4/V3/V4/V4/w3 ));
 OR2_X1 \V4/V3/V4/_0_  (.A1(\V4/V3/V4/c1 ),
    .A2(\V4/V3/V4/c2 ),
    .ZN(\V4/V3/V4/c3 ));
 OR2_X1 \V4/V3/_0_  (.A1(\V4/V3/c1 ),
    .A2(\V4/V3/c2 ),
    .ZN(\V4/V3/c3 ));
 AND2_X1 \V4/V4/A1/A1/M1/M1/_0_  (.A1(\V4/V4/v2 [0]),
    .A2(\V4/V4/v3 [0]),
    .ZN(\V4/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M1/M1/_1_  (.A(\V4/V4/v2 [0]),
    .B(\V4/V4/v3 [0]),
    .Z(\V4/V4/A1/A1/M1/s1 ));
 AND2_X1 \V4/V4/A1/A1/M1/M2/_0_  (.A1(\V4/V4/A1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M1/M2/_1_  (.A(\V4/V4/A1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/s1 [0]));
 OR2_X1 \V4/V4/A1/A1/M1/_0_  (.A1(\V4/V4/A1/A1/M1/c1 ),
    .A2(\V4/V4/A1/A1/M1/c2 ),
    .ZN(\V4/V4/A1/A1/c1 ));
 AND2_X1 \V4/V4/A1/A1/M2/M1/_0_  (.A1(\V4/V4/v2 [1]),
    .A2(\V4/V4/v3 [1]),
    .ZN(\V4/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M2/M1/_1_  (.A(\V4/V4/v2 [1]),
    .B(\V4/V4/v3 [1]),
    .Z(\V4/V4/A1/A1/M2/s1 ));
 AND2_X1 \V4/V4/A1/A1/M2/M2/_0_  (.A1(\V4/V4/A1/A1/M2/s1 ),
    .A2(\V4/V4/A1/A1/c1 ),
    .ZN(\V4/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M2/M2/_1_  (.A(\V4/V4/A1/A1/M2/s1 ),
    .B(\V4/V4/A1/A1/c1 ),
    .Z(\V4/V4/s1 [1]));
 OR2_X1 \V4/V4/A1/A1/M2/_0_  (.A1(\V4/V4/A1/A1/M2/c1 ),
    .A2(\V4/V4/A1/A1/M2/c2 ),
    .ZN(\V4/V4/A1/A1/c2 ));
 AND2_X1 \V4/V4/A1/A1/M3/M1/_0_  (.A1(\V4/V4/v2 [2]),
    .A2(\V4/V4/v3 [2]),
    .ZN(\V4/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M3/M1/_1_  (.A(\V4/V4/v2 [2]),
    .B(\V4/V4/v3 [2]),
    .Z(\V4/V4/A1/A1/M3/s1 ));
 AND2_X1 \V4/V4/A1/A1/M3/M2/_0_  (.A1(\V4/V4/A1/A1/M3/s1 ),
    .A2(\V4/V4/A1/A1/c2 ),
    .ZN(\V4/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M3/M2/_1_  (.A(\V4/V4/A1/A1/M3/s1 ),
    .B(\V4/V4/A1/A1/c2 ),
    .Z(\V4/V4/s1 [2]));
 OR2_X1 \V4/V4/A1/A1/M3/_0_  (.A1(\V4/V4/A1/A1/M3/c1 ),
    .A2(\V4/V4/A1/A1/M3/c2 ),
    .ZN(\V4/V4/A1/A1/c3 ));
 AND2_X1 \V4/V4/A1/A1/M4/M1/_0_  (.A1(\V4/V4/v2 [3]),
    .A2(\V4/V4/v3 [3]),
    .ZN(\V4/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M4/M1/_1_  (.A(\V4/V4/v2 [3]),
    .B(\V4/V4/v3 [3]),
    .Z(\V4/V4/A1/A1/M4/s1 ));
 AND2_X1 \V4/V4/A1/A1/M4/M2/_0_  (.A1(\V4/V4/A1/A1/M4/s1 ),
    .A2(\V4/V4/A1/A1/c3 ),
    .ZN(\V4/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M4/M2/_1_  (.A(\V4/V4/A1/A1/M4/s1 ),
    .B(\V4/V4/A1/A1/c3 ),
    .Z(\V4/V4/s1 [3]));
 OR2_X1 \V4/V4/A1/A1/M4/_0_  (.A1(\V4/V4/A1/A1/M4/c1 ),
    .A2(\V4/V4/A1/A1/M4/c2 ),
    .ZN(\V4/V4/A1/c1 ));
 AND2_X1 \V4/V4/A1/A2/M1/M1/_0_  (.A1(\V4/V4/v2 [4]),
    .A2(\V4/V4/v3 [4]),
    .ZN(\V4/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M1/M1/_1_  (.A(\V4/V4/v2 [4]),
    .B(\V4/V4/v3 [4]),
    .Z(\V4/V4/A1/A2/M1/s1 ));
 AND2_X1 \V4/V4/A1/A2/M1/M2/_0_  (.A1(\V4/V4/A1/A2/M1/s1 ),
    .A2(\V4/V4/A1/c1 ),
    .ZN(\V4/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M1/M2/_1_  (.A(\V4/V4/A1/A2/M1/s1 ),
    .B(\V4/V4/A1/c1 ),
    .Z(\V4/V4/s1 [4]));
 OR2_X1 \V4/V4/A1/A2/M1/_0_  (.A1(\V4/V4/A1/A2/M1/c1 ),
    .A2(\V4/V4/A1/A2/M1/c2 ),
    .ZN(\V4/V4/A1/A2/c1 ));
 AND2_X1 \V4/V4/A1/A2/M2/M1/_0_  (.A1(\V4/V4/v2 [5]),
    .A2(\V4/V4/v3 [5]),
    .ZN(\V4/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M2/M1/_1_  (.A(\V4/V4/v2 [5]),
    .B(\V4/V4/v3 [5]),
    .Z(\V4/V4/A1/A2/M2/s1 ));
 AND2_X1 \V4/V4/A1/A2/M2/M2/_0_  (.A1(\V4/V4/A1/A2/M2/s1 ),
    .A2(\V4/V4/A1/A2/c1 ),
    .ZN(\V4/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M2/M2/_1_  (.A(\V4/V4/A1/A2/M2/s1 ),
    .B(\V4/V4/A1/A2/c1 ),
    .Z(\V4/V4/s1 [5]));
 OR2_X1 \V4/V4/A1/A2/M2/_0_  (.A1(\V4/V4/A1/A2/M2/c1 ),
    .A2(\V4/V4/A1/A2/M2/c2 ),
    .ZN(\V4/V4/A1/A2/c2 ));
 AND2_X1 \V4/V4/A1/A2/M3/M1/_0_  (.A1(\V4/V4/v2 [6]),
    .A2(\V4/V4/v3 [6]),
    .ZN(\V4/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M3/M1/_1_  (.A(\V4/V4/v2 [6]),
    .B(\V4/V4/v3 [6]),
    .Z(\V4/V4/A1/A2/M3/s1 ));
 AND2_X1 \V4/V4/A1/A2/M3/M2/_0_  (.A1(\V4/V4/A1/A2/M3/s1 ),
    .A2(\V4/V4/A1/A2/c2 ),
    .ZN(\V4/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M3/M2/_1_  (.A(\V4/V4/A1/A2/M3/s1 ),
    .B(\V4/V4/A1/A2/c2 ),
    .Z(\V4/V4/s1 [6]));
 OR2_X1 \V4/V4/A1/A2/M3/_0_  (.A1(\V4/V4/A1/A2/M3/c1 ),
    .A2(\V4/V4/A1/A2/M3/c2 ),
    .ZN(\V4/V4/A1/A2/c3 ));
 AND2_X1 \V4/V4/A1/A2/M4/M1/_0_  (.A1(\V4/V4/v2 [7]),
    .A2(\V4/V4/v3 [7]),
    .ZN(\V4/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M4/M1/_1_  (.A(\V4/V4/v2 [7]),
    .B(\V4/V4/v3 [7]),
    .Z(\V4/V4/A1/A2/M4/s1 ));
 AND2_X1 \V4/V4/A1/A2/M4/M2/_0_  (.A1(\V4/V4/A1/A2/M4/s1 ),
    .A2(\V4/V4/A1/A2/c3 ),
    .ZN(\V4/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M4/M2/_1_  (.A(\V4/V4/A1/A2/M4/s1 ),
    .B(\V4/V4/A1/A2/c3 ),
    .Z(\V4/V4/s1 [7]));
 OR2_X1 \V4/V4/A1/A2/M4/_0_  (.A1(\V4/V4/A1/A2/M4/c1 ),
    .A2(\V4/V4/A1/A2/M4/c2 ),
    .ZN(\V4/V4/c1 ));
 AND2_X1 \V4/V4/A2/A1/M1/M1/_0_  (.A1(\V4/V4/s1 [0]),
    .A2(\V4/V4/v1 [4]),
    .ZN(\V4/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M1/M1/_1_  (.A(\V4/V4/s1 [0]),
    .B(\V4/V4/v1 [4]),
    .Z(\V4/V4/A2/A1/M1/s1 ));
 AND2_X1 \V4/V4/A2/A1/M1/M2/_0_  (.A1(\V4/V4/A2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M1/M2/_1_  (.A(\V4/V4/A2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v4 [4]));
 OR2_X1 \V4/V4/A2/A1/M1/_0_  (.A1(\V4/V4/A2/A1/M1/c1 ),
    .A2(\V4/V4/A2/A1/M1/c2 ),
    .ZN(\V4/V4/A2/A1/c1 ));
 AND2_X1 \V4/V4/A2/A1/M2/M1/_0_  (.A1(\V4/V4/s1 [1]),
    .A2(\V4/V4/v1 [5]),
    .ZN(\V4/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M2/M1/_1_  (.A(\V4/V4/s1 [1]),
    .B(\V4/V4/v1 [5]),
    .Z(\V4/V4/A2/A1/M2/s1 ));
 AND2_X1 \V4/V4/A2/A1/M2/M2/_0_  (.A1(\V4/V4/A2/A1/M2/s1 ),
    .A2(\V4/V4/A2/A1/c1 ),
    .ZN(\V4/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M2/M2/_1_  (.A(\V4/V4/A2/A1/M2/s1 ),
    .B(\V4/V4/A2/A1/c1 ),
    .Z(\V4/v4 [5]));
 OR2_X1 \V4/V4/A2/A1/M2/_0_  (.A1(\V4/V4/A2/A1/M2/c1 ),
    .A2(\V4/V4/A2/A1/M2/c2 ),
    .ZN(\V4/V4/A2/A1/c2 ));
 AND2_X1 \V4/V4/A2/A1/M3/M1/_0_  (.A1(\V4/V4/s1 [2]),
    .A2(\V4/V4/v1 [6]),
    .ZN(\V4/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M3/M1/_1_  (.A(\V4/V4/s1 [2]),
    .B(\V4/V4/v1 [6]),
    .Z(\V4/V4/A2/A1/M3/s1 ));
 AND2_X1 \V4/V4/A2/A1/M3/M2/_0_  (.A1(\V4/V4/A2/A1/M3/s1 ),
    .A2(\V4/V4/A2/A1/c2 ),
    .ZN(\V4/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M3/M2/_1_  (.A(\V4/V4/A2/A1/M3/s1 ),
    .B(\V4/V4/A2/A1/c2 ),
    .Z(\V4/v4 [6]));
 OR2_X1 \V4/V4/A2/A1/M3/_0_  (.A1(\V4/V4/A2/A1/M3/c1 ),
    .A2(\V4/V4/A2/A1/M3/c2 ),
    .ZN(\V4/V4/A2/A1/c3 ));
 AND2_X1 \V4/V4/A2/A1/M4/M1/_0_  (.A1(\V4/V4/s1 [3]),
    .A2(\V4/V4/v1 [7]),
    .ZN(\V4/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M4/M1/_1_  (.A(\V4/V4/s1 [3]),
    .B(\V4/V4/v1 [7]),
    .Z(\V4/V4/A2/A1/M4/s1 ));
 AND2_X1 \V4/V4/A2/A1/M4/M2/_0_  (.A1(\V4/V4/A2/A1/M4/s1 ),
    .A2(\V4/V4/A2/A1/c3 ),
    .ZN(\V4/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M4/M2/_1_  (.A(\V4/V4/A2/A1/M4/s1 ),
    .B(\V4/V4/A2/A1/c3 ),
    .Z(\V4/v4 [7]));
 OR2_X1 \V4/V4/A2/A1/M4/_0_  (.A1(\V4/V4/A2/A1/M4/c1 ),
    .A2(\V4/V4/A2/A1/M4/c2 ),
    .ZN(\V4/V4/A2/c1 ));
 AND2_X1 \V4/V4/A2/A2/M1/M1/_0_  (.A1(\V4/V4/s1 [4]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M1/M1/_1_  (.A(\V4/V4/s1 [4]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M1/s1 ));
 AND2_X1 \V4/V4/A2/A2/M1/M2/_0_  (.A1(\V4/V4/A2/A2/M1/s1 ),
    .A2(\V4/V4/A2/c1 ),
    .ZN(\V4/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M1/M2/_1_  (.A(\V4/V4/A2/A2/M1/s1 ),
    .B(\V4/V4/A2/c1 ),
    .Z(\V4/V4/s2 [4]));
 OR2_X1 \V4/V4/A2/A2/M1/_0_  (.A1(\V4/V4/A2/A2/M1/c1 ),
    .A2(\V4/V4/A2/A2/M1/c2 ),
    .ZN(\V4/V4/A2/A2/c1 ));
 AND2_X1 \V4/V4/A2/A2/M2/M1/_0_  (.A1(\V4/V4/s1 [5]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M2/M1/_1_  (.A(\V4/V4/s1 [5]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M2/s1 ));
 AND2_X1 \V4/V4/A2/A2/M2/M2/_0_  (.A1(\V4/V4/A2/A2/M2/s1 ),
    .A2(\V4/V4/A2/A2/c1 ),
    .ZN(\V4/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M2/M2/_1_  (.A(\V4/V4/A2/A2/M2/s1 ),
    .B(\V4/V4/A2/A2/c1 ),
    .Z(\V4/V4/s2 [5]));
 OR2_X1 \V4/V4/A2/A2/M2/_0_  (.A1(\V4/V4/A2/A2/M2/c1 ),
    .A2(\V4/V4/A2/A2/M2/c2 ),
    .ZN(\V4/V4/A2/A2/c2 ));
 AND2_X1 \V4/V4/A2/A2/M3/M1/_0_  (.A1(\V4/V4/s1 [6]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M3/M1/_1_  (.A(\V4/V4/s1 [6]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M3/s1 ));
 AND2_X1 \V4/V4/A2/A2/M3/M2/_0_  (.A1(\V4/V4/A2/A2/M3/s1 ),
    .A2(\V4/V4/A2/A2/c2 ),
    .ZN(\V4/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M3/M2/_1_  (.A(\V4/V4/A2/A2/M3/s1 ),
    .B(\V4/V4/A2/A2/c2 ),
    .Z(\V4/V4/s2 [6]));
 OR2_X1 \V4/V4/A2/A2/M3/_0_  (.A1(\V4/V4/A2/A2/M3/c1 ),
    .A2(\V4/V4/A2/A2/M3/c2 ),
    .ZN(\V4/V4/A2/A2/c3 ));
 AND2_X1 \V4/V4/A2/A2/M4/M1/_0_  (.A1(\V4/V4/s1 [7]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M4/M1/_1_  (.A(\V4/V4/s1 [7]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M4/s1 ));
 AND2_X1 \V4/V4/A2/A2/M4/M2/_0_  (.A1(\V4/V4/A2/A2/M4/s1 ),
    .A2(\V4/V4/A2/A2/c3 ),
    .ZN(\V4/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M4/M2/_1_  (.A(\V4/V4/A2/A2/M4/s1 ),
    .B(\V4/V4/A2/A2/c3 ),
    .Z(\V4/V4/s2 [7]));
 OR2_X1 \V4/V4/A2/A2/M4/_0_  (.A1(\V4/V4/A2/A2/M4/c1 ),
    .A2(\V4/V4/A2/A2/M4/c2 ),
    .ZN(\V4/V4/c2 ));
 AND2_X1 \V4/V4/A3/A1/M1/M1/_0_  (.A1(\V4/V4/v4 [0]),
    .A2(\V4/V4/s2 [4]),
    .ZN(\V4/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M1/M1/_1_  (.A(\V4/V4/v4 [0]),
    .B(\V4/V4/s2 [4]),
    .Z(\V4/V4/A3/A1/M1/s1 ));
 AND2_X1 \V4/V4/A3/A1/M1/M2/_0_  (.A1(\V4/V4/A3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M1/M2/_1_  (.A(\V4/V4/A3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/v4 [8]));
 OR2_X1 \V4/V4/A3/A1/M1/_0_  (.A1(\V4/V4/A3/A1/M1/c1 ),
    .A2(\V4/V4/A3/A1/M1/c2 ),
    .ZN(\V4/V4/A3/A1/c1 ));
 AND2_X1 \V4/V4/A3/A1/M2/M1/_0_  (.A1(\V4/V4/v4 [1]),
    .A2(\V4/V4/s2 [5]),
    .ZN(\V4/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M2/M1/_1_  (.A(\V4/V4/v4 [1]),
    .B(\V4/V4/s2 [5]),
    .Z(\V4/V4/A3/A1/M2/s1 ));
 AND2_X1 \V4/V4/A3/A1/M2/M2/_0_  (.A1(\V4/V4/A3/A1/M2/s1 ),
    .A2(\V4/V4/A3/A1/c1 ),
    .ZN(\V4/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M2/M2/_1_  (.A(\V4/V4/A3/A1/M2/s1 ),
    .B(\V4/V4/A3/A1/c1 ),
    .Z(\V4/v4 [9]));
 OR2_X1 \V4/V4/A3/A1/M2/_0_  (.A1(\V4/V4/A3/A1/M2/c1 ),
    .A2(\V4/V4/A3/A1/M2/c2 ),
    .ZN(\V4/V4/A3/A1/c2 ));
 AND2_X1 \V4/V4/A3/A1/M3/M1/_0_  (.A1(\V4/V4/v4 [2]),
    .A2(\V4/V4/s2 [6]),
    .ZN(\V4/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M3/M1/_1_  (.A(\V4/V4/v4 [2]),
    .B(\V4/V4/s2 [6]),
    .Z(\V4/V4/A3/A1/M3/s1 ));
 AND2_X1 \V4/V4/A3/A1/M3/M2/_0_  (.A1(\V4/V4/A3/A1/M3/s1 ),
    .A2(\V4/V4/A3/A1/c2 ),
    .ZN(\V4/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M3/M2/_1_  (.A(\V4/V4/A3/A1/M3/s1 ),
    .B(\V4/V4/A3/A1/c2 ),
    .Z(\V4/v4 [10]));
 OR2_X1 \V4/V4/A3/A1/M3/_0_  (.A1(\V4/V4/A3/A1/M3/c1 ),
    .A2(\V4/V4/A3/A1/M3/c2 ),
    .ZN(\V4/V4/A3/A1/c3 ));
 AND2_X1 \V4/V4/A3/A1/M4/M1/_0_  (.A1(\V4/V4/v4 [3]),
    .A2(\V4/V4/s2 [7]),
    .ZN(\V4/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M4/M1/_1_  (.A(\V4/V4/v4 [3]),
    .B(\V4/V4/s2 [7]),
    .Z(\V4/V4/A3/A1/M4/s1 ));
 AND2_X1 \V4/V4/A3/A1/M4/M2/_0_  (.A1(\V4/V4/A3/A1/M4/s1 ),
    .A2(\V4/V4/A3/A1/c3 ),
    .ZN(\V4/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M4/M2/_1_  (.A(\V4/V4/A3/A1/M4/s1 ),
    .B(\V4/V4/A3/A1/c3 ),
    .Z(\V4/v4 [11]));
 OR2_X1 \V4/V4/A3/A1/M4/_0_  (.A1(\V4/V4/A3/A1/M4/c1 ),
    .A2(\V4/V4/A3/A1/M4/c2 ),
    .ZN(\V4/V4/A3/c1 ));
 AND2_X1 \V4/V4/A3/A2/M1/M1/_0_  (.A1(\V4/V4/v4 [4]),
    .A2(\V4/V4/c3 ),
    .ZN(\V4/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M1/M1/_1_  (.A(\V4/V4/v4 [4]),
    .B(\V4/V4/c3 ),
    .Z(\V4/V4/A3/A2/M1/s1 ));
 AND2_X1 \V4/V4/A3/A2/M1/M2/_0_  (.A1(\V4/V4/A3/A2/M1/s1 ),
    .A2(\V4/V4/A3/c1 ),
    .ZN(\V4/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M1/M2/_1_  (.A(\V4/V4/A3/A2/M1/s1 ),
    .B(\V4/V4/A3/c1 ),
    .Z(\V4/v4 [12]));
 OR2_X1 \V4/V4/A3/A2/M1/_0_  (.A1(\V4/V4/A3/A2/M1/c1 ),
    .A2(\V4/V4/A3/A2/M1/c2 ),
    .ZN(\V4/V4/A3/A2/c1 ));
 AND2_X1 \V4/V4/A3/A2/M2/M1/_0_  (.A1(\V4/V4/v4 [5]),
    .A2(ground),
    .ZN(\V4/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M2/M1/_1_  (.A(\V4/V4/v4 [5]),
    .B(ground),
    .Z(\V4/V4/A3/A2/M2/s1 ));
 AND2_X1 \V4/V4/A3/A2/M2/M2/_0_  (.A1(\V4/V4/A3/A2/M2/s1 ),
    .A2(\V4/V4/A3/A2/c1 ),
    .ZN(\V4/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M2/M2/_1_  (.A(\V4/V4/A3/A2/M2/s1 ),
    .B(\V4/V4/A3/A2/c1 ),
    .Z(\V4/v4 [13]));
 OR2_X1 \V4/V4/A3/A2/M2/_0_  (.A1(\V4/V4/A3/A2/M2/c1 ),
    .A2(\V4/V4/A3/A2/M2/c2 ),
    .ZN(\V4/V4/A3/A2/c2 ));
 AND2_X1 \V4/V4/A3/A2/M3/M1/_0_  (.A1(\V4/V4/v4 [6]),
    .A2(ground),
    .ZN(\V4/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M3/M1/_1_  (.A(\V4/V4/v4 [6]),
    .B(ground),
    .Z(\V4/V4/A3/A2/M3/s1 ));
 AND2_X1 \V4/V4/A3/A2/M3/M2/_0_  (.A1(\V4/V4/A3/A2/M3/s1 ),
    .A2(\V4/V4/A3/A2/c2 ),
    .ZN(\V4/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M3/M2/_1_  (.A(\V4/V4/A3/A2/M3/s1 ),
    .B(\V4/V4/A3/A2/c2 ),
    .Z(\V4/v4 [14]));
 OR2_X1 \V4/V4/A3/A2/M3/_0_  (.A1(\V4/V4/A3/A2/M3/c1 ),
    .A2(\V4/V4/A3/A2/M3/c2 ),
    .ZN(\V4/V4/A3/A2/c3 ));
 AND2_X1 \V4/V4/A3/A2/M4/M1/_0_  (.A1(\V4/V4/v4 [7]),
    .A2(ground),
    .ZN(\V4/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M4/M1/_1_  (.A(\V4/V4/v4 [7]),
    .B(ground),
    .Z(\V4/V4/A3/A2/M4/s1 ));
 AND2_X1 \V4/V4/A3/A2/M4/M2/_0_  (.A1(\V4/V4/A3/A2/M4/s1 ),
    .A2(\V4/V4/A3/A2/c3 ),
    .ZN(\V4/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M4/M2/_1_  (.A(\V4/V4/A3/A2/M4/s1 ),
    .B(\V4/V4/A3/A2/c3 ),
    .Z(\V4/v4 [15]));
 OR2_X1 \V4/V4/A3/A2/M4/_0_  (.A1(\V4/V4/A3/A2/M4/c1 ),
    .A2(\V4/V4/A3/A2/M4/c2 ),
    .ZN(\V4/V4/overflow ));
 AND2_X1 \V4/V4/V1/A1/M1/M1/_0_  (.A1(\V4/V4/V1/v2 [0]),
    .A2(\V4/V4/V1/v3 [0]),
    .ZN(\V4/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M1/M1/_1_  (.A(\V4/V4/V1/v2 [0]),
    .B(\V4/V4/V1/v3 [0]),
    .Z(\V4/V4/V1/A1/M1/s1 ));
 AND2_X1 \V4/V4/V1/A1/M1/M2/_0_  (.A1(\V4/V4/V1/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M1/M2/_1_  (.A(\V4/V4/V1/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/V1/s1 [0]));
 OR2_X1 \V4/V4/V1/A1/M1/_0_  (.A1(\V4/V4/V1/A1/M1/c1 ),
    .A2(\V4/V4/V1/A1/M1/c2 ),
    .ZN(\V4/V4/V1/A1/c1 ));
 AND2_X1 \V4/V4/V1/A1/M2/M1/_0_  (.A1(\V4/V4/V1/v2 [1]),
    .A2(\V4/V4/V1/v3 [1]),
    .ZN(\V4/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M2/M1/_1_  (.A(\V4/V4/V1/v2 [1]),
    .B(\V4/V4/V1/v3 [1]),
    .Z(\V4/V4/V1/A1/M2/s1 ));
 AND2_X1 \V4/V4/V1/A1/M2/M2/_0_  (.A1(\V4/V4/V1/A1/M2/s1 ),
    .A2(\V4/V4/V1/A1/c1 ),
    .ZN(\V4/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M2/M2/_1_  (.A(\V4/V4/V1/A1/M2/s1 ),
    .B(\V4/V4/V1/A1/c1 ),
    .Z(\V4/V4/V1/s1 [1]));
 OR2_X1 \V4/V4/V1/A1/M2/_0_  (.A1(\V4/V4/V1/A1/M2/c1 ),
    .A2(\V4/V4/V1/A1/M2/c2 ),
    .ZN(\V4/V4/V1/A1/c2 ));
 AND2_X1 \V4/V4/V1/A1/M3/M1/_0_  (.A1(\V4/V4/V1/v2 [2]),
    .A2(\V4/V4/V1/v3 [2]),
    .ZN(\V4/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M3/M1/_1_  (.A(\V4/V4/V1/v2 [2]),
    .B(\V4/V4/V1/v3 [2]),
    .Z(\V4/V4/V1/A1/M3/s1 ));
 AND2_X1 \V4/V4/V1/A1/M3/M2/_0_  (.A1(\V4/V4/V1/A1/M3/s1 ),
    .A2(\V4/V4/V1/A1/c2 ),
    .ZN(\V4/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M3/M2/_1_  (.A(\V4/V4/V1/A1/M3/s1 ),
    .B(\V4/V4/V1/A1/c2 ),
    .Z(\V4/V4/V1/s1 [2]));
 OR2_X1 \V4/V4/V1/A1/M3/_0_  (.A1(\V4/V4/V1/A1/M3/c1 ),
    .A2(\V4/V4/V1/A1/M3/c2 ),
    .ZN(\V4/V4/V1/A1/c3 ));
 AND2_X1 \V4/V4/V1/A1/M4/M1/_0_  (.A1(\V4/V4/V1/v2 [3]),
    .A2(\V4/V4/V1/v3 [3]),
    .ZN(\V4/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M4/M1/_1_  (.A(\V4/V4/V1/v2 [3]),
    .B(\V4/V4/V1/v3 [3]),
    .Z(\V4/V4/V1/A1/M4/s1 ));
 AND2_X1 \V4/V4/V1/A1/M4/M2/_0_  (.A1(\V4/V4/V1/A1/M4/s1 ),
    .A2(\V4/V4/V1/A1/c3 ),
    .ZN(\V4/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M4/M2/_1_  (.A(\V4/V4/V1/A1/M4/s1 ),
    .B(\V4/V4/V1/A1/c3 ),
    .Z(\V4/V4/V1/s1 [3]));
 OR2_X1 \V4/V4/V1/A1/M4/_0_  (.A1(\V4/V4/V1/A1/M4/c1 ),
    .A2(\V4/V4/V1/A1/M4/c2 ),
    .ZN(\V4/V4/V1/c1 ));
 AND2_X1 \V4/V4/V1/A2/M1/M1/_0_  (.A1(\V4/V4/V1/s1 [0]),
    .A2(\V4/V4/V1/v1 [2]),
    .ZN(\V4/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M1/M1/_1_  (.A(\V4/V4/V1/s1 [0]),
    .B(\V4/V4/V1/v1 [2]),
    .Z(\V4/V4/V1/A2/M1/s1 ));
 AND2_X1 \V4/V4/V1/A2/M1/M2/_0_  (.A1(\V4/V4/V1/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M1/M2/_1_  (.A(\V4/V4/V1/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/v4 [2]));
 OR2_X1 \V4/V4/V1/A2/M1/_0_  (.A1(\V4/V4/V1/A2/M1/c1 ),
    .A2(\V4/V4/V1/A2/M1/c2 ),
    .ZN(\V4/V4/V1/A2/c1 ));
 AND2_X1 \V4/V4/V1/A2/M2/M1/_0_  (.A1(\V4/V4/V1/s1 [1]),
    .A2(\V4/V4/V1/v1 [3]),
    .ZN(\V4/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M2/M1/_1_  (.A(\V4/V4/V1/s1 [1]),
    .B(\V4/V4/V1/v1 [3]),
    .Z(\V4/V4/V1/A2/M2/s1 ));
 AND2_X1 \V4/V4/V1/A2/M2/M2/_0_  (.A1(\V4/V4/V1/A2/M2/s1 ),
    .A2(\V4/V4/V1/A2/c1 ),
    .ZN(\V4/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M2/M2/_1_  (.A(\V4/V4/V1/A2/M2/s1 ),
    .B(\V4/V4/V1/A2/c1 ),
    .Z(\V4/v4 [3]));
 OR2_X1 \V4/V4/V1/A2/M2/_0_  (.A1(\V4/V4/V1/A2/M2/c1 ),
    .A2(\V4/V4/V1/A2/M2/c2 ),
    .ZN(\V4/V4/V1/A2/c2 ));
 AND2_X1 \V4/V4/V1/A2/M3/M1/_0_  (.A1(\V4/V4/V1/s1 [2]),
    .A2(ground),
    .ZN(\V4/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M3/M1/_1_  (.A(\V4/V4/V1/s1 [2]),
    .B(ground),
    .Z(\V4/V4/V1/A2/M3/s1 ));
 AND2_X1 \V4/V4/V1/A2/M3/M2/_0_  (.A1(\V4/V4/V1/A2/M3/s1 ),
    .A2(\V4/V4/V1/A2/c2 ),
    .ZN(\V4/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M3/M2/_1_  (.A(\V4/V4/V1/A2/M3/s1 ),
    .B(\V4/V4/V1/A2/c2 ),
    .Z(\V4/V4/V1/s2 [2]));
 OR2_X1 \V4/V4/V1/A2/M3/_0_  (.A1(\V4/V4/V1/A2/M3/c1 ),
    .A2(\V4/V4/V1/A2/M3/c2 ),
    .ZN(\V4/V4/V1/A2/c3 ));
 AND2_X1 \V4/V4/V1/A2/M4/M1/_0_  (.A1(\V4/V4/V1/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M4/M1/_1_  (.A(\V4/V4/V1/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V1/A2/M4/s1 ));
 AND2_X1 \V4/V4/V1/A2/M4/M2/_0_  (.A1(\V4/V4/V1/A2/M4/s1 ),
    .A2(\V4/V4/V1/A2/c3 ),
    .ZN(\V4/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M4/M2/_1_  (.A(\V4/V4/V1/A2/M4/s1 ),
    .B(\V4/V4/V1/A2/c3 ),
    .Z(\V4/V4/V1/s2 [3]));
 OR2_X1 \V4/V4/V1/A2/M4/_0_  (.A1(\V4/V4/V1/A2/M4/c1 ),
    .A2(\V4/V4/V1/A2/M4/c2 ),
    .ZN(\V4/V4/V1/c2 ));
 AND2_X1 \V4/V4/V1/A3/M1/M1/_0_  (.A1(\V4/V4/V1/v4 [0]),
    .A2(\V4/V4/V1/s2 [2]),
    .ZN(\V4/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M1/M1/_1_  (.A(\V4/V4/V1/v4 [0]),
    .B(\V4/V4/V1/s2 [2]),
    .Z(\V4/V4/V1/A3/M1/s1 ));
 AND2_X1 \V4/V4/V1/A3/M1/M2/_0_  (.A1(\V4/V4/V1/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M1/M2/_1_  (.A(\V4/V4/V1/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v1 [4]));
 OR2_X1 \V4/V4/V1/A3/M1/_0_  (.A1(\V4/V4/V1/A3/M1/c1 ),
    .A2(\V4/V4/V1/A3/M1/c2 ),
    .ZN(\V4/V4/V1/A3/c1 ));
 AND2_X1 \V4/V4/V1/A3/M2/M1/_0_  (.A1(\V4/V4/V1/v4 [1]),
    .A2(\V4/V4/V1/s2 [3]),
    .ZN(\V4/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M2/M1/_1_  (.A(\V4/V4/V1/v4 [1]),
    .B(\V4/V4/V1/s2 [3]),
    .Z(\V4/V4/V1/A3/M2/s1 ));
 AND2_X1 \V4/V4/V1/A3/M2/M2/_0_  (.A1(\V4/V4/V1/A3/M2/s1 ),
    .A2(\V4/V4/V1/A3/c1 ),
    .ZN(\V4/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M2/M2/_1_  (.A(\V4/V4/V1/A3/M2/s1 ),
    .B(\V4/V4/V1/A3/c1 ),
    .Z(\V4/V4/v1 [5]));
 OR2_X1 \V4/V4/V1/A3/M2/_0_  (.A1(\V4/V4/V1/A3/M2/c1 ),
    .A2(\V4/V4/V1/A3/M2/c2 ),
    .ZN(\V4/V4/V1/A3/c2 ));
 AND2_X1 \V4/V4/V1/A3/M3/M1/_0_  (.A1(\V4/V4/V1/v4 [2]),
    .A2(\V4/V4/V1/c3 ),
    .ZN(\V4/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M3/M1/_1_  (.A(\V4/V4/V1/v4 [2]),
    .B(\V4/V4/V1/c3 ),
    .Z(\V4/V4/V1/A3/M3/s1 ));
 AND2_X1 \V4/V4/V1/A3/M3/M2/_0_  (.A1(\V4/V4/V1/A3/M3/s1 ),
    .A2(\V4/V4/V1/A3/c2 ),
    .ZN(\V4/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M3/M2/_1_  (.A(\V4/V4/V1/A3/M3/s1 ),
    .B(\V4/V4/V1/A3/c2 ),
    .Z(\V4/V4/v1 [6]));
 OR2_X1 \V4/V4/V1/A3/M3/_0_  (.A1(\V4/V4/V1/A3/M3/c1 ),
    .A2(\V4/V4/V1/A3/M3/c2 ),
    .ZN(\V4/V4/V1/A3/c3 ));
 AND2_X1 \V4/V4/V1/A3/M4/M1/_0_  (.A1(\V4/V4/V1/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M4/M1/_1_  (.A(\V4/V4/V1/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V1/A3/M4/s1 ));
 AND2_X1 \V4/V4/V1/A3/M4/M2/_0_  (.A1(\V4/V4/V1/A3/M4/s1 ),
    .A2(\V4/V4/V1/A3/c3 ),
    .ZN(\V4/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M4/M2/_1_  (.A(\V4/V4/V1/A3/M4/s1 ),
    .B(\V4/V4/V1/A3/c3 ),
    .Z(\V4/V4/v1 [7]));
 OR2_X1 \V4/V4/V1/A3/M4/_0_  (.A1(\V4/V4/V1/A3/M4/c1 ),
    .A2(\V4/V4/V1/A3/M4/c2 ),
    .ZN(\V4/V4/V1/overflow ));
 AND2_X1 \V4/V4/V1/V1/HA1/_0_  (.A1(\V4/V4/V1/V1/w2 ),
    .A2(\V4/V4/V1/V1/w1 ),
    .ZN(\V4/V4/V1/V1/w4 ));
 XOR2_X2 \V4/V4/V1/V1/HA1/_1_  (.A(\V4/V4/V1/V1/w2 ),
    .B(\V4/V4/V1/V1/w1 ),
    .Z(\V4/v4 [1]));
 AND2_X1 \V4/V4/V1/V1/HA2/_0_  (.A1(\V4/V4/V1/V1/w4 ),
    .A2(\V4/V4/V1/V1/w3 ),
    .ZN(\V4/V4/V1/v1 [3]));
 XOR2_X2 \V4/V4/V1/V1/HA2/_1_  (.A(\V4/V4/V1/V1/w4 ),
    .B(\V4/V4/V1/V1/w3 ),
    .Z(\V4/V4/V1/v1 [2]));
 AND2_X1 \V4/V4/V1/V1/_0_  (.A1(A[24]),
    .A2(B[24]),
    .ZN(\V4/v4 [0]));
 AND2_X1 \V4/V4/V1/V1/_1_  (.A1(A[24]),
    .A2(B[25]),
    .ZN(\V4/V4/V1/V1/w1 ));
 AND2_X1 \V4/V4/V1/V1/_2_  (.A1(B[24]),
    .A2(A[25]),
    .ZN(\V4/V4/V1/V1/w2 ));
 AND2_X1 \V4/V4/V1/V1/_3_  (.A1(B[25]),
    .A2(A[25]),
    .ZN(\V4/V4/V1/V1/w3 ));
 AND2_X1 \V4/V4/V1/V2/HA1/_0_  (.A1(\V4/V4/V1/V2/w2 ),
    .A2(\V4/V4/V1/V2/w1 ),
    .ZN(\V4/V4/V1/V2/w4 ));
 XOR2_X2 \V4/V4/V1/V2/HA1/_1_  (.A(\V4/V4/V1/V2/w2 ),
    .B(\V4/V4/V1/V2/w1 ),
    .Z(\V4/V4/V1/v2 [1]));
 AND2_X1 \V4/V4/V1/V2/HA2/_0_  (.A1(\V4/V4/V1/V2/w4 ),
    .A2(\V4/V4/V1/V2/w3 ),
    .ZN(\V4/V4/V1/v2 [3]));
 XOR2_X2 \V4/V4/V1/V2/HA2/_1_  (.A(\V4/V4/V1/V2/w4 ),
    .B(\V4/V4/V1/V2/w3 ),
    .Z(\V4/V4/V1/v2 [2]));
 AND2_X1 \V4/V4/V1/V2/_0_  (.A1(A[26]),
    .A2(B[24]),
    .ZN(\V4/V4/V1/v2 [0]));
 AND2_X1 \V4/V4/V1/V2/_1_  (.A1(A[26]),
    .A2(B[25]),
    .ZN(\V4/V4/V1/V2/w1 ));
 AND2_X1 \V4/V4/V1/V2/_2_  (.A1(B[24]),
    .A2(A[27]),
    .ZN(\V4/V4/V1/V2/w2 ));
 AND2_X1 \V4/V4/V1/V2/_3_  (.A1(B[25]),
    .A2(A[27]),
    .ZN(\V4/V4/V1/V2/w3 ));
 AND2_X1 \V4/V4/V1/V3/HA1/_0_  (.A1(\V4/V4/V1/V3/w2 ),
    .A2(\V4/V4/V1/V3/w1 ),
    .ZN(\V4/V4/V1/V3/w4 ));
 XOR2_X2 \V4/V4/V1/V3/HA1/_1_  (.A(\V4/V4/V1/V3/w2 ),
    .B(\V4/V4/V1/V3/w1 ),
    .Z(\V4/V4/V1/v3 [1]));
 AND2_X1 \V4/V4/V1/V3/HA2/_0_  (.A1(\V4/V4/V1/V3/w4 ),
    .A2(\V4/V4/V1/V3/w3 ),
    .ZN(\V4/V4/V1/v3 [3]));
 XOR2_X2 \V4/V4/V1/V3/HA2/_1_  (.A(\V4/V4/V1/V3/w4 ),
    .B(\V4/V4/V1/V3/w3 ),
    .Z(\V4/V4/V1/v3 [2]));
 AND2_X1 \V4/V4/V1/V3/_0_  (.A1(A[24]),
    .A2(B[26]),
    .ZN(\V4/V4/V1/v3 [0]));
 AND2_X1 \V4/V4/V1/V3/_1_  (.A1(A[24]),
    .A2(B[27]),
    .ZN(\V4/V4/V1/V3/w1 ));
 AND2_X1 \V4/V4/V1/V3/_2_  (.A1(B[26]),
    .A2(A[25]),
    .ZN(\V4/V4/V1/V3/w2 ));
 AND2_X1 \V4/V4/V1/V3/_3_  (.A1(B[27]),
    .A2(A[25]),
    .ZN(\V4/V4/V1/V3/w3 ));
 AND2_X1 \V4/V4/V1/V4/HA1/_0_  (.A1(\V4/V4/V1/V4/w2 ),
    .A2(\V4/V4/V1/V4/w1 ),
    .ZN(\V4/V4/V1/V4/w4 ));
 XOR2_X2 \V4/V4/V1/V4/HA1/_1_  (.A(\V4/V4/V1/V4/w2 ),
    .B(\V4/V4/V1/V4/w1 ),
    .Z(\V4/V4/V1/v4 [1]));
 AND2_X1 \V4/V4/V1/V4/HA2/_0_  (.A1(\V4/V4/V1/V4/w4 ),
    .A2(\V4/V4/V1/V4/w3 ),
    .ZN(\V4/V4/V1/v4 [3]));
 XOR2_X2 \V4/V4/V1/V4/HA2/_1_  (.A(\V4/V4/V1/V4/w4 ),
    .B(\V4/V4/V1/V4/w3 ),
    .Z(\V4/V4/V1/v4 [2]));
 AND2_X1 \V4/V4/V1/V4/_0_  (.A1(A[26]),
    .A2(B[26]),
    .ZN(\V4/V4/V1/v4 [0]));
 AND2_X1 \V4/V4/V1/V4/_1_  (.A1(A[26]),
    .A2(B[27]),
    .ZN(\V4/V4/V1/V4/w1 ));
 AND2_X1 \V4/V4/V1/V4/_2_  (.A1(B[26]),
    .A2(A[27]),
    .ZN(\V4/V4/V1/V4/w2 ));
 AND2_X1 \V4/V4/V1/V4/_3_  (.A1(B[27]),
    .A2(A[27]),
    .ZN(\V4/V4/V1/V4/w3 ));
 OR2_X1 \V4/V4/V1/_0_  (.A1(\V4/V4/V1/c1 ),
    .A2(\V4/V4/V1/c2 ),
    .ZN(\V4/V4/V1/c3 ));
 AND2_X1 \V4/V4/V2/A1/M1/M1/_0_  (.A1(\V4/V4/V2/v2 [0]),
    .A2(\V4/V4/V2/v3 [0]),
    .ZN(\V4/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M1/M1/_1_  (.A(\V4/V4/V2/v2 [0]),
    .B(\V4/V4/V2/v3 [0]),
    .Z(\V4/V4/V2/A1/M1/s1 ));
 AND2_X1 \V4/V4/V2/A1/M1/M2/_0_  (.A1(\V4/V4/V2/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M1/M2/_1_  (.A(\V4/V4/V2/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/V2/s1 [0]));
 OR2_X1 \V4/V4/V2/A1/M1/_0_  (.A1(\V4/V4/V2/A1/M1/c1 ),
    .A2(\V4/V4/V2/A1/M1/c2 ),
    .ZN(\V4/V4/V2/A1/c1 ));
 AND2_X1 \V4/V4/V2/A1/M2/M1/_0_  (.A1(\V4/V4/V2/v2 [1]),
    .A2(\V4/V4/V2/v3 [1]),
    .ZN(\V4/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M2/M1/_1_  (.A(\V4/V4/V2/v2 [1]),
    .B(\V4/V4/V2/v3 [1]),
    .Z(\V4/V4/V2/A1/M2/s1 ));
 AND2_X1 \V4/V4/V2/A1/M2/M2/_0_  (.A1(\V4/V4/V2/A1/M2/s1 ),
    .A2(\V4/V4/V2/A1/c1 ),
    .ZN(\V4/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M2/M2/_1_  (.A(\V4/V4/V2/A1/M2/s1 ),
    .B(\V4/V4/V2/A1/c1 ),
    .Z(\V4/V4/V2/s1 [1]));
 OR2_X1 \V4/V4/V2/A1/M2/_0_  (.A1(\V4/V4/V2/A1/M2/c1 ),
    .A2(\V4/V4/V2/A1/M2/c2 ),
    .ZN(\V4/V4/V2/A1/c2 ));
 AND2_X1 \V4/V4/V2/A1/M3/M1/_0_  (.A1(\V4/V4/V2/v2 [2]),
    .A2(\V4/V4/V2/v3 [2]),
    .ZN(\V4/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M3/M1/_1_  (.A(\V4/V4/V2/v2 [2]),
    .B(\V4/V4/V2/v3 [2]),
    .Z(\V4/V4/V2/A1/M3/s1 ));
 AND2_X1 \V4/V4/V2/A1/M3/M2/_0_  (.A1(\V4/V4/V2/A1/M3/s1 ),
    .A2(\V4/V4/V2/A1/c2 ),
    .ZN(\V4/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M3/M2/_1_  (.A(\V4/V4/V2/A1/M3/s1 ),
    .B(\V4/V4/V2/A1/c2 ),
    .Z(\V4/V4/V2/s1 [2]));
 OR2_X1 \V4/V4/V2/A1/M3/_0_  (.A1(\V4/V4/V2/A1/M3/c1 ),
    .A2(\V4/V4/V2/A1/M3/c2 ),
    .ZN(\V4/V4/V2/A1/c3 ));
 AND2_X1 \V4/V4/V2/A1/M4/M1/_0_  (.A1(\V4/V4/V2/v2 [3]),
    .A2(\V4/V4/V2/v3 [3]),
    .ZN(\V4/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M4/M1/_1_  (.A(\V4/V4/V2/v2 [3]),
    .B(\V4/V4/V2/v3 [3]),
    .Z(\V4/V4/V2/A1/M4/s1 ));
 AND2_X1 \V4/V4/V2/A1/M4/M2/_0_  (.A1(\V4/V4/V2/A1/M4/s1 ),
    .A2(\V4/V4/V2/A1/c3 ),
    .ZN(\V4/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M4/M2/_1_  (.A(\V4/V4/V2/A1/M4/s1 ),
    .B(\V4/V4/V2/A1/c3 ),
    .Z(\V4/V4/V2/s1 [3]));
 OR2_X1 \V4/V4/V2/A1/M4/_0_  (.A1(\V4/V4/V2/A1/M4/c1 ),
    .A2(\V4/V4/V2/A1/M4/c2 ),
    .ZN(\V4/V4/V2/c1 ));
 AND2_X1 \V4/V4/V2/A2/M1/M1/_0_  (.A1(\V4/V4/V2/s1 [0]),
    .A2(\V4/V4/V2/v1 [2]),
    .ZN(\V4/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M1/M1/_1_  (.A(\V4/V4/V2/s1 [0]),
    .B(\V4/V4/V2/v1 [2]),
    .Z(\V4/V4/V2/A2/M1/s1 ));
 AND2_X1 \V4/V4/V2/A2/M1/M2/_0_  (.A1(\V4/V4/V2/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M1/M2/_1_  (.A(\V4/V4/V2/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v2 [2]));
 OR2_X1 \V4/V4/V2/A2/M1/_0_  (.A1(\V4/V4/V2/A2/M1/c1 ),
    .A2(\V4/V4/V2/A2/M1/c2 ),
    .ZN(\V4/V4/V2/A2/c1 ));
 AND2_X1 \V4/V4/V2/A2/M2/M1/_0_  (.A1(\V4/V4/V2/s1 [1]),
    .A2(\V4/V4/V2/v1 [3]),
    .ZN(\V4/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M2/M1/_1_  (.A(\V4/V4/V2/s1 [1]),
    .B(\V4/V4/V2/v1 [3]),
    .Z(\V4/V4/V2/A2/M2/s1 ));
 AND2_X1 \V4/V4/V2/A2/M2/M2/_0_  (.A1(\V4/V4/V2/A2/M2/s1 ),
    .A2(\V4/V4/V2/A2/c1 ),
    .ZN(\V4/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M2/M2/_1_  (.A(\V4/V4/V2/A2/M2/s1 ),
    .B(\V4/V4/V2/A2/c1 ),
    .Z(\V4/V4/v2 [3]));
 OR2_X1 \V4/V4/V2/A2/M2/_0_  (.A1(\V4/V4/V2/A2/M2/c1 ),
    .A2(\V4/V4/V2/A2/M2/c2 ),
    .ZN(\V4/V4/V2/A2/c2 ));
 AND2_X1 \V4/V4/V2/A2/M3/M1/_0_  (.A1(\V4/V4/V2/s1 [2]),
    .A2(ground),
    .ZN(\V4/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M3/M1/_1_  (.A(\V4/V4/V2/s1 [2]),
    .B(ground),
    .Z(\V4/V4/V2/A2/M3/s1 ));
 AND2_X1 \V4/V4/V2/A2/M3/M2/_0_  (.A1(\V4/V4/V2/A2/M3/s1 ),
    .A2(\V4/V4/V2/A2/c2 ),
    .ZN(\V4/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M3/M2/_1_  (.A(\V4/V4/V2/A2/M3/s1 ),
    .B(\V4/V4/V2/A2/c2 ),
    .Z(\V4/V4/V2/s2 [2]));
 OR2_X1 \V4/V4/V2/A2/M3/_0_  (.A1(\V4/V4/V2/A2/M3/c1 ),
    .A2(\V4/V4/V2/A2/M3/c2 ),
    .ZN(\V4/V4/V2/A2/c3 ));
 AND2_X1 \V4/V4/V2/A2/M4/M1/_0_  (.A1(\V4/V4/V2/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M4/M1/_1_  (.A(\V4/V4/V2/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V2/A2/M4/s1 ));
 AND2_X1 \V4/V4/V2/A2/M4/M2/_0_  (.A1(\V4/V4/V2/A2/M4/s1 ),
    .A2(\V4/V4/V2/A2/c3 ),
    .ZN(\V4/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M4/M2/_1_  (.A(\V4/V4/V2/A2/M4/s1 ),
    .B(\V4/V4/V2/A2/c3 ),
    .Z(\V4/V4/V2/s2 [3]));
 OR2_X1 \V4/V4/V2/A2/M4/_0_  (.A1(\V4/V4/V2/A2/M4/c1 ),
    .A2(\V4/V4/V2/A2/M4/c2 ),
    .ZN(\V4/V4/V2/c2 ));
 AND2_X1 \V4/V4/V2/A3/M1/M1/_0_  (.A1(\V4/V4/V2/v4 [0]),
    .A2(\V4/V4/V2/s2 [2]),
    .ZN(\V4/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M1/M1/_1_  (.A(\V4/V4/V2/v4 [0]),
    .B(\V4/V4/V2/s2 [2]),
    .Z(\V4/V4/V2/A3/M1/s1 ));
 AND2_X1 \V4/V4/V2/A3/M1/M2/_0_  (.A1(\V4/V4/V2/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M1/M2/_1_  (.A(\V4/V4/V2/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v2 [4]));
 OR2_X1 \V4/V4/V2/A3/M1/_0_  (.A1(\V4/V4/V2/A3/M1/c1 ),
    .A2(\V4/V4/V2/A3/M1/c2 ),
    .ZN(\V4/V4/V2/A3/c1 ));
 AND2_X1 \V4/V4/V2/A3/M2/M1/_0_  (.A1(\V4/V4/V2/v4 [1]),
    .A2(\V4/V4/V2/s2 [3]),
    .ZN(\V4/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M2/M1/_1_  (.A(\V4/V4/V2/v4 [1]),
    .B(\V4/V4/V2/s2 [3]),
    .Z(\V4/V4/V2/A3/M2/s1 ));
 AND2_X1 \V4/V4/V2/A3/M2/M2/_0_  (.A1(\V4/V4/V2/A3/M2/s1 ),
    .A2(\V4/V4/V2/A3/c1 ),
    .ZN(\V4/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M2/M2/_1_  (.A(\V4/V4/V2/A3/M2/s1 ),
    .B(\V4/V4/V2/A3/c1 ),
    .Z(\V4/V4/v2 [5]));
 OR2_X1 \V4/V4/V2/A3/M2/_0_  (.A1(\V4/V4/V2/A3/M2/c1 ),
    .A2(\V4/V4/V2/A3/M2/c2 ),
    .ZN(\V4/V4/V2/A3/c2 ));
 AND2_X1 \V4/V4/V2/A3/M3/M1/_0_  (.A1(\V4/V4/V2/v4 [2]),
    .A2(\V4/V4/V2/c3 ),
    .ZN(\V4/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M3/M1/_1_  (.A(\V4/V4/V2/v4 [2]),
    .B(\V4/V4/V2/c3 ),
    .Z(\V4/V4/V2/A3/M3/s1 ));
 AND2_X1 \V4/V4/V2/A3/M3/M2/_0_  (.A1(\V4/V4/V2/A3/M3/s1 ),
    .A2(\V4/V4/V2/A3/c2 ),
    .ZN(\V4/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M3/M2/_1_  (.A(\V4/V4/V2/A3/M3/s1 ),
    .B(\V4/V4/V2/A3/c2 ),
    .Z(\V4/V4/v2 [6]));
 OR2_X1 \V4/V4/V2/A3/M3/_0_  (.A1(\V4/V4/V2/A3/M3/c1 ),
    .A2(\V4/V4/V2/A3/M3/c2 ),
    .ZN(\V4/V4/V2/A3/c3 ));
 AND2_X1 \V4/V4/V2/A3/M4/M1/_0_  (.A1(\V4/V4/V2/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M4/M1/_1_  (.A(\V4/V4/V2/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V2/A3/M4/s1 ));
 AND2_X1 \V4/V4/V2/A3/M4/M2/_0_  (.A1(\V4/V4/V2/A3/M4/s1 ),
    .A2(\V4/V4/V2/A3/c3 ),
    .ZN(\V4/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M4/M2/_1_  (.A(\V4/V4/V2/A3/M4/s1 ),
    .B(\V4/V4/V2/A3/c3 ),
    .Z(\V4/V4/v2 [7]));
 OR2_X1 \V4/V4/V2/A3/M4/_0_  (.A1(\V4/V4/V2/A3/M4/c1 ),
    .A2(\V4/V4/V2/A3/M4/c2 ),
    .ZN(\V4/V4/V2/overflow ));
 AND2_X1 \V4/V4/V2/V1/HA1/_0_  (.A1(\V4/V4/V2/V1/w2 ),
    .A2(\V4/V4/V2/V1/w1 ),
    .ZN(\V4/V4/V2/V1/w4 ));
 XOR2_X2 \V4/V4/V2/V1/HA1/_1_  (.A(\V4/V4/V2/V1/w2 ),
    .B(\V4/V4/V2/V1/w1 ),
    .Z(\V4/V4/v2 [1]));
 AND2_X1 \V4/V4/V2/V1/HA2/_0_  (.A1(\V4/V4/V2/V1/w4 ),
    .A2(\V4/V4/V2/V1/w3 ),
    .ZN(\V4/V4/V2/v1 [3]));
 XOR2_X2 \V4/V4/V2/V1/HA2/_1_  (.A(\V4/V4/V2/V1/w4 ),
    .B(\V4/V4/V2/V1/w3 ),
    .Z(\V4/V4/V2/v1 [2]));
 AND2_X1 \V4/V4/V2/V1/_0_  (.A1(A[28]),
    .A2(B[24]),
    .ZN(\V4/V4/v2 [0]));
 AND2_X1 \V4/V4/V2/V1/_1_  (.A1(A[28]),
    .A2(B[25]),
    .ZN(\V4/V4/V2/V1/w1 ));
 AND2_X1 \V4/V4/V2/V1/_2_  (.A1(B[24]),
    .A2(A[29]),
    .ZN(\V4/V4/V2/V1/w2 ));
 AND2_X1 \V4/V4/V2/V1/_3_  (.A1(B[25]),
    .A2(A[29]),
    .ZN(\V4/V4/V2/V1/w3 ));
 AND2_X1 \V4/V4/V2/V2/HA1/_0_  (.A1(\V4/V4/V2/V2/w2 ),
    .A2(\V4/V4/V2/V2/w1 ),
    .ZN(\V4/V4/V2/V2/w4 ));
 XOR2_X2 \V4/V4/V2/V2/HA1/_1_  (.A(\V4/V4/V2/V2/w2 ),
    .B(\V4/V4/V2/V2/w1 ),
    .Z(\V4/V4/V2/v2 [1]));
 AND2_X1 \V4/V4/V2/V2/HA2/_0_  (.A1(\V4/V4/V2/V2/w4 ),
    .A2(\V4/V4/V2/V2/w3 ),
    .ZN(\V4/V4/V2/v2 [3]));
 XOR2_X2 \V4/V4/V2/V2/HA2/_1_  (.A(\V4/V4/V2/V2/w4 ),
    .B(\V4/V4/V2/V2/w3 ),
    .Z(\V4/V4/V2/v2 [2]));
 AND2_X1 \V4/V4/V2/V2/_0_  (.A1(A[30]),
    .A2(B[24]),
    .ZN(\V4/V4/V2/v2 [0]));
 AND2_X1 \V4/V4/V2/V2/_1_  (.A1(A[30]),
    .A2(B[25]),
    .ZN(\V4/V4/V2/V2/w1 ));
 AND2_X1 \V4/V4/V2/V2/_2_  (.A1(B[24]),
    .A2(A[31]),
    .ZN(\V4/V4/V2/V2/w2 ));
 AND2_X1 \V4/V4/V2/V2/_3_  (.A1(B[25]),
    .A2(A[31]),
    .ZN(\V4/V4/V2/V2/w3 ));
 AND2_X1 \V4/V4/V2/V3/HA1/_0_  (.A1(\V4/V4/V2/V3/w2 ),
    .A2(\V4/V4/V2/V3/w1 ),
    .ZN(\V4/V4/V2/V3/w4 ));
 XOR2_X2 \V4/V4/V2/V3/HA1/_1_  (.A(\V4/V4/V2/V3/w2 ),
    .B(\V4/V4/V2/V3/w1 ),
    .Z(\V4/V4/V2/v3 [1]));
 AND2_X1 \V4/V4/V2/V3/HA2/_0_  (.A1(\V4/V4/V2/V3/w4 ),
    .A2(\V4/V4/V2/V3/w3 ),
    .ZN(\V4/V4/V2/v3 [3]));
 XOR2_X2 \V4/V4/V2/V3/HA2/_1_  (.A(\V4/V4/V2/V3/w4 ),
    .B(\V4/V4/V2/V3/w3 ),
    .Z(\V4/V4/V2/v3 [2]));
 AND2_X1 \V4/V4/V2/V3/_0_  (.A1(A[28]),
    .A2(B[26]),
    .ZN(\V4/V4/V2/v3 [0]));
 AND2_X1 \V4/V4/V2/V3/_1_  (.A1(A[28]),
    .A2(B[27]),
    .ZN(\V4/V4/V2/V3/w1 ));
 AND2_X1 \V4/V4/V2/V3/_2_  (.A1(B[26]),
    .A2(A[29]),
    .ZN(\V4/V4/V2/V3/w2 ));
 AND2_X1 \V4/V4/V2/V3/_3_  (.A1(B[27]),
    .A2(A[29]),
    .ZN(\V4/V4/V2/V3/w3 ));
 AND2_X1 \V4/V4/V2/V4/HA1/_0_  (.A1(\V4/V4/V2/V4/w2 ),
    .A2(\V4/V4/V2/V4/w1 ),
    .ZN(\V4/V4/V2/V4/w4 ));
 XOR2_X2 \V4/V4/V2/V4/HA1/_1_  (.A(\V4/V4/V2/V4/w2 ),
    .B(\V4/V4/V2/V4/w1 ),
    .Z(\V4/V4/V2/v4 [1]));
 AND2_X1 \V4/V4/V2/V4/HA2/_0_  (.A1(\V4/V4/V2/V4/w4 ),
    .A2(\V4/V4/V2/V4/w3 ),
    .ZN(\V4/V4/V2/v4 [3]));
 XOR2_X2 \V4/V4/V2/V4/HA2/_1_  (.A(\V4/V4/V2/V4/w4 ),
    .B(\V4/V4/V2/V4/w3 ),
    .Z(\V4/V4/V2/v4 [2]));
 AND2_X1 \V4/V4/V2/V4/_0_  (.A1(A[30]),
    .A2(B[26]),
    .ZN(\V4/V4/V2/v4 [0]));
 AND2_X1 \V4/V4/V2/V4/_1_  (.A1(A[30]),
    .A2(B[27]),
    .ZN(\V4/V4/V2/V4/w1 ));
 AND2_X1 \V4/V4/V2/V4/_2_  (.A1(B[26]),
    .A2(A[31]),
    .ZN(\V4/V4/V2/V4/w2 ));
 AND2_X1 \V4/V4/V2/V4/_3_  (.A1(B[27]),
    .A2(A[31]),
    .ZN(\V4/V4/V2/V4/w3 ));
 OR2_X1 \V4/V4/V2/_0_  (.A1(\V4/V4/V2/c1 ),
    .A2(\V4/V4/V2/c2 ),
    .ZN(\V4/V4/V2/c3 ));
 AND2_X1 \V4/V4/V3/A1/M1/M1/_0_  (.A1(\V4/V4/V3/v2 [0]),
    .A2(\V4/V4/V3/v3 [0]),
    .ZN(\V4/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M1/M1/_1_  (.A(\V4/V4/V3/v2 [0]),
    .B(\V4/V4/V3/v3 [0]),
    .Z(\V4/V4/V3/A1/M1/s1 ));
 AND2_X1 \V4/V4/V3/A1/M1/M2/_0_  (.A1(\V4/V4/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M1/M2/_1_  (.A(\V4/V4/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/V3/s1 [0]));
 OR2_X1 \V4/V4/V3/A1/M1/_0_  (.A1(\V4/V4/V3/A1/M1/c1 ),
    .A2(\V4/V4/V3/A1/M1/c2 ),
    .ZN(\V4/V4/V3/A1/c1 ));
 AND2_X1 \V4/V4/V3/A1/M2/M1/_0_  (.A1(\V4/V4/V3/v2 [1]),
    .A2(\V4/V4/V3/v3 [1]),
    .ZN(\V4/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M2/M1/_1_  (.A(\V4/V4/V3/v2 [1]),
    .B(\V4/V4/V3/v3 [1]),
    .Z(\V4/V4/V3/A1/M2/s1 ));
 AND2_X1 \V4/V4/V3/A1/M2/M2/_0_  (.A1(\V4/V4/V3/A1/M2/s1 ),
    .A2(\V4/V4/V3/A1/c1 ),
    .ZN(\V4/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M2/M2/_1_  (.A(\V4/V4/V3/A1/M2/s1 ),
    .B(\V4/V4/V3/A1/c1 ),
    .Z(\V4/V4/V3/s1 [1]));
 OR2_X1 \V4/V4/V3/A1/M2/_0_  (.A1(\V4/V4/V3/A1/M2/c1 ),
    .A2(\V4/V4/V3/A1/M2/c2 ),
    .ZN(\V4/V4/V3/A1/c2 ));
 AND2_X1 \V4/V4/V3/A1/M3/M1/_0_  (.A1(\V4/V4/V3/v2 [2]),
    .A2(\V4/V4/V3/v3 [2]),
    .ZN(\V4/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M3/M1/_1_  (.A(\V4/V4/V3/v2 [2]),
    .B(\V4/V4/V3/v3 [2]),
    .Z(\V4/V4/V3/A1/M3/s1 ));
 AND2_X1 \V4/V4/V3/A1/M3/M2/_0_  (.A1(\V4/V4/V3/A1/M3/s1 ),
    .A2(\V4/V4/V3/A1/c2 ),
    .ZN(\V4/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M3/M2/_1_  (.A(\V4/V4/V3/A1/M3/s1 ),
    .B(\V4/V4/V3/A1/c2 ),
    .Z(\V4/V4/V3/s1 [2]));
 OR2_X1 \V4/V4/V3/A1/M3/_0_  (.A1(\V4/V4/V3/A1/M3/c1 ),
    .A2(\V4/V4/V3/A1/M3/c2 ),
    .ZN(\V4/V4/V3/A1/c3 ));
 AND2_X1 \V4/V4/V3/A1/M4/M1/_0_  (.A1(\V4/V4/V3/v2 [3]),
    .A2(\V4/V4/V3/v3 [3]),
    .ZN(\V4/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M4/M1/_1_  (.A(\V4/V4/V3/v2 [3]),
    .B(\V4/V4/V3/v3 [3]),
    .Z(\V4/V4/V3/A1/M4/s1 ));
 AND2_X1 \V4/V4/V3/A1/M4/M2/_0_  (.A1(\V4/V4/V3/A1/M4/s1 ),
    .A2(\V4/V4/V3/A1/c3 ),
    .ZN(\V4/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M4/M2/_1_  (.A(\V4/V4/V3/A1/M4/s1 ),
    .B(\V4/V4/V3/A1/c3 ),
    .Z(\V4/V4/V3/s1 [3]));
 OR2_X1 \V4/V4/V3/A1/M4/_0_  (.A1(\V4/V4/V3/A1/M4/c1 ),
    .A2(\V4/V4/V3/A1/M4/c2 ),
    .ZN(\V4/V4/V3/c1 ));
 AND2_X1 \V4/V4/V3/A2/M1/M1/_0_  (.A1(\V4/V4/V3/s1 [0]),
    .A2(\V4/V4/V3/v1 [2]),
    .ZN(\V4/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M1/M1/_1_  (.A(\V4/V4/V3/s1 [0]),
    .B(\V4/V4/V3/v1 [2]),
    .Z(\V4/V4/V3/A2/M1/s1 ));
 AND2_X1 \V4/V4/V3/A2/M1/M2/_0_  (.A1(\V4/V4/V3/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M1/M2/_1_  (.A(\V4/V4/V3/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v3 [2]));
 OR2_X1 \V4/V4/V3/A2/M1/_0_  (.A1(\V4/V4/V3/A2/M1/c1 ),
    .A2(\V4/V4/V3/A2/M1/c2 ),
    .ZN(\V4/V4/V3/A2/c1 ));
 AND2_X1 \V4/V4/V3/A2/M2/M1/_0_  (.A1(\V4/V4/V3/s1 [1]),
    .A2(\V4/V4/V3/v1 [3]),
    .ZN(\V4/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M2/M1/_1_  (.A(\V4/V4/V3/s1 [1]),
    .B(\V4/V4/V3/v1 [3]),
    .Z(\V4/V4/V3/A2/M2/s1 ));
 AND2_X1 \V4/V4/V3/A2/M2/M2/_0_  (.A1(\V4/V4/V3/A2/M2/s1 ),
    .A2(\V4/V4/V3/A2/c1 ),
    .ZN(\V4/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M2/M2/_1_  (.A(\V4/V4/V3/A2/M2/s1 ),
    .B(\V4/V4/V3/A2/c1 ),
    .Z(\V4/V4/v3 [3]));
 OR2_X1 \V4/V4/V3/A2/M2/_0_  (.A1(\V4/V4/V3/A2/M2/c1 ),
    .A2(\V4/V4/V3/A2/M2/c2 ),
    .ZN(\V4/V4/V3/A2/c2 ));
 AND2_X1 \V4/V4/V3/A2/M3/M1/_0_  (.A1(\V4/V4/V3/s1 [2]),
    .A2(ground),
    .ZN(\V4/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M3/M1/_1_  (.A(\V4/V4/V3/s1 [2]),
    .B(ground),
    .Z(\V4/V4/V3/A2/M3/s1 ));
 AND2_X1 \V4/V4/V3/A2/M3/M2/_0_  (.A1(\V4/V4/V3/A2/M3/s1 ),
    .A2(\V4/V4/V3/A2/c2 ),
    .ZN(\V4/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M3/M2/_1_  (.A(\V4/V4/V3/A2/M3/s1 ),
    .B(\V4/V4/V3/A2/c2 ),
    .Z(\V4/V4/V3/s2 [2]));
 OR2_X1 \V4/V4/V3/A2/M3/_0_  (.A1(\V4/V4/V3/A2/M3/c1 ),
    .A2(\V4/V4/V3/A2/M3/c2 ),
    .ZN(\V4/V4/V3/A2/c3 ));
 AND2_X1 \V4/V4/V3/A2/M4/M1/_0_  (.A1(\V4/V4/V3/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M4/M1/_1_  (.A(\V4/V4/V3/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V3/A2/M4/s1 ));
 AND2_X1 \V4/V4/V3/A2/M4/M2/_0_  (.A1(\V4/V4/V3/A2/M4/s1 ),
    .A2(\V4/V4/V3/A2/c3 ),
    .ZN(\V4/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M4/M2/_1_  (.A(\V4/V4/V3/A2/M4/s1 ),
    .B(\V4/V4/V3/A2/c3 ),
    .Z(\V4/V4/V3/s2 [3]));
 OR2_X1 \V4/V4/V3/A2/M4/_0_  (.A1(\V4/V4/V3/A2/M4/c1 ),
    .A2(\V4/V4/V3/A2/M4/c2 ),
    .ZN(\V4/V4/V3/c2 ));
 AND2_X1 \V4/V4/V3/A3/M1/M1/_0_  (.A1(\V4/V4/V3/v4 [0]),
    .A2(\V4/V4/V3/s2 [2]),
    .ZN(\V4/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M1/M1/_1_  (.A(\V4/V4/V3/v4 [0]),
    .B(\V4/V4/V3/s2 [2]),
    .Z(\V4/V4/V3/A3/M1/s1 ));
 AND2_X1 \V4/V4/V3/A3/M1/M2/_0_  (.A1(\V4/V4/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M1/M2/_1_  (.A(\V4/V4/V3/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v3 [4]));
 OR2_X1 \V4/V4/V3/A3/M1/_0_  (.A1(\V4/V4/V3/A3/M1/c1 ),
    .A2(\V4/V4/V3/A3/M1/c2 ),
    .ZN(\V4/V4/V3/A3/c1 ));
 AND2_X1 \V4/V4/V3/A3/M2/M1/_0_  (.A1(\V4/V4/V3/v4 [1]),
    .A2(\V4/V4/V3/s2 [3]),
    .ZN(\V4/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M2/M1/_1_  (.A(\V4/V4/V3/v4 [1]),
    .B(\V4/V4/V3/s2 [3]),
    .Z(\V4/V4/V3/A3/M2/s1 ));
 AND2_X1 \V4/V4/V3/A3/M2/M2/_0_  (.A1(\V4/V4/V3/A3/M2/s1 ),
    .A2(\V4/V4/V3/A3/c1 ),
    .ZN(\V4/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M2/M2/_1_  (.A(\V4/V4/V3/A3/M2/s1 ),
    .B(\V4/V4/V3/A3/c1 ),
    .Z(\V4/V4/v3 [5]));
 OR2_X1 \V4/V4/V3/A3/M2/_0_  (.A1(\V4/V4/V3/A3/M2/c1 ),
    .A2(\V4/V4/V3/A3/M2/c2 ),
    .ZN(\V4/V4/V3/A3/c2 ));
 AND2_X1 \V4/V4/V3/A3/M3/M1/_0_  (.A1(\V4/V4/V3/v4 [2]),
    .A2(\V4/V4/V3/c3 ),
    .ZN(\V4/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M3/M1/_1_  (.A(\V4/V4/V3/v4 [2]),
    .B(\V4/V4/V3/c3 ),
    .Z(\V4/V4/V3/A3/M3/s1 ));
 AND2_X1 \V4/V4/V3/A3/M3/M2/_0_  (.A1(\V4/V4/V3/A3/M3/s1 ),
    .A2(\V4/V4/V3/A3/c2 ),
    .ZN(\V4/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M3/M2/_1_  (.A(\V4/V4/V3/A3/M3/s1 ),
    .B(\V4/V4/V3/A3/c2 ),
    .Z(\V4/V4/v3 [6]));
 OR2_X1 \V4/V4/V3/A3/M3/_0_  (.A1(\V4/V4/V3/A3/M3/c1 ),
    .A2(\V4/V4/V3/A3/M3/c2 ),
    .ZN(\V4/V4/V3/A3/c3 ));
 AND2_X1 \V4/V4/V3/A3/M4/M1/_0_  (.A1(\V4/V4/V3/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M4/M1/_1_  (.A(\V4/V4/V3/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V3/A3/M4/s1 ));
 AND2_X1 \V4/V4/V3/A3/M4/M2/_0_  (.A1(\V4/V4/V3/A3/M4/s1 ),
    .A2(\V4/V4/V3/A3/c3 ),
    .ZN(\V4/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M4/M2/_1_  (.A(\V4/V4/V3/A3/M4/s1 ),
    .B(\V4/V4/V3/A3/c3 ),
    .Z(\V4/V4/v3 [7]));
 OR2_X1 \V4/V4/V3/A3/M4/_0_  (.A1(\V4/V4/V3/A3/M4/c1 ),
    .A2(\V4/V4/V3/A3/M4/c2 ),
    .ZN(\V4/V4/V3/overflow ));
 AND2_X1 \V4/V4/V3/V1/HA1/_0_  (.A1(\V4/V4/V3/V1/w2 ),
    .A2(\V4/V4/V3/V1/w1 ),
    .ZN(\V4/V4/V3/V1/w4 ));
 XOR2_X2 \V4/V4/V3/V1/HA1/_1_  (.A(\V4/V4/V3/V1/w2 ),
    .B(\V4/V4/V3/V1/w1 ),
    .Z(\V4/V4/v3 [1]));
 AND2_X1 \V4/V4/V3/V1/HA2/_0_  (.A1(\V4/V4/V3/V1/w4 ),
    .A2(\V4/V4/V3/V1/w3 ),
    .ZN(\V4/V4/V3/v1 [3]));
 XOR2_X2 \V4/V4/V3/V1/HA2/_1_  (.A(\V4/V4/V3/V1/w4 ),
    .B(\V4/V4/V3/V1/w3 ),
    .Z(\V4/V4/V3/v1 [2]));
 AND2_X1 \V4/V4/V3/V1/_0_  (.A1(A[24]),
    .A2(B[28]),
    .ZN(\V4/V4/v3 [0]));
 AND2_X1 \V4/V4/V3/V1/_1_  (.A1(A[24]),
    .A2(B[29]),
    .ZN(\V4/V4/V3/V1/w1 ));
 AND2_X1 \V4/V4/V3/V1/_2_  (.A1(B[28]),
    .A2(A[25]),
    .ZN(\V4/V4/V3/V1/w2 ));
 AND2_X1 \V4/V4/V3/V1/_3_  (.A1(B[29]),
    .A2(A[25]),
    .ZN(\V4/V4/V3/V1/w3 ));
 AND2_X1 \V4/V4/V3/V2/HA1/_0_  (.A1(\V4/V4/V3/V2/w2 ),
    .A2(\V4/V4/V3/V2/w1 ),
    .ZN(\V4/V4/V3/V2/w4 ));
 XOR2_X2 \V4/V4/V3/V2/HA1/_1_  (.A(\V4/V4/V3/V2/w2 ),
    .B(\V4/V4/V3/V2/w1 ),
    .Z(\V4/V4/V3/v2 [1]));
 AND2_X1 \V4/V4/V3/V2/HA2/_0_  (.A1(\V4/V4/V3/V2/w4 ),
    .A2(\V4/V4/V3/V2/w3 ),
    .ZN(\V4/V4/V3/v2 [3]));
 XOR2_X2 \V4/V4/V3/V2/HA2/_1_  (.A(\V4/V4/V3/V2/w4 ),
    .B(\V4/V4/V3/V2/w3 ),
    .Z(\V4/V4/V3/v2 [2]));
 AND2_X1 \V4/V4/V3/V2/_0_  (.A1(A[26]),
    .A2(B[28]),
    .ZN(\V4/V4/V3/v2 [0]));
 AND2_X1 \V4/V4/V3/V2/_1_  (.A1(A[26]),
    .A2(B[29]),
    .ZN(\V4/V4/V3/V2/w1 ));
 AND2_X1 \V4/V4/V3/V2/_2_  (.A1(B[28]),
    .A2(A[27]),
    .ZN(\V4/V4/V3/V2/w2 ));
 AND2_X1 \V4/V4/V3/V2/_3_  (.A1(B[29]),
    .A2(A[27]),
    .ZN(\V4/V4/V3/V2/w3 ));
 AND2_X1 \V4/V4/V3/V3/HA1/_0_  (.A1(\V4/V4/V3/V3/w2 ),
    .A2(\V4/V4/V3/V3/w1 ),
    .ZN(\V4/V4/V3/V3/w4 ));
 XOR2_X2 \V4/V4/V3/V3/HA1/_1_  (.A(\V4/V4/V3/V3/w2 ),
    .B(\V4/V4/V3/V3/w1 ),
    .Z(\V4/V4/V3/v3 [1]));
 AND2_X1 \V4/V4/V3/V3/HA2/_0_  (.A1(\V4/V4/V3/V3/w4 ),
    .A2(\V4/V4/V3/V3/w3 ),
    .ZN(\V4/V4/V3/v3 [3]));
 XOR2_X2 \V4/V4/V3/V3/HA2/_1_  (.A(\V4/V4/V3/V3/w4 ),
    .B(\V4/V4/V3/V3/w3 ),
    .Z(\V4/V4/V3/v3 [2]));
 AND2_X1 \V4/V4/V3/V3/_0_  (.A1(A[24]),
    .A2(B[30]),
    .ZN(\V4/V4/V3/v3 [0]));
 AND2_X1 \V4/V4/V3/V3/_1_  (.A1(A[24]),
    .A2(B[31]),
    .ZN(\V4/V4/V3/V3/w1 ));
 AND2_X1 \V4/V4/V3/V3/_2_  (.A1(B[30]),
    .A2(A[25]),
    .ZN(\V4/V4/V3/V3/w2 ));
 AND2_X1 \V4/V4/V3/V3/_3_  (.A1(B[31]),
    .A2(A[25]),
    .ZN(\V4/V4/V3/V3/w3 ));
 AND2_X1 \V4/V4/V3/V4/HA1/_0_  (.A1(\V4/V4/V3/V4/w2 ),
    .A2(\V4/V4/V3/V4/w1 ),
    .ZN(\V4/V4/V3/V4/w4 ));
 XOR2_X2 \V4/V4/V3/V4/HA1/_1_  (.A(\V4/V4/V3/V4/w2 ),
    .B(\V4/V4/V3/V4/w1 ),
    .Z(\V4/V4/V3/v4 [1]));
 AND2_X1 \V4/V4/V3/V4/HA2/_0_  (.A1(\V4/V4/V3/V4/w4 ),
    .A2(\V4/V4/V3/V4/w3 ),
    .ZN(\V4/V4/V3/v4 [3]));
 XOR2_X2 \V4/V4/V3/V4/HA2/_1_  (.A(\V4/V4/V3/V4/w4 ),
    .B(\V4/V4/V3/V4/w3 ),
    .Z(\V4/V4/V3/v4 [2]));
 AND2_X1 \V4/V4/V3/V4/_0_  (.A1(A[26]),
    .A2(B[30]),
    .ZN(\V4/V4/V3/v4 [0]));
 AND2_X1 \V4/V4/V3/V4/_1_  (.A1(A[26]),
    .A2(B[31]),
    .ZN(\V4/V4/V3/V4/w1 ));
 AND2_X1 \V4/V4/V3/V4/_2_  (.A1(B[30]),
    .A2(A[27]),
    .ZN(\V4/V4/V3/V4/w2 ));
 AND2_X1 \V4/V4/V3/V4/_3_  (.A1(B[31]),
    .A2(A[27]),
    .ZN(\V4/V4/V3/V4/w3 ));
 OR2_X1 \V4/V4/V3/_0_  (.A1(\V4/V4/V3/c1 ),
    .A2(\V4/V4/V3/c2 ),
    .ZN(\V4/V4/V3/c3 ));
 AND2_X1 \V4/V4/V4/A1/M1/M1/_0_  (.A1(\V4/V4/V4/v2 [0]),
    .A2(\V4/V4/V4/v3 [0]),
    .ZN(\V4/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M1/M1/_1_  (.A(\V4/V4/V4/v2 [0]),
    .B(\V4/V4/V4/v3 [0]),
    .Z(\V4/V4/V4/A1/M1/s1 ));
 AND2_X1 \V4/V4/V4/A1/M1/M2/_0_  (.A1(\V4/V4/V4/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M1/M2/_1_  (.A(\V4/V4/V4/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/V4/s1 [0]));
 OR2_X1 \V4/V4/V4/A1/M1/_0_  (.A1(\V4/V4/V4/A1/M1/c1 ),
    .A2(\V4/V4/V4/A1/M1/c2 ),
    .ZN(\V4/V4/V4/A1/c1 ));
 AND2_X1 \V4/V4/V4/A1/M2/M1/_0_  (.A1(\V4/V4/V4/v2 [1]),
    .A2(\V4/V4/V4/v3 [1]),
    .ZN(\V4/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M2/M1/_1_  (.A(\V4/V4/V4/v2 [1]),
    .B(\V4/V4/V4/v3 [1]),
    .Z(\V4/V4/V4/A1/M2/s1 ));
 AND2_X1 \V4/V4/V4/A1/M2/M2/_0_  (.A1(\V4/V4/V4/A1/M2/s1 ),
    .A2(\V4/V4/V4/A1/c1 ),
    .ZN(\V4/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M2/M2/_1_  (.A(\V4/V4/V4/A1/M2/s1 ),
    .B(\V4/V4/V4/A1/c1 ),
    .Z(\V4/V4/V4/s1 [1]));
 OR2_X1 \V4/V4/V4/A1/M2/_0_  (.A1(\V4/V4/V4/A1/M2/c1 ),
    .A2(\V4/V4/V4/A1/M2/c2 ),
    .ZN(\V4/V4/V4/A1/c2 ));
 AND2_X1 \V4/V4/V4/A1/M3/M1/_0_  (.A1(\V4/V4/V4/v2 [2]),
    .A2(\V4/V4/V4/v3 [2]),
    .ZN(\V4/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M3/M1/_1_  (.A(\V4/V4/V4/v2 [2]),
    .B(\V4/V4/V4/v3 [2]),
    .Z(\V4/V4/V4/A1/M3/s1 ));
 AND2_X1 \V4/V4/V4/A1/M3/M2/_0_  (.A1(\V4/V4/V4/A1/M3/s1 ),
    .A2(\V4/V4/V4/A1/c2 ),
    .ZN(\V4/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M3/M2/_1_  (.A(\V4/V4/V4/A1/M3/s1 ),
    .B(\V4/V4/V4/A1/c2 ),
    .Z(\V4/V4/V4/s1 [2]));
 OR2_X1 \V4/V4/V4/A1/M3/_0_  (.A1(\V4/V4/V4/A1/M3/c1 ),
    .A2(\V4/V4/V4/A1/M3/c2 ),
    .ZN(\V4/V4/V4/A1/c3 ));
 AND2_X1 \V4/V4/V4/A1/M4/M1/_0_  (.A1(\V4/V4/V4/v2 [3]),
    .A2(\V4/V4/V4/v3 [3]),
    .ZN(\V4/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M4/M1/_1_  (.A(\V4/V4/V4/v2 [3]),
    .B(\V4/V4/V4/v3 [3]),
    .Z(\V4/V4/V4/A1/M4/s1 ));
 AND2_X1 \V4/V4/V4/A1/M4/M2/_0_  (.A1(\V4/V4/V4/A1/M4/s1 ),
    .A2(\V4/V4/V4/A1/c3 ),
    .ZN(\V4/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M4/M2/_1_  (.A(\V4/V4/V4/A1/M4/s1 ),
    .B(\V4/V4/V4/A1/c3 ),
    .Z(\V4/V4/V4/s1 [3]));
 OR2_X1 \V4/V4/V4/A1/M4/_0_  (.A1(\V4/V4/V4/A1/M4/c1 ),
    .A2(\V4/V4/V4/A1/M4/c2 ),
    .ZN(\V4/V4/V4/c1 ));
 AND2_X1 \V4/V4/V4/A2/M1/M1/_0_  (.A1(\V4/V4/V4/s1 [0]),
    .A2(\V4/V4/V4/v1 [2]),
    .ZN(\V4/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M1/M1/_1_  (.A(\V4/V4/V4/s1 [0]),
    .B(\V4/V4/V4/v1 [2]),
    .Z(\V4/V4/V4/A2/M1/s1 ));
 AND2_X1 \V4/V4/V4/A2/M1/M2/_0_  (.A1(\V4/V4/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M1/M2/_1_  (.A(\V4/V4/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v4 [2]));
 OR2_X1 \V4/V4/V4/A2/M1/_0_  (.A1(\V4/V4/V4/A2/M1/c1 ),
    .A2(\V4/V4/V4/A2/M1/c2 ),
    .ZN(\V4/V4/V4/A2/c1 ));
 AND2_X1 \V4/V4/V4/A2/M2/M1/_0_  (.A1(\V4/V4/V4/s1 [1]),
    .A2(\V4/V4/V4/v1 [3]),
    .ZN(\V4/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M2/M1/_1_  (.A(\V4/V4/V4/s1 [1]),
    .B(\V4/V4/V4/v1 [3]),
    .Z(\V4/V4/V4/A2/M2/s1 ));
 AND2_X1 \V4/V4/V4/A2/M2/M2/_0_  (.A1(\V4/V4/V4/A2/M2/s1 ),
    .A2(\V4/V4/V4/A2/c1 ),
    .ZN(\V4/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M2/M2/_1_  (.A(\V4/V4/V4/A2/M2/s1 ),
    .B(\V4/V4/V4/A2/c1 ),
    .Z(\V4/V4/v4 [3]));
 OR2_X1 \V4/V4/V4/A2/M2/_0_  (.A1(\V4/V4/V4/A2/M2/c1 ),
    .A2(\V4/V4/V4/A2/M2/c2 ),
    .ZN(\V4/V4/V4/A2/c2 ));
 AND2_X1 \V4/V4/V4/A2/M3/M1/_0_  (.A1(\V4/V4/V4/s1 [2]),
    .A2(ground),
    .ZN(\V4/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M3/M1/_1_  (.A(\V4/V4/V4/s1 [2]),
    .B(ground),
    .Z(\V4/V4/V4/A2/M3/s1 ));
 AND2_X1 \V4/V4/V4/A2/M3/M2/_0_  (.A1(\V4/V4/V4/A2/M3/s1 ),
    .A2(\V4/V4/V4/A2/c2 ),
    .ZN(\V4/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M3/M2/_1_  (.A(\V4/V4/V4/A2/M3/s1 ),
    .B(\V4/V4/V4/A2/c2 ),
    .Z(\V4/V4/V4/s2 [2]));
 OR2_X1 \V4/V4/V4/A2/M3/_0_  (.A1(\V4/V4/V4/A2/M3/c1 ),
    .A2(\V4/V4/V4/A2/M3/c2 ),
    .ZN(\V4/V4/V4/A2/c3 ));
 AND2_X1 \V4/V4/V4/A2/M4/M1/_0_  (.A1(\V4/V4/V4/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M4/M1/_1_  (.A(\V4/V4/V4/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V4/A2/M4/s1 ));
 AND2_X1 \V4/V4/V4/A2/M4/M2/_0_  (.A1(\V4/V4/V4/A2/M4/s1 ),
    .A2(\V4/V4/V4/A2/c3 ),
    .ZN(\V4/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M4/M2/_1_  (.A(\V4/V4/V4/A2/M4/s1 ),
    .B(\V4/V4/V4/A2/c3 ),
    .Z(\V4/V4/V4/s2 [3]));
 OR2_X1 \V4/V4/V4/A2/M4/_0_  (.A1(\V4/V4/V4/A2/M4/c1 ),
    .A2(\V4/V4/V4/A2/M4/c2 ),
    .ZN(\V4/V4/V4/c2 ));
 AND2_X1 \V4/V4/V4/A3/M1/M1/_0_  (.A1(\V4/V4/V4/v4 [0]),
    .A2(\V4/V4/V4/s2 [2]),
    .ZN(\V4/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M1/M1/_1_  (.A(\V4/V4/V4/v4 [0]),
    .B(\V4/V4/V4/s2 [2]),
    .Z(\V4/V4/V4/A3/M1/s1 ));
 AND2_X1 \V4/V4/V4/A3/M1/M2/_0_  (.A1(\V4/V4/V4/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M1/M2/_1_  (.A(\V4/V4/V4/A3/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v4 [4]));
 OR2_X1 \V4/V4/V4/A3/M1/_0_  (.A1(\V4/V4/V4/A3/M1/c1 ),
    .A2(\V4/V4/V4/A3/M1/c2 ),
    .ZN(\V4/V4/V4/A3/c1 ));
 AND2_X1 \V4/V4/V4/A3/M2/M1/_0_  (.A1(\V4/V4/V4/v4 [1]),
    .A2(\V4/V4/V4/s2 [3]),
    .ZN(\V4/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M2/M1/_1_  (.A(\V4/V4/V4/v4 [1]),
    .B(\V4/V4/V4/s2 [3]),
    .Z(\V4/V4/V4/A3/M2/s1 ));
 AND2_X1 \V4/V4/V4/A3/M2/M2/_0_  (.A1(\V4/V4/V4/A3/M2/s1 ),
    .A2(\V4/V4/V4/A3/c1 ),
    .ZN(\V4/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M2/M2/_1_  (.A(\V4/V4/V4/A3/M2/s1 ),
    .B(\V4/V4/V4/A3/c1 ),
    .Z(\V4/V4/v4 [5]));
 OR2_X1 \V4/V4/V4/A3/M2/_0_  (.A1(\V4/V4/V4/A3/M2/c1 ),
    .A2(\V4/V4/V4/A3/M2/c2 ),
    .ZN(\V4/V4/V4/A3/c2 ));
 AND2_X1 \V4/V4/V4/A3/M3/M1/_0_  (.A1(\V4/V4/V4/v4 [2]),
    .A2(\V4/V4/V4/c3 ),
    .ZN(\V4/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M3/M1/_1_  (.A(\V4/V4/V4/v4 [2]),
    .B(\V4/V4/V4/c3 ),
    .Z(\V4/V4/V4/A3/M3/s1 ));
 AND2_X1 \V4/V4/V4/A3/M3/M2/_0_  (.A1(\V4/V4/V4/A3/M3/s1 ),
    .A2(\V4/V4/V4/A3/c2 ),
    .ZN(\V4/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M3/M2/_1_  (.A(\V4/V4/V4/A3/M3/s1 ),
    .B(\V4/V4/V4/A3/c2 ),
    .Z(\V4/V4/v4 [6]));
 OR2_X1 \V4/V4/V4/A3/M3/_0_  (.A1(\V4/V4/V4/A3/M3/c1 ),
    .A2(\V4/V4/V4/A3/M3/c2 ),
    .ZN(\V4/V4/V4/A3/c3 ));
 AND2_X1 \V4/V4/V4/A3/M4/M1/_0_  (.A1(\V4/V4/V4/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M4/M1/_1_  (.A(\V4/V4/V4/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V4/A3/M4/s1 ));
 AND2_X1 \V4/V4/V4/A3/M4/M2/_0_  (.A1(\V4/V4/V4/A3/M4/s1 ),
    .A2(\V4/V4/V4/A3/c3 ),
    .ZN(\V4/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M4/M2/_1_  (.A(\V4/V4/V4/A3/M4/s1 ),
    .B(\V4/V4/V4/A3/c3 ),
    .Z(\V4/V4/v4 [7]));
 OR2_X1 \V4/V4/V4/A3/M4/_0_  (.A1(\V4/V4/V4/A3/M4/c1 ),
    .A2(\V4/V4/V4/A3/M4/c2 ),
    .ZN(\V4/V4/V4/overflow ));
 AND2_X1 \V4/V4/V4/V1/HA1/_0_  (.A1(\V4/V4/V4/V1/w2 ),
    .A2(\V4/V4/V4/V1/w1 ),
    .ZN(\V4/V4/V4/V1/w4 ));
 XOR2_X2 \V4/V4/V4/V1/HA1/_1_  (.A(\V4/V4/V4/V1/w2 ),
    .B(\V4/V4/V4/V1/w1 ),
    .Z(\V4/V4/v4 [1]));
 AND2_X1 \V4/V4/V4/V1/HA2/_0_  (.A1(\V4/V4/V4/V1/w4 ),
    .A2(\V4/V4/V4/V1/w3 ),
    .ZN(\V4/V4/V4/v1 [3]));
 XOR2_X2 \V4/V4/V4/V1/HA2/_1_  (.A(\V4/V4/V4/V1/w4 ),
    .B(\V4/V4/V4/V1/w3 ),
    .Z(\V4/V4/V4/v1 [2]));
 AND2_X1 \V4/V4/V4/V1/_0_  (.A1(A[28]),
    .A2(B[28]),
    .ZN(\V4/V4/v4 [0]));
 AND2_X1 \V4/V4/V4/V1/_1_  (.A1(A[28]),
    .A2(B[29]),
    .ZN(\V4/V4/V4/V1/w1 ));
 AND2_X1 \V4/V4/V4/V1/_2_  (.A1(B[28]),
    .A2(A[29]),
    .ZN(\V4/V4/V4/V1/w2 ));
 AND2_X1 \V4/V4/V4/V1/_3_  (.A1(B[29]),
    .A2(A[29]),
    .ZN(\V4/V4/V4/V1/w3 ));
 AND2_X1 \V4/V4/V4/V2/HA1/_0_  (.A1(\V4/V4/V4/V2/w2 ),
    .A2(\V4/V4/V4/V2/w1 ),
    .ZN(\V4/V4/V4/V2/w4 ));
 XOR2_X2 \V4/V4/V4/V2/HA1/_1_  (.A(\V4/V4/V4/V2/w2 ),
    .B(\V4/V4/V4/V2/w1 ),
    .Z(\V4/V4/V4/v2 [1]));
 AND2_X1 \V4/V4/V4/V2/HA2/_0_  (.A1(\V4/V4/V4/V2/w4 ),
    .A2(\V4/V4/V4/V2/w3 ),
    .ZN(\V4/V4/V4/v2 [3]));
 XOR2_X2 \V4/V4/V4/V2/HA2/_1_  (.A(\V4/V4/V4/V2/w4 ),
    .B(\V4/V4/V4/V2/w3 ),
    .Z(\V4/V4/V4/v2 [2]));
 AND2_X1 \V4/V4/V4/V2/_0_  (.A1(A[30]),
    .A2(B[28]),
    .ZN(\V4/V4/V4/v2 [0]));
 AND2_X1 \V4/V4/V4/V2/_1_  (.A1(A[30]),
    .A2(B[29]),
    .ZN(\V4/V4/V4/V2/w1 ));
 AND2_X1 \V4/V4/V4/V2/_2_  (.A1(B[28]),
    .A2(A[31]),
    .ZN(\V4/V4/V4/V2/w2 ));
 AND2_X1 \V4/V4/V4/V2/_3_  (.A1(B[29]),
    .A2(A[31]),
    .ZN(\V4/V4/V4/V2/w3 ));
 AND2_X1 \V4/V4/V4/V3/HA1/_0_  (.A1(\V4/V4/V4/V3/w2 ),
    .A2(\V4/V4/V4/V3/w1 ),
    .ZN(\V4/V4/V4/V3/w4 ));
 XOR2_X2 \V4/V4/V4/V3/HA1/_1_  (.A(\V4/V4/V4/V3/w2 ),
    .B(\V4/V4/V4/V3/w1 ),
    .Z(\V4/V4/V4/v3 [1]));
 AND2_X1 \V4/V4/V4/V3/HA2/_0_  (.A1(\V4/V4/V4/V3/w4 ),
    .A2(\V4/V4/V4/V3/w3 ),
    .ZN(\V4/V4/V4/v3 [3]));
 XOR2_X2 \V4/V4/V4/V3/HA2/_1_  (.A(\V4/V4/V4/V3/w4 ),
    .B(\V4/V4/V4/V3/w3 ),
    .Z(\V4/V4/V4/v3 [2]));
 AND2_X1 \V4/V4/V4/V3/_0_  (.A1(A[28]),
    .A2(B[30]),
    .ZN(\V4/V4/V4/v3 [0]));
 AND2_X1 \V4/V4/V4/V3/_1_  (.A1(A[28]),
    .A2(B[31]),
    .ZN(\V4/V4/V4/V3/w1 ));
 AND2_X1 \V4/V4/V4/V3/_2_  (.A1(B[30]),
    .A2(A[29]),
    .ZN(\V4/V4/V4/V3/w2 ));
 AND2_X1 \V4/V4/V4/V3/_3_  (.A1(B[31]),
    .A2(A[29]),
    .ZN(\V4/V4/V4/V3/w3 ));
 AND2_X1 \V4/V4/V4/V4/HA1/_0_  (.A1(\V4/V4/V4/V4/w2 ),
    .A2(\V4/V4/V4/V4/w1 ),
    .ZN(\V4/V4/V4/V4/w4 ));
 XOR2_X2 \V4/V4/V4/V4/HA1/_1_  (.A(\V4/V4/V4/V4/w2 ),
    .B(\V4/V4/V4/V4/w1 ),
    .Z(\V4/V4/V4/v4 [1]));
 AND2_X1 \V4/V4/V4/V4/HA2/_0_  (.A1(\V4/V4/V4/V4/w4 ),
    .A2(\V4/V4/V4/V4/w3 ),
    .ZN(\V4/V4/V4/v4 [3]));
 XOR2_X2 \V4/V4/V4/V4/HA2/_1_  (.A(\V4/V4/V4/V4/w4 ),
    .B(\V4/V4/V4/V4/w3 ),
    .Z(\V4/V4/V4/v4 [2]));
 AND2_X1 \V4/V4/V4/V4/_0_  (.A1(A[30]),
    .A2(B[30]),
    .ZN(\V4/V4/V4/v4 [0]));
 AND2_X1 \V4/V4/V4/V4/_1_  (.A1(A[30]),
    .A2(B[31]),
    .ZN(\V4/V4/V4/V4/w1 ));
 AND2_X1 \V4/V4/V4/V4/_2_  (.A1(B[30]),
    .A2(A[31]),
    .ZN(\V4/V4/V4/V4/w2 ));
 AND2_X1 \V4/V4/V4/V4/_3_  (.A1(B[31]),
    .A2(A[31]),
    .ZN(\V4/V4/V4/V4/w3 ));
 OR2_X1 \V4/V4/V4/_0_  (.A1(\V4/V4/V4/c1 ),
    .A2(\V4/V4/V4/c2 ),
    .ZN(\V4/V4/V4/c3 ));
 OR2_X1 \V4/V4/_0_  (.A1(\V4/V4/c1 ),
    .A2(\V4/V4/c2 ),
    .ZN(\V4/V4/c3 ));
 OR2_X1 \V4/_0_  (.A1(\V4/c1 ),
    .A2(\V4/c2 ),
    .ZN(\V4/c3 ));
 OR2_X2 _0_ (.A1(c1),
    .A2(c2),
    .ZN(c3));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_682 ();
 assign Prod[16] = s2[0];
 assign Prod[26] = s2[10];
 assign Prod[27] = s2[11];
 assign Prod[28] = s2[12];
 assign Prod[29] = s2[13];
 assign Prod[30] = s2[14];
 assign Prod[31] = s2[15];
 assign Prod[17] = s2[1];
 assign Prod[18] = s2[2];
 assign Prod[19] = s2[3];
 assign Prod[20] = s2[4];
 assign Prod[21] = s2[5];
 assign Prod[22] = s2[6];
 assign Prod[23] = s2[7];
 assign Prod[24] = s2[8];
 assign Prod[25] = s2[9];
 assign Prod[0] = v1[0];
 assign Prod[10] = v1[10];
 assign Prod[11] = v1[11];
 assign Prod[12] = v1[12];
 assign Prod[13] = v1[13];
 assign Prod[14] = v1[14];
 assign Prod[15] = v1[15];
 assign Prod[1] = v1[1];
 assign Prod[2] = v1[2];
 assign Prod[3] = v1[3];
 assign Prod[4] = v1[4];
 assign Prod[5] = v1[5];
 assign Prod[6] = v1[6];
 assign Prod[7] = v1[7];
 assign Prod[8] = v1[8];
 assign Prod[9] = v1[9];
endmodule
