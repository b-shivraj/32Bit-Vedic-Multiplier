module vedic32x32 (ground,
    overflow,
    A,
    B,
    Prod);
 input ground;
 output overflow;
 input [31:0] A;
 input [31:0] B;
 output [63:0] Prod;

 wire c1;
 wire c2;
 wire c3;
 wire \A1/c1 ;
 wire \A1/A1/c1 ;
 wire \A1/A1/A1/c1 ;
 wire \A1/A1/A1/A1/c1 ;
 wire \A1/A1/A1/A1/c2 ;
 wire \A1/A1/A1/A1/c3 ;
 wire \A1/A1/A1/A1/M1/c1 ;
 wire \A1/A1/A1/A1/M1/c2 ;
 wire \A1/A1/A1/A1/M1/s1 ;
 wire \A1/A1/A1/A1/M2/c1 ;
 wire \A1/A1/A1/A1/M2/c2 ;
 wire \A1/A1/A1/A1/M2/s1 ;
 wire \A1/A1/A1/A1/M3/c1 ;
 wire \A1/A1/A1/A1/M3/c2 ;
 wire \A1/A1/A1/A1/M3/s1 ;
 wire \A1/A1/A1/A1/M4/c1 ;
 wire \A1/A1/A1/A1/M4/c2 ;
 wire \A1/A1/A1/A1/M4/s1 ;
 wire \A1/A1/A1/A2/c1 ;
 wire \A1/A1/A1/A2/c2 ;
 wire \A1/A1/A1/A2/c3 ;
 wire \A1/A1/A1/A2/M1/c1 ;
 wire \A1/A1/A1/A2/M1/c2 ;
 wire \A1/A1/A1/A2/M1/s1 ;
 wire \A1/A1/A1/A2/M2/c1 ;
 wire \A1/A1/A1/A2/M2/c2 ;
 wire \A1/A1/A1/A2/M2/s1 ;
 wire \A1/A1/A1/A2/M3/c1 ;
 wire \A1/A1/A1/A2/M3/c2 ;
 wire \A1/A1/A1/A2/M3/s1 ;
 wire \A1/A1/A1/A2/M4/c1 ;
 wire \A1/A1/A1/A2/M4/c2 ;
 wire \A1/A1/A1/A2/M4/s1 ;
 wire \A1/A1/A2/c1 ;
 wire \A1/A1/A2/A1/c1 ;
 wire \A1/A1/A2/A1/c2 ;
 wire \A1/A1/A2/A1/c3 ;
 wire \A1/A1/A2/A1/M1/c1 ;
 wire \A1/A1/A2/A1/M1/c2 ;
 wire \A1/A1/A2/A1/M1/s1 ;
 wire \A1/A1/A2/A1/M2/c1 ;
 wire \A1/A1/A2/A1/M2/c2 ;
 wire \A1/A1/A2/A1/M2/s1 ;
 wire \A1/A1/A2/A1/M3/c1 ;
 wire \A1/A1/A2/A1/M3/c2 ;
 wire \A1/A1/A2/A1/M3/s1 ;
 wire \A1/A1/A2/A1/M4/c1 ;
 wire \A1/A1/A2/A1/M4/c2 ;
 wire \A1/A1/A2/A1/M4/s1 ;
 wire \A1/A1/A2/A2/c1 ;
 wire \A1/A1/A2/A2/c2 ;
 wire \A1/A1/A2/A2/c3 ;
 wire \A1/A1/A2/A2/M1/c1 ;
 wire \A1/A1/A2/A2/M1/c2 ;
 wire \A1/A1/A2/A2/M1/s1 ;
 wire \A1/A1/A2/A2/M2/c1 ;
 wire \A1/A1/A2/A2/M2/c2 ;
 wire \A1/A1/A2/A2/M2/s1 ;
 wire \A1/A1/A2/A2/M3/c1 ;
 wire \A1/A1/A2/A2/M3/c2 ;
 wire \A1/A1/A2/A2/M3/s1 ;
 wire \A1/A1/A2/A2/M4/c1 ;
 wire \A1/A1/A2/A2/M4/c2 ;
 wire \A1/A1/A2/A2/M4/s1 ;
 wire \A1/A2/c1 ;
 wire \A1/A2/A1/c1 ;
 wire \A1/A2/A1/A1/c1 ;
 wire \A1/A2/A1/A1/c2 ;
 wire \A1/A2/A1/A1/c3 ;
 wire \A1/A2/A1/A1/M1/c1 ;
 wire \A1/A2/A1/A1/M1/c2 ;
 wire \A1/A2/A1/A1/M1/s1 ;
 wire \A1/A2/A1/A1/M2/c1 ;
 wire \A1/A2/A1/A1/M2/c2 ;
 wire \A1/A2/A1/A1/M2/s1 ;
 wire \A1/A2/A1/A1/M3/c1 ;
 wire \A1/A2/A1/A1/M3/c2 ;
 wire \A1/A2/A1/A1/M3/s1 ;
 wire \A1/A2/A1/A1/M4/c1 ;
 wire \A1/A2/A1/A1/M4/c2 ;
 wire \A1/A2/A1/A1/M4/s1 ;
 wire \A1/A2/A1/A2/c1 ;
 wire \A1/A2/A1/A2/c2 ;
 wire \A1/A2/A1/A2/c3 ;
 wire \A1/A2/A1/A2/M1/c1 ;
 wire \A1/A2/A1/A2/M1/c2 ;
 wire \A1/A2/A1/A2/M1/s1 ;
 wire \A1/A2/A1/A2/M2/c1 ;
 wire \A1/A2/A1/A2/M2/c2 ;
 wire \A1/A2/A1/A2/M2/s1 ;
 wire \A1/A2/A1/A2/M3/c1 ;
 wire \A1/A2/A1/A2/M3/c2 ;
 wire \A1/A2/A1/A2/M3/s1 ;
 wire \A1/A2/A1/A2/M4/c1 ;
 wire \A1/A2/A1/A2/M4/c2 ;
 wire \A1/A2/A1/A2/M4/s1 ;
 wire \A1/A2/A2/c1 ;
 wire \A1/A2/A2/A1/c1 ;
 wire \A1/A2/A2/A1/c2 ;
 wire \A1/A2/A2/A1/c3 ;
 wire \A1/A2/A2/A1/M1/c1 ;
 wire \A1/A2/A2/A1/M1/c2 ;
 wire \A1/A2/A2/A1/M1/s1 ;
 wire \A1/A2/A2/A1/M2/c1 ;
 wire \A1/A2/A2/A1/M2/c2 ;
 wire \A1/A2/A2/A1/M2/s1 ;
 wire \A1/A2/A2/A1/M3/c1 ;
 wire \A1/A2/A2/A1/M3/c2 ;
 wire \A1/A2/A2/A1/M3/s1 ;
 wire \A1/A2/A2/A1/M4/c1 ;
 wire \A1/A2/A2/A1/M4/c2 ;
 wire \A1/A2/A2/A1/M4/s1 ;
 wire \A1/A2/A2/A2/c1 ;
 wire \A1/A2/A2/A2/c2 ;
 wire \A1/A2/A2/A2/c3 ;
 wire \A1/A2/A2/A2/M1/c1 ;
 wire \A1/A2/A2/A2/M1/c2 ;
 wire \A1/A2/A2/A2/M1/s1 ;
 wire \A1/A2/A2/A2/M2/c1 ;
 wire \A1/A2/A2/A2/M2/c2 ;
 wire \A1/A2/A2/A2/M2/s1 ;
 wire \A1/A2/A2/A2/M3/c1 ;
 wire \A1/A2/A2/A2/M3/c2 ;
 wire \A1/A2/A2/A2/M3/s1 ;
 wire \A1/A2/A2/A2/M4/c1 ;
 wire \A1/A2/A2/A2/M4/c2 ;
 wire \A1/A2/A2/A2/M4/s1 ;
 wire \A2/c1 ;
 wire \A2/A1/c1 ;
 wire \A2/A1/A1/c1 ;
 wire \A2/A1/A1/A1/c1 ;
 wire \A2/A1/A1/A1/c2 ;
 wire \A2/A1/A1/A1/c3 ;
 wire \A2/A1/A1/A1/M1/c1 ;
 wire \A2/A1/A1/A1/M1/c2 ;
 wire \A2/A1/A1/A1/M1/s1 ;
 wire \A2/A1/A1/A1/M2/c1 ;
 wire \A2/A1/A1/A1/M2/c2 ;
 wire \A2/A1/A1/A1/M2/s1 ;
 wire \A2/A1/A1/A1/M3/c1 ;
 wire \A2/A1/A1/A1/M3/c2 ;
 wire \A2/A1/A1/A1/M3/s1 ;
 wire \A2/A1/A1/A1/M4/c1 ;
 wire \A2/A1/A1/A1/M4/c2 ;
 wire \A2/A1/A1/A1/M4/s1 ;
 wire \A2/A1/A1/A2/c1 ;
 wire \A2/A1/A1/A2/c2 ;
 wire \A2/A1/A1/A2/c3 ;
 wire \A2/A1/A1/A2/M1/c1 ;
 wire \A2/A1/A1/A2/M1/c2 ;
 wire \A2/A1/A1/A2/M1/s1 ;
 wire \A2/A1/A1/A2/M2/c1 ;
 wire \A2/A1/A1/A2/M2/c2 ;
 wire \A2/A1/A1/A2/M2/s1 ;
 wire \A2/A1/A1/A2/M3/c1 ;
 wire \A2/A1/A1/A2/M3/c2 ;
 wire \A2/A1/A1/A2/M3/s1 ;
 wire \A2/A1/A1/A2/M4/c1 ;
 wire \A2/A1/A1/A2/M4/c2 ;
 wire \A2/A1/A1/A2/M4/s1 ;
 wire \A2/A1/A2/c1 ;
 wire \A2/A1/A2/A1/c1 ;
 wire \A2/A1/A2/A1/c2 ;
 wire \A2/A1/A2/A1/c3 ;
 wire \A2/A1/A2/A1/M1/c1 ;
 wire \A2/A1/A2/A1/M1/c2 ;
 wire \A2/A1/A2/A1/M1/s1 ;
 wire \A2/A1/A2/A1/M2/c1 ;
 wire \A2/A1/A2/A1/M2/c2 ;
 wire \A2/A1/A2/A1/M2/s1 ;
 wire \A2/A1/A2/A1/M3/c1 ;
 wire \A2/A1/A2/A1/M3/c2 ;
 wire \A2/A1/A2/A1/M3/s1 ;
 wire \A2/A1/A2/A1/M4/c1 ;
 wire \A2/A1/A2/A1/M4/c2 ;
 wire \A2/A1/A2/A1/M4/s1 ;
 wire \A2/A1/A2/A2/c1 ;
 wire \A2/A1/A2/A2/c2 ;
 wire \A2/A1/A2/A2/c3 ;
 wire \A2/A1/A2/A2/M1/c1 ;
 wire \A2/A1/A2/A2/M1/c2 ;
 wire \A2/A1/A2/A2/M1/s1 ;
 wire \A2/A1/A2/A2/M2/c1 ;
 wire \A2/A1/A2/A2/M2/c2 ;
 wire \A2/A1/A2/A2/M2/s1 ;
 wire \A2/A1/A2/A2/M3/c1 ;
 wire \A2/A1/A2/A2/M3/c2 ;
 wire \A2/A1/A2/A2/M3/s1 ;
 wire \A2/A1/A2/A2/M4/c1 ;
 wire \A2/A1/A2/A2/M4/c2 ;
 wire \A2/A1/A2/A2/M4/s1 ;
 wire \A2/A2/c1 ;
 wire \A2/A2/A1/c1 ;
 wire \A2/A2/A1/A1/c1 ;
 wire \A2/A2/A1/A1/c2 ;
 wire \A2/A2/A1/A1/c3 ;
 wire \A2/A2/A1/A1/M1/c1 ;
 wire \A2/A2/A1/A1/M1/c2 ;
 wire \A2/A2/A1/A1/M1/s1 ;
 wire \A2/A2/A1/A1/M2/c1 ;
 wire \A2/A2/A1/A1/M2/c2 ;
 wire \A2/A2/A1/A1/M2/s1 ;
 wire \A2/A2/A1/A1/M3/c1 ;
 wire \A2/A2/A1/A1/M3/c2 ;
 wire \A2/A2/A1/A1/M3/s1 ;
 wire \A2/A2/A1/A1/M4/c1 ;
 wire \A2/A2/A1/A1/M4/c2 ;
 wire \A2/A2/A1/A1/M4/s1 ;
 wire \A2/A2/A1/A2/c1 ;
 wire \A2/A2/A1/A2/c2 ;
 wire \A2/A2/A1/A2/c3 ;
 wire \A2/A2/A1/A2/M1/c1 ;
 wire \A2/A2/A1/A2/M1/c2 ;
 wire \A2/A2/A1/A2/M1/s1 ;
 wire \A2/A2/A1/A2/M2/c1 ;
 wire \A2/A2/A1/A2/M2/c2 ;
 wire \A2/A2/A1/A2/M2/s1 ;
 wire \A2/A2/A1/A2/M3/c1 ;
 wire \A2/A2/A1/A2/M3/c2 ;
 wire \A2/A2/A1/A2/M3/s1 ;
 wire \A2/A2/A1/A2/M4/c1 ;
 wire \A2/A2/A1/A2/M4/c2 ;
 wire \A2/A2/A1/A2/M4/s1 ;
 wire \A2/A2/A2/c1 ;
 wire \A2/A2/A2/A1/c1 ;
 wire \A2/A2/A2/A1/c2 ;
 wire \A2/A2/A2/A1/c3 ;
 wire \A2/A2/A2/A1/M1/c1 ;
 wire \A2/A2/A2/A1/M1/c2 ;
 wire \A2/A2/A2/A1/M1/s1 ;
 wire \A2/A2/A2/A1/M2/c1 ;
 wire \A2/A2/A2/A1/M2/c2 ;
 wire \A2/A2/A2/A1/M2/s1 ;
 wire \A2/A2/A2/A1/M3/c1 ;
 wire \A2/A2/A2/A1/M3/c2 ;
 wire \A2/A2/A2/A1/M3/s1 ;
 wire \A2/A2/A2/A1/M4/c1 ;
 wire \A2/A2/A2/A1/M4/c2 ;
 wire \A2/A2/A2/A1/M4/s1 ;
 wire \A2/A2/A2/A2/c1 ;
 wire \A2/A2/A2/A2/c2 ;
 wire \A2/A2/A2/A2/c3 ;
 wire \A2/A2/A2/A2/M1/c1 ;
 wire \A2/A2/A2/A2/M1/c2 ;
 wire \A2/A2/A2/A2/M1/s1 ;
 wire \A2/A2/A2/A2/M2/c1 ;
 wire \A2/A2/A2/A2/M2/c2 ;
 wire \A2/A2/A2/A2/M2/s1 ;
 wire \A2/A2/A2/A2/M3/c1 ;
 wire \A2/A2/A2/A2/M3/c2 ;
 wire \A2/A2/A2/A2/M3/s1 ;
 wire \A2/A2/A2/A2/M4/c1 ;
 wire \A2/A2/A2/A2/M4/c2 ;
 wire \A2/A2/A2/A2/M4/s1 ;
 wire \A3/c1 ;
 wire \A3/A1/c1 ;
 wire \A3/A1/A1/c1 ;
 wire \A3/A1/A1/A1/c1 ;
 wire \A3/A1/A1/A1/c2 ;
 wire \A3/A1/A1/A1/c3 ;
 wire \A3/A1/A1/A1/M1/c1 ;
 wire \A3/A1/A1/A1/M1/c2 ;
 wire \A3/A1/A1/A1/M1/s1 ;
 wire \A3/A1/A1/A1/M2/c1 ;
 wire \A3/A1/A1/A1/M2/c2 ;
 wire \A3/A1/A1/A1/M2/s1 ;
 wire \A3/A1/A1/A1/M3/c1 ;
 wire \A3/A1/A1/A1/M3/c2 ;
 wire \A3/A1/A1/A1/M3/s1 ;
 wire \A3/A1/A1/A1/M4/c1 ;
 wire \A3/A1/A1/A1/M4/c2 ;
 wire \A3/A1/A1/A1/M4/s1 ;
 wire \A3/A1/A1/A2/c1 ;
 wire \A3/A1/A1/A2/c2 ;
 wire \A3/A1/A1/A2/c3 ;
 wire \A3/A1/A1/A2/M1/c1 ;
 wire \A3/A1/A1/A2/M1/c2 ;
 wire \A3/A1/A1/A2/M1/s1 ;
 wire \A3/A1/A1/A2/M2/c1 ;
 wire \A3/A1/A1/A2/M2/c2 ;
 wire \A3/A1/A1/A2/M2/s1 ;
 wire \A3/A1/A1/A2/M3/c1 ;
 wire \A3/A1/A1/A2/M3/c2 ;
 wire \A3/A1/A1/A2/M3/s1 ;
 wire \A3/A1/A1/A2/M4/c1 ;
 wire \A3/A1/A1/A2/M4/c2 ;
 wire \A3/A1/A1/A2/M4/s1 ;
 wire \A3/A1/A2/c1 ;
 wire \A3/A1/A2/A1/c1 ;
 wire \A3/A1/A2/A1/c2 ;
 wire \A3/A1/A2/A1/c3 ;
 wire \A3/A1/A2/A1/M1/c1 ;
 wire \A3/A1/A2/A1/M1/c2 ;
 wire \A3/A1/A2/A1/M1/s1 ;
 wire \A3/A1/A2/A1/M2/c1 ;
 wire \A3/A1/A2/A1/M2/c2 ;
 wire \A3/A1/A2/A1/M2/s1 ;
 wire \A3/A1/A2/A1/M3/c1 ;
 wire \A3/A1/A2/A1/M3/c2 ;
 wire \A3/A1/A2/A1/M3/s1 ;
 wire \A3/A1/A2/A1/M4/c1 ;
 wire \A3/A1/A2/A1/M4/c2 ;
 wire \A3/A1/A2/A1/M4/s1 ;
 wire \A3/A1/A2/A2/c1 ;
 wire \A3/A1/A2/A2/c2 ;
 wire \A3/A1/A2/A2/c3 ;
 wire \A3/A1/A2/A2/M1/c1 ;
 wire \A3/A1/A2/A2/M1/c2 ;
 wire \A3/A1/A2/A2/M1/s1 ;
 wire \A3/A1/A2/A2/M2/c1 ;
 wire \A3/A1/A2/A2/M2/c2 ;
 wire \A3/A1/A2/A2/M2/s1 ;
 wire \A3/A1/A2/A2/M3/c1 ;
 wire \A3/A1/A2/A2/M3/c2 ;
 wire \A3/A1/A2/A2/M3/s1 ;
 wire \A3/A1/A2/A2/M4/c1 ;
 wire \A3/A1/A2/A2/M4/c2 ;
 wire \A3/A1/A2/A2/M4/s1 ;
 wire \A3/A2/c1 ;
 wire \A3/A2/A1/c1 ;
 wire \A3/A2/A1/A1/c1 ;
 wire \A3/A2/A1/A1/c2 ;
 wire \A3/A2/A1/A1/c3 ;
 wire \A3/A2/A1/A1/M1/c1 ;
 wire \A3/A2/A1/A1/M1/c2 ;
 wire \A3/A2/A1/A1/M1/s1 ;
 wire \A3/A2/A1/A1/M2/c1 ;
 wire \A3/A2/A1/A1/M2/c2 ;
 wire \A3/A2/A1/A1/M2/s1 ;
 wire \A3/A2/A1/A1/M3/c1 ;
 wire \A3/A2/A1/A1/M3/c2 ;
 wire \A3/A2/A1/A1/M3/s1 ;
 wire \A3/A2/A1/A1/M4/c1 ;
 wire \A3/A2/A1/A1/M4/c2 ;
 wire \A3/A2/A1/A1/M4/s1 ;
 wire \A3/A2/A1/A2/c1 ;
 wire \A3/A2/A1/A2/c2 ;
 wire \A3/A2/A1/A2/c3 ;
 wire \A3/A2/A1/A2/M1/c1 ;
 wire \A3/A2/A1/A2/M1/c2 ;
 wire \A3/A2/A1/A2/M1/s1 ;
 wire \A3/A2/A1/A2/M2/c1 ;
 wire \A3/A2/A1/A2/M2/c2 ;
 wire \A3/A2/A1/A2/M2/s1 ;
 wire \A3/A2/A1/A2/M3/c1 ;
 wire \A3/A2/A1/A2/M3/c2 ;
 wire \A3/A2/A1/A2/M3/s1 ;
 wire \A3/A2/A1/A2/M4/c1 ;
 wire \A3/A2/A1/A2/M4/c2 ;
 wire \A3/A2/A1/A2/M4/s1 ;
 wire \A3/A2/A2/c1 ;
 wire \A3/A2/A2/A1/c1 ;
 wire \A3/A2/A2/A1/c2 ;
 wire \A3/A2/A2/A1/c3 ;
 wire \A3/A2/A2/A1/M1/c1 ;
 wire \A3/A2/A2/A1/M1/c2 ;
 wire \A3/A2/A2/A1/M1/s1 ;
 wire \A3/A2/A2/A1/M2/c1 ;
 wire \A3/A2/A2/A1/M2/c2 ;
 wire \A3/A2/A2/A1/M2/s1 ;
 wire \A3/A2/A2/A1/M3/c1 ;
 wire \A3/A2/A2/A1/M3/c2 ;
 wire \A3/A2/A2/A1/M3/s1 ;
 wire \A3/A2/A2/A1/M4/c1 ;
 wire \A3/A2/A2/A1/M4/c2 ;
 wire \A3/A2/A2/A1/M4/s1 ;
 wire \A3/A2/A2/A2/c1 ;
 wire \A3/A2/A2/A2/c2 ;
 wire \A3/A2/A2/A2/c3 ;
 wire \A3/A2/A2/A2/M1/c1 ;
 wire \A3/A2/A2/A2/M1/c2 ;
 wire \A3/A2/A2/A2/M1/s1 ;
 wire \A3/A2/A2/A2/M2/c1 ;
 wire \A3/A2/A2/A2/M2/c2 ;
 wire \A3/A2/A2/A2/M2/s1 ;
 wire \A3/A2/A2/A2/M3/c1 ;
 wire \A3/A2/A2/A2/M3/c2 ;
 wire \A3/A2/A2/A2/M3/s1 ;
 wire \A3/A2/A2/A2/M4/c1 ;
 wire \A3/A2/A2/A2/M4/c2 ;
 wire \A3/A2/A2/A2/M4/s1 ;
 wire \V1/c1 ;
 wire \V1/c2 ;
 wire \V1/c3 ;
 wire \V1/overflow ;
 wire \V1/A1/c1 ;
 wire \V1/A1/A1/c1 ;
 wire \V1/A1/A1/A1/c1 ;
 wire \V1/A1/A1/A1/c2 ;
 wire \V1/A1/A1/A1/c3 ;
 wire \V1/A1/A1/A1/M1/c1 ;
 wire \V1/A1/A1/A1/M1/c2 ;
 wire \V1/A1/A1/A1/M1/s1 ;
 wire \V1/A1/A1/A1/M2/c1 ;
 wire \V1/A1/A1/A1/M2/c2 ;
 wire \V1/A1/A1/A1/M2/s1 ;
 wire \V1/A1/A1/A1/M3/c1 ;
 wire \V1/A1/A1/A1/M3/c2 ;
 wire \V1/A1/A1/A1/M3/s1 ;
 wire \V1/A1/A1/A1/M4/c1 ;
 wire \V1/A1/A1/A1/M4/c2 ;
 wire \V1/A1/A1/A1/M4/s1 ;
 wire \V1/A1/A1/A2/c1 ;
 wire \V1/A1/A1/A2/c2 ;
 wire \V1/A1/A1/A2/c3 ;
 wire \V1/A1/A1/A2/M1/c1 ;
 wire \V1/A1/A1/A2/M1/c2 ;
 wire \V1/A1/A1/A2/M1/s1 ;
 wire \V1/A1/A1/A2/M2/c1 ;
 wire \V1/A1/A1/A2/M2/c2 ;
 wire \V1/A1/A1/A2/M2/s1 ;
 wire \V1/A1/A1/A2/M3/c1 ;
 wire \V1/A1/A1/A2/M3/c2 ;
 wire \V1/A1/A1/A2/M3/s1 ;
 wire \V1/A1/A1/A2/M4/c1 ;
 wire \V1/A1/A1/A2/M4/c2 ;
 wire \V1/A1/A1/A2/M4/s1 ;
 wire \V1/A1/A2/c1 ;
 wire \V1/A1/A2/A1/c1 ;
 wire \V1/A1/A2/A1/c2 ;
 wire \V1/A1/A2/A1/c3 ;
 wire \V1/A1/A2/A1/M1/c1 ;
 wire \V1/A1/A2/A1/M1/c2 ;
 wire \V1/A1/A2/A1/M1/s1 ;
 wire \V1/A1/A2/A1/M2/c1 ;
 wire \V1/A1/A2/A1/M2/c2 ;
 wire \V1/A1/A2/A1/M2/s1 ;
 wire \V1/A1/A2/A1/M3/c1 ;
 wire \V1/A1/A2/A1/M3/c2 ;
 wire \V1/A1/A2/A1/M3/s1 ;
 wire \V1/A1/A2/A1/M4/c1 ;
 wire \V1/A1/A2/A1/M4/c2 ;
 wire \V1/A1/A2/A1/M4/s1 ;
 wire \V1/A1/A2/A2/c1 ;
 wire \V1/A1/A2/A2/c2 ;
 wire \V1/A1/A2/A2/c3 ;
 wire \V1/A1/A2/A2/M1/c1 ;
 wire \V1/A1/A2/A2/M1/c2 ;
 wire \V1/A1/A2/A2/M1/s1 ;
 wire \V1/A1/A2/A2/M2/c1 ;
 wire \V1/A1/A2/A2/M2/c2 ;
 wire \V1/A1/A2/A2/M2/s1 ;
 wire \V1/A1/A2/A2/M3/c1 ;
 wire \V1/A1/A2/A2/M3/c2 ;
 wire \V1/A1/A2/A2/M3/s1 ;
 wire \V1/A1/A2/A2/M4/c1 ;
 wire \V1/A1/A2/A2/M4/c2 ;
 wire \V1/A1/A2/A2/M4/s1 ;
 wire \V1/A2/c1 ;
 wire \V1/A2/A1/c1 ;
 wire \V1/A2/A1/A1/c1 ;
 wire \V1/A2/A1/A1/c2 ;
 wire \V1/A2/A1/A1/c3 ;
 wire \V1/A2/A1/A1/M1/c1 ;
 wire \V1/A2/A1/A1/M1/c2 ;
 wire \V1/A2/A1/A1/M1/s1 ;
 wire \V1/A2/A1/A1/M2/c1 ;
 wire \V1/A2/A1/A1/M2/c2 ;
 wire \V1/A2/A1/A1/M2/s1 ;
 wire \V1/A2/A1/A1/M3/c1 ;
 wire \V1/A2/A1/A1/M3/c2 ;
 wire \V1/A2/A1/A1/M3/s1 ;
 wire \V1/A2/A1/A1/M4/c1 ;
 wire \V1/A2/A1/A1/M4/c2 ;
 wire \V1/A2/A1/A1/M4/s1 ;
 wire \V1/A2/A1/A2/c1 ;
 wire \V1/A2/A1/A2/c2 ;
 wire \V1/A2/A1/A2/c3 ;
 wire \V1/A2/A1/A2/M1/c1 ;
 wire \V1/A2/A1/A2/M1/c2 ;
 wire \V1/A2/A1/A2/M1/s1 ;
 wire \V1/A2/A1/A2/M2/c1 ;
 wire \V1/A2/A1/A2/M2/c2 ;
 wire \V1/A2/A1/A2/M2/s1 ;
 wire \V1/A2/A1/A2/M3/c1 ;
 wire \V1/A2/A1/A2/M3/c2 ;
 wire \V1/A2/A1/A2/M3/s1 ;
 wire \V1/A2/A1/A2/M4/c1 ;
 wire \V1/A2/A1/A2/M4/c2 ;
 wire \V1/A2/A1/A2/M4/s1 ;
 wire \V1/A2/A2/c1 ;
 wire \V1/A2/A2/A1/c1 ;
 wire \V1/A2/A2/A1/c2 ;
 wire \V1/A2/A2/A1/c3 ;
 wire \V1/A2/A2/A1/M1/c1 ;
 wire \V1/A2/A2/A1/M1/c2 ;
 wire \V1/A2/A2/A1/M1/s1 ;
 wire \V1/A2/A2/A1/M2/c1 ;
 wire \V1/A2/A2/A1/M2/c2 ;
 wire \V1/A2/A2/A1/M2/s1 ;
 wire \V1/A2/A2/A1/M3/c1 ;
 wire \V1/A2/A2/A1/M3/c2 ;
 wire \V1/A2/A2/A1/M3/s1 ;
 wire \V1/A2/A2/A1/M4/c1 ;
 wire \V1/A2/A2/A1/M4/c2 ;
 wire \V1/A2/A2/A1/M4/s1 ;
 wire \V1/A2/A2/A2/c1 ;
 wire \V1/A2/A2/A2/c2 ;
 wire \V1/A2/A2/A2/c3 ;
 wire \V1/A2/A2/A2/M1/c1 ;
 wire \V1/A2/A2/A2/M1/c2 ;
 wire \V1/A2/A2/A2/M1/s1 ;
 wire \V1/A2/A2/A2/M2/c1 ;
 wire \V1/A2/A2/A2/M2/c2 ;
 wire \V1/A2/A2/A2/M2/s1 ;
 wire \V1/A2/A2/A2/M3/c1 ;
 wire \V1/A2/A2/A2/M3/c2 ;
 wire \V1/A2/A2/A2/M3/s1 ;
 wire \V1/A2/A2/A2/M4/c1 ;
 wire \V1/A2/A2/A2/M4/c2 ;
 wire \V1/A2/A2/A2/M4/s1 ;
 wire \V1/A3/c1 ;
 wire \V1/A3/A1/c1 ;
 wire \V1/A3/A1/A1/c1 ;
 wire \V1/A3/A1/A1/c2 ;
 wire \V1/A3/A1/A1/c3 ;
 wire \V1/A3/A1/A1/M1/c1 ;
 wire \V1/A3/A1/A1/M1/c2 ;
 wire \V1/A3/A1/A1/M1/s1 ;
 wire \V1/A3/A1/A1/M2/c1 ;
 wire \V1/A3/A1/A1/M2/c2 ;
 wire \V1/A3/A1/A1/M2/s1 ;
 wire \V1/A3/A1/A1/M3/c1 ;
 wire \V1/A3/A1/A1/M3/c2 ;
 wire \V1/A3/A1/A1/M3/s1 ;
 wire \V1/A3/A1/A1/M4/c1 ;
 wire \V1/A3/A1/A1/M4/c2 ;
 wire \V1/A3/A1/A1/M4/s1 ;
 wire \V1/A3/A1/A2/c1 ;
 wire \V1/A3/A1/A2/c2 ;
 wire \V1/A3/A1/A2/c3 ;
 wire \V1/A3/A1/A2/M1/c1 ;
 wire \V1/A3/A1/A2/M1/c2 ;
 wire \V1/A3/A1/A2/M1/s1 ;
 wire \V1/A3/A1/A2/M2/c1 ;
 wire \V1/A3/A1/A2/M2/c2 ;
 wire \V1/A3/A1/A2/M2/s1 ;
 wire \V1/A3/A1/A2/M3/c1 ;
 wire \V1/A3/A1/A2/M3/c2 ;
 wire \V1/A3/A1/A2/M3/s1 ;
 wire \V1/A3/A1/A2/M4/c1 ;
 wire \V1/A3/A1/A2/M4/c2 ;
 wire \V1/A3/A1/A2/M4/s1 ;
 wire \V1/A3/A2/c1 ;
 wire \V1/A3/A2/A1/c1 ;
 wire \V1/A3/A2/A1/c2 ;
 wire \V1/A3/A2/A1/c3 ;
 wire \V1/A3/A2/A1/M1/c1 ;
 wire \V1/A3/A2/A1/M1/c2 ;
 wire \V1/A3/A2/A1/M1/s1 ;
 wire \V1/A3/A2/A1/M2/c1 ;
 wire \V1/A3/A2/A1/M2/c2 ;
 wire \V1/A3/A2/A1/M2/s1 ;
 wire \V1/A3/A2/A1/M3/c1 ;
 wire \V1/A3/A2/A1/M3/c2 ;
 wire \V1/A3/A2/A1/M3/s1 ;
 wire \V1/A3/A2/A1/M4/c1 ;
 wire \V1/A3/A2/A1/M4/c2 ;
 wire \V1/A3/A2/A1/M4/s1 ;
 wire \V1/A3/A2/A2/c1 ;
 wire \V1/A3/A2/A2/c2 ;
 wire \V1/A3/A2/A2/c3 ;
 wire \V1/A3/A2/A2/M1/c1 ;
 wire \V1/A3/A2/A2/M1/c2 ;
 wire \V1/A3/A2/A2/M1/s1 ;
 wire \V1/A3/A2/A2/M2/c1 ;
 wire \V1/A3/A2/A2/M2/c2 ;
 wire \V1/A3/A2/A2/M2/s1 ;
 wire \V1/A3/A2/A2/M3/c1 ;
 wire \V1/A3/A2/A2/M3/c2 ;
 wire \V1/A3/A2/A2/M3/s1 ;
 wire \V1/A3/A2/A2/M4/c1 ;
 wire \V1/A3/A2/A2/M4/c2 ;
 wire \V1/A3/A2/A2/M4/s1 ;
 wire \V1/V1/c1 ;
 wire \V1/V1/c2 ;
 wire \V1/V1/c3 ;
 wire \V1/V1/overflow ;
 wire \V1/V1/A1/c1 ;
 wire \V1/V1/A1/A1/c1 ;
 wire \V1/V1/A1/A1/c2 ;
 wire \V1/V1/A1/A1/c3 ;
 wire \V1/V1/A1/A1/M1/c1 ;
 wire \V1/V1/A1/A1/M1/c2 ;
 wire \V1/V1/A1/A1/M1/s1 ;
 wire \V1/V1/A1/A1/M2/c1 ;
 wire \V1/V1/A1/A1/M2/c2 ;
 wire \V1/V1/A1/A1/M2/s1 ;
 wire \V1/V1/A1/A1/M3/c1 ;
 wire \V1/V1/A1/A1/M3/c2 ;
 wire \V1/V1/A1/A1/M3/s1 ;
 wire \V1/V1/A1/A1/M4/c1 ;
 wire \V1/V1/A1/A1/M4/c2 ;
 wire \V1/V1/A1/A1/M4/s1 ;
 wire \V1/V1/A1/A2/c1 ;
 wire \V1/V1/A1/A2/c2 ;
 wire \V1/V1/A1/A2/c3 ;
 wire \V1/V1/A1/A2/M1/c1 ;
 wire \V1/V1/A1/A2/M1/c2 ;
 wire \V1/V1/A1/A2/M1/s1 ;
 wire \V1/V1/A1/A2/M2/c1 ;
 wire \V1/V1/A1/A2/M2/c2 ;
 wire \V1/V1/A1/A2/M2/s1 ;
 wire \V1/V1/A1/A2/M3/c1 ;
 wire \V1/V1/A1/A2/M3/c2 ;
 wire \V1/V1/A1/A2/M3/s1 ;
 wire \V1/V1/A1/A2/M4/c1 ;
 wire \V1/V1/A1/A2/M4/c2 ;
 wire \V1/V1/A1/A2/M4/s1 ;
 wire \V1/V1/A2/c1 ;
 wire \V1/V1/A2/A1/c1 ;
 wire \V1/V1/A2/A1/c2 ;
 wire \V1/V1/A2/A1/c3 ;
 wire \V1/V1/A2/A1/M1/c1 ;
 wire \V1/V1/A2/A1/M1/c2 ;
 wire \V1/V1/A2/A1/M1/s1 ;
 wire \V1/V1/A2/A1/M2/c1 ;
 wire \V1/V1/A2/A1/M2/c2 ;
 wire \V1/V1/A2/A1/M2/s1 ;
 wire \V1/V1/A2/A1/M3/c1 ;
 wire \V1/V1/A2/A1/M3/c2 ;
 wire \V1/V1/A2/A1/M3/s1 ;
 wire \V1/V1/A2/A1/M4/c1 ;
 wire \V1/V1/A2/A1/M4/c2 ;
 wire \V1/V1/A2/A1/M4/s1 ;
 wire \V1/V1/A2/A2/c1 ;
 wire \V1/V1/A2/A2/c2 ;
 wire \V1/V1/A2/A2/c3 ;
 wire \V1/V1/A2/A2/M1/c1 ;
 wire \V1/V1/A2/A2/M1/c2 ;
 wire \V1/V1/A2/A2/M1/s1 ;
 wire \V1/V1/A2/A2/M2/c1 ;
 wire \V1/V1/A2/A2/M2/c2 ;
 wire \V1/V1/A2/A2/M2/s1 ;
 wire \V1/V1/A2/A2/M3/c1 ;
 wire \V1/V1/A2/A2/M3/c2 ;
 wire \V1/V1/A2/A2/M3/s1 ;
 wire \V1/V1/A2/A2/M4/c1 ;
 wire \V1/V1/A2/A2/M4/c2 ;
 wire \V1/V1/A2/A2/M4/s1 ;
 wire \V1/V1/A3/c1 ;
 wire \V1/V1/A3/A1/c1 ;
 wire \V1/V1/A3/A1/c2 ;
 wire \V1/V1/A3/A1/c3 ;
 wire \V1/V1/A3/A1/M1/c1 ;
 wire \V1/V1/A3/A1/M1/c2 ;
 wire \V1/V1/A3/A1/M1/s1 ;
 wire \V1/V1/A3/A1/M2/c1 ;
 wire \V1/V1/A3/A1/M2/c2 ;
 wire \V1/V1/A3/A1/M2/s1 ;
 wire \V1/V1/A3/A1/M3/c1 ;
 wire \V1/V1/A3/A1/M3/c2 ;
 wire \V1/V1/A3/A1/M3/s1 ;
 wire \V1/V1/A3/A1/M4/c1 ;
 wire \V1/V1/A3/A1/M4/c2 ;
 wire \V1/V1/A3/A1/M4/s1 ;
 wire \V1/V1/A3/A2/c1 ;
 wire \V1/V1/A3/A2/c2 ;
 wire \V1/V1/A3/A2/c3 ;
 wire \V1/V1/A3/A2/M1/c1 ;
 wire \V1/V1/A3/A2/M1/c2 ;
 wire \V1/V1/A3/A2/M1/s1 ;
 wire \V1/V1/A3/A2/M2/c1 ;
 wire \V1/V1/A3/A2/M2/c2 ;
 wire \V1/V1/A3/A2/M2/s1 ;
 wire \V1/V1/A3/A2/M3/c1 ;
 wire \V1/V1/A3/A2/M3/c2 ;
 wire \V1/V1/A3/A2/M3/s1 ;
 wire \V1/V1/A3/A2/M4/c1 ;
 wire \V1/V1/A3/A2/M4/c2 ;
 wire \V1/V1/A3/A2/M4/s1 ;
 wire \V1/V1/V1/c1 ;
 wire \V1/V1/V1/c2 ;
 wire \V1/V1/V1/c3 ;
 wire \V1/V1/V1/overflow ;
 wire \V1/V1/V1/A1/c1 ;
 wire \V1/V1/V1/A1/c2 ;
 wire \V1/V1/V1/A1/c3 ;
 wire \V1/V1/V1/A1/M1/c1 ;
 wire \V1/V1/V1/A1/M1/c2 ;
 wire \V1/V1/V1/A1/M1/s1 ;
 wire \V1/V1/V1/A1/M2/c1 ;
 wire \V1/V1/V1/A1/M2/c2 ;
 wire \V1/V1/V1/A1/M2/s1 ;
 wire \V1/V1/V1/A1/M3/c1 ;
 wire \V1/V1/V1/A1/M3/c2 ;
 wire \V1/V1/V1/A1/M3/s1 ;
 wire \V1/V1/V1/A1/M4/c1 ;
 wire \V1/V1/V1/A1/M4/c2 ;
 wire \V1/V1/V1/A1/M4/s1 ;
 wire \V1/V1/V1/A2/c1 ;
 wire \V1/V1/V1/A2/c2 ;
 wire \V1/V1/V1/A2/c3 ;
 wire \V1/V1/V1/A2/M1/c1 ;
 wire \V1/V1/V1/A2/M1/c2 ;
 wire \V1/V1/V1/A2/M1/s1 ;
 wire \V1/V1/V1/A2/M2/c1 ;
 wire \V1/V1/V1/A2/M2/c2 ;
 wire \V1/V1/V1/A2/M2/s1 ;
 wire \V1/V1/V1/A2/M3/c1 ;
 wire \V1/V1/V1/A2/M3/c2 ;
 wire \V1/V1/V1/A2/M3/s1 ;
 wire \V1/V1/V1/A2/M4/c1 ;
 wire \V1/V1/V1/A2/M4/c2 ;
 wire \V1/V1/V1/A2/M4/s1 ;
 wire \V1/V1/V1/A3/c1 ;
 wire \V1/V1/V1/A3/c2 ;
 wire \V1/V1/V1/A3/c3 ;
 wire \V1/V1/V1/A3/M1/c1 ;
 wire \V1/V1/V1/A3/M1/c2 ;
 wire \V1/V1/V1/A3/M1/s1 ;
 wire \V1/V1/V1/A3/M2/c1 ;
 wire \V1/V1/V1/A3/M2/c2 ;
 wire \V1/V1/V1/A3/M2/s1 ;
 wire \V1/V1/V1/A3/M3/c1 ;
 wire \V1/V1/V1/A3/M3/c2 ;
 wire \V1/V1/V1/A3/M3/s1 ;
 wire \V1/V1/V1/A3/M4/c1 ;
 wire \V1/V1/V1/A3/M4/c2 ;
 wire \V1/V1/V1/A3/M4/s1 ;
 wire \V1/V1/V1/V1/w1 ;
 wire \V1/V1/V1/V1/w2 ;
 wire \V1/V1/V1/V1/w3 ;
 wire \V1/V1/V1/V1/w4 ;
 wire \V1/V1/V1/V2/w1 ;
 wire \V1/V1/V1/V2/w2 ;
 wire \V1/V1/V1/V2/w3 ;
 wire \V1/V1/V1/V2/w4 ;
 wire \V1/V1/V1/V3/w1 ;
 wire \V1/V1/V1/V3/w2 ;
 wire \V1/V1/V1/V3/w3 ;
 wire \V1/V1/V1/V3/w4 ;
 wire \V1/V1/V1/V4/w1 ;
 wire \V1/V1/V1/V4/w2 ;
 wire \V1/V1/V1/V4/w3 ;
 wire \V1/V1/V1/V4/w4 ;
 wire \V1/V1/V2/c1 ;
 wire \V1/V1/V2/c2 ;
 wire \V1/V1/V2/c3 ;
 wire \V1/V1/V2/overflow ;
 wire \V1/V1/V2/A1/c1 ;
 wire \V1/V1/V2/A1/c2 ;
 wire \V1/V1/V2/A1/c3 ;
 wire \V1/V1/V2/A1/M1/c1 ;
 wire \V1/V1/V2/A1/M1/c2 ;
 wire \V1/V1/V2/A1/M1/s1 ;
 wire \V1/V1/V2/A1/M2/c1 ;
 wire \V1/V1/V2/A1/M2/c2 ;
 wire \V1/V1/V2/A1/M2/s1 ;
 wire \V1/V1/V2/A1/M3/c1 ;
 wire \V1/V1/V2/A1/M3/c2 ;
 wire \V1/V1/V2/A1/M3/s1 ;
 wire \V1/V1/V2/A1/M4/c1 ;
 wire \V1/V1/V2/A1/M4/c2 ;
 wire \V1/V1/V2/A1/M4/s1 ;
 wire \V1/V1/V2/A2/c1 ;
 wire \V1/V1/V2/A2/c2 ;
 wire \V1/V1/V2/A2/c3 ;
 wire \V1/V1/V2/A2/M1/c1 ;
 wire \V1/V1/V2/A2/M1/c2 ;
 wire \V1/V1/V2/A2/M1/s1 ;
 wire \V1/V1/V2/A2/M2/c1 ;
 wire \V1/V1/V2/A2/M2/c2 ;
 wire \V1/V1/V2/A2/M2/s1 ;
 wire \V1/V1/V2/A2/M3/c1 ;
 wire \V1/V1/V2/A2/M3/c2 ;
 wire \V1/V1/V2/A2/M3/s1 ;
 wire \V1/V1/V2/A2/M4/c1 ;
 wire \V1/V1/V2/A2/M4/c2 ;
 wire \V1/V1/V2/A2/M4/s1 ;
 wire \V1/V1/V2/A3/c1 ;
 wire \V1/V1/V2/A3/c2 ;
 wire \V1/V1/V2/A3/c3 ;
 wire \V1/V1/V2/A3/M1/c1 ;
 wire \V1/V1/V2/A3/M1/c2 ;
 wire \V1/V1/V2/A3/M1/s1 ;
 wire \V1/V1/V2/A3/M2/c1 ;
 wire \V1/V1/V2/A3/M2/c2 ;
 wire \V1/V1/V2/A3/M2/s1 ;
 wire \V1/V1/V2/A3/M3/c1 ;
 wire \V1/V1/V2/A3/M3/c2 ;
 wire \V1/V1/V2/A3/M3/s1 ;
 wire \V1/V1/V2/A3/M4/c1 ;
 wire \V1/V1/V2/A3/M4/c2 ;
 wire \V1/V1/V2/A3/M4/s1 ;
 wire \V1/V1/V2/V1/w1 ;
 wire \V1/V1/V2/V1/w2 ;
 wire \V1/V1/V2/V1/w3 ;
 wire \V1/V1/V2/V1/w4 ;
 wire \V1/V1/V2/V2/w1 ;
 wire \V1/V1/V2/V2/w2 ;
 wire \V1/V1/V2/V2/w3 ;
 wire \V1/V1/V2/V2/w4 ;
 wire \V1/V1/V2/V3/w1 ;
 wire \V1/V1/V2/V3/w2 ;
 wire \V1/V1/V2/V3/w3 ;
 wire \V1/V1/V2/V3/w4 ;
 wire \V1/V1/V2/V4/w1 ;
 wire \V1/V1/V2/V4/w2 ;
 wire \V1/V1/V2/V4/w3 ;
 wire \V1/V1/V2/V4/w4 ;
 wire \V1/V1/V3/c1 ;
 wire \V1/V1/V3/c2 ;
 wire \V1/V1/V3/c3 ;
 wire \V1/V1/V3/overflow ;
 wire \V1/V1/V3/A1/c1 ;
 wire \V1/V1/V3/A1/c2 ;
 wire \V1/V1/V3/A1/c3 ;
 wire \V1/V1/V3/A1/M1/c1 ;
 wire \V1/V1/V3/A1/M1/c2 ;
 wire \V1/V1/V3/A1/M1/s1 ;
 wire \V1/V1/V3/A1/M2/c1 ;
 wire \V1/V1/V3/A1/M2/c2 ;
 wire \V1/V1/V3/A1/M2/s1 ;
 wire \V1/V1/V3/A1/M3/c1 ;
 wire \V1/V1/V3/A1/M3/c2 ;
 wire \V1/V1/V3/A1/M3/s1 ;
 wire \V1/V1/V3/A1/M4/c1 ;
 wire \V1/V1/V3/A1/M4/c2 ;
 wire \V1/V1/V3/A1/M4/s1 ;
 wire \V1/V1/V3/A2/c1 ;
 wire \V1/V1/V3/A2/c2 ;
 wire \V1/V1/V3/A2/c3 ;
 wire \V1/V1/V3/A2/M1/c1 ;
 wire \V1/V1/V3/A2/M1/c2 ;
 wire \V1/V1/V3/A2/M1/s1 ;
 wire \V1/V1/V3/A2/M2/c1 ;
 wire \V1/V1/V3/A2/M2/c2 ;
 wire \V1/V1/V3/A2/M2/s1 ;
 wire \V1/V1/V3/A2/M3/c1 ;
 wire \V1/V1/V3/A2/M3/c2 ;
 wire \V1/V1/V3/A2/M3/s1 ;
 wire \V1/V1/V3/A2/M4/c1 ;
 wire \V1/V1/V3/A2/M4/c2 ;
 wire \V1/V1/V3/A2/M4/s1 ;
 wire \V1/V1/V3/A3/c1 ;
 wire \V1/V1/V3/A3/c2 ;
 wire \V1/V1/V3/A3/c3 ;
 wire \V1/V1/V3/A3/M1/c1 ;
 wire \V1/V1/V3/A3/M1/c2 ;
 wire \V1/V1/V3/A3/M1/s1 ;
 wire \V1/V1/V3/A3/M2/c1 ;
 wire \V1/V1/V3/A3/M2/c2 ;
 wire \V1/V1/V3/A3/M2/s1 ;
 wire \V1/V1/V3/A3/M3/c1 ;
 wire \V1/V1/V3/A3/M3/c2 ;
 wire \V1/V1/V3/A3/M3/s1 ;
 wire \V1/V1/V3/A3/M4/c1 ;
 wire \V1/V1/V3/A3/M4/c2 ;
 wire \V1/V1/V3/A3/M4/s1 ;
 wire \V1/V1/V3/V1/w1 ;
 wire \V1/V1/V3/V1/w2 ;
 wire \V1/V1/V3/V1/w3 ;
 wire \V1/V1/V3/V1/w4 ;
 wire \V1/V1/V3/V2/w1 ;
 wire \V1/V1/V3/V2/w2 ;
 wire \V1/V1/V3/V2/w3 ;
 wire \V1/V1/V3/V2/w4 ;
 wire \V1/V1/V3/V3/w1 ;
 wire \V1/V1/V3/V3/w2 ;
 wire \V1/V1/V3/V3/w3 ;
 wire \V1/V1/V3/V3/w4 ;
 wire \V1/V1/V3/V4/w1 ;
 wire \V1/V1/V3/V4/w2 ;
 wire \V1/V1/V3/V4/w3 ;
 wire \V1/V1/V3/V4/w4 ;
 wire \V1/V1/V4/c1 ;
 wire \V1/V1/V4/c2 ;
 wire \V1/V1/V4/c3 ;
 wire \V1/V1/V4/overflow ;
 wire \V1/V1/V4/A1/c1 ;
 wire \V1/V1/V4/A1/c2 ;
 wire \V1/V1/V4/A1/c3 ;
 wire \V1/V1/V4/A1/M1/c1 ;
 wire \V1/V1/V4/A1/M1/c2 ;
 wire \V1/V1/V4/A1/M1/s1 ;
 wire \V1/V1/V4/A1/M2/c1 ;
 wire \V1/V1/V4/A1/M2/c2 ;
 wire \V1/V1/V4/A1/M2/s1 ;
 wire \V1/V1/V4/A1/M3/c1 ;
 wire \V1/V1/V4/A1/M3/c2 ;
 wire \V1/V1/V4/A1/M3/s1 ;
 wire \V1/V1/V4/A1/M4/c1 ;
 wire \V1/V1/V4/A1/M4/c2 ;
 wire \V1/V1/V4/A1/M4/s1 ;
 wire \V1/V1/V4/A2/c1 ;
 wire \V1/V1/V4/A2/c2 ;
 wire \V1/V1/V4/A2/c3 ;
 wire \V1/V1/V4/A2/M1/c1 ;
 wire \V1/V1/V4/A2/M1/c2 ;
 wire \V1/V1/V4/A2/M1/s1 ;
 wire \V1/V1/V4/A2/M2/c1 ;
 wire \V1/V1/V4/A2/M2/c2 ;
 wire \V1/V1/V4/A2/M2/s1 ;
 wire \V1/V1/V4/A2/M3/c1 ;
 wire \V1/V1/V4/A2/M3/c2 ;
 wire \V1/V1/V4/A2/M3/s1 ;
 wire \V1/V1/V4/A2/M4/c1 ;
 wire \V1/V1/V4/A2/M4/c2 ;
 wire \V1/V1/V4/A2/M4/s1 ;
 wire \V1/V1/V4/A3/c1 ;
 wire \V1/V1/V4/A3/c2 ;
 wire \V1/V1/V4/A3/c3 ;
 wire \V1/V1/V4/A3/M1/c1 ;
 wire \V1/V1/V4/A3/M1/c2 ;
 wire \V1/V1/V4/A3/M1/s1 ;
 wire \V1/V1/V4/A3/M2/c1 ;
 wire \V1/V1/V4/A3/M2/c2 ;
 wire \V1/V1/V4/A3/M2/s1 ;
 wire \V1/V1/V4/A3/M3/c1 ;
 wire \V1/V1/V4/A3/M3/c2 ;
 wire \V1/V1/V4/A3/M3/s1 ;
 wire \V1/V1/V4/A3/M4/c1 ;
 wire \V1/V1/V4/A3/M4/c2 ;
 wire \V1/V1/V4/A3/M4/s1 ;
 wire \V1/V1/V4/V1/w1 ;
 wire \V1/V1/V4/V1/w2 ;
 wire \V1/V1/V4/V1/w3 ;
 wire \V1/V1/V4/V1/w4 ;
 wire \V1/V1/V4/V2/w1 ;
 wire \V1/V1/V4/V2/w2 ;
 wire \V1/V1/V4/V2/w3 ;
 wire \V1/V1/V4/V2/w4 ;
 wire \V1/V1/V4/V3/w1 ;
 wire \V1/V1/V4/V3/w2 ;
 wire \V1/V1/V4/V3/w3 ;
 wire \V1/V1/V4/V3/w4 ;
 wire \V1/V1/V4/V4/w1 ;
 wire \V1/V1/V4/V4/w2 ;
 wire \V1/V1/V4/V4/w3 ;
 wire \V1/V1/V4/V4/w4 ;
 wire \V1/V2/c1 ;
 wire \V1/V2/c2 ;
 wire \V1/V2/c3 ;
 wire \V1/V2/overflow ;
 wire \V1/V2/A1/c1 ;
 wire \V1/V2/A1/A1/c1 ;
 wire \V1/V2/A1/A1/c2 ;
 wire \V1/V2/A1/A1/c3 ;
 wire \V1/V2/A1/A1/M1/c1 ;
 wire \V1/V2/A1/A1/M1/c2 ;
 wire \V1/V2/A1/A1/M1/s1 ;
 wire \V1/V2/A1/A1/M2/c1 ;
 wire \V1/V2/A1/A1/M2/c2 ;
 wire \V1/V2/A1/A1/M2/s1 ;
 wire \V1/V2/A1/A1/M3/c1 ;
 wire \V1/V2/A1/A1/M3/c2 ;
 wire \V1/V2/A1/A1/M3/s1 ;
 wire \V1/V2/A1/A1/M4/c1 ;
 wire \V1/V2/A1/A1/M4/c2 ;
 wire \V1/V2/A1/A1/M4/s1 ;
 wire \V1/V2/A1/A2/c1 ;
 wire \V1/V2/A1/A2/c2 ;
 wire \V1/V2/A1/A2/c3 ;
 wire \V1/V2/A1/A2/M1/c1 ;
 wire \V1/V2/A1/A2/M1/c2 ;
 wire \V1/V2/A1/A2/M1/s1 ;
 wire \V1/V2/A1/A2/M2/c1 ;
 wire \V1/V2/A1/A2/M2/c2 ;
 wire \V1/V2/A1/A2/M2/s1 ;
 wire \V1/V2/A1/A2/M3/c1 ;
 wire \V1/V2/A1/A2/M3/c2 ;
 wire \V1/V2/A1/A2/M3/s1 ;
 wire \V1/V2/A1/A2/M4/c1 ;
 wire \V1/V2/A1/A2/M4/c2 ;
 wire \V1/V2/A1/A2/M4/s1 ;
 wire \V1/V2/A2/c1 ;
 wire \V1/V2/A2/A1/c1 ;
 wire \V1/V2/A2/A1/c2 ;
 wire \V1/V2/A2/A1/c3 ;
 wire \V1/V2/A2/A1/M1/c1 ;
 wire \V1/V2/A2/A1/M1/c2 ;
 wire \V1/V2/A2/A1/M1/s1 ;
 wire \V1/V2/A2/A1/M2/c1 ;
 wire \V1/V2/A2/A1/M2/c2 ;
 wire \V1/V2/A2/A1/M2/s1 ;
 wire \V1/V2/A2/A1/M3/c1 ;
 wire \V1/V2/A2/A1/M3/c2 ;
 wire \V1/V2/A2/A1/M3/s1 ;
 wire \V1/V2/A2/A1/M4/c1 ;
 wire \V1/V2/A2/A1/M4/c2 ;
 wire \V1/V2/A2/A1/M4/s1 ;
 wire \V1/V2/A2/A2/c1 ;
 wire \V1/V2/A2/A2/c2 ;
 wire \V1/V2/A2/A2/c3 ;
 wire \V1/V2/A2/A2/M1/c1 ;
 wire \V1/V2/A2/A2/M1/c2 ;
 wire \V1/V2/A2/A2/M1/s1 ;
 wire \V1/V2/A2/A2/M2/c1 ;
 wire \V1/V2/A2/A2/M2/c2 ;
 wire \V1/V2/A2/A2/M2/s1 ;
 wire \V1/V2/A2/A2/M3/c1 ;
 wire \V1/V2/A2/A2/M3/c2 ;
 wire \V1/V2/A2/A2/M3/s1 ;
 wire \V1/V2/A2/A2/M4/c1 ;
 wire \V1/V2/A2/A2/M4/c2 ;
 wire \V1/V2/A2/A2/M4/s1 ;
 wire \V1/V2/A3/c1 ;
 wire \V1/V2/A3/A1/c1 ;
 wire \V1/V2/A3/A1/c2 ;
 wire \V1/V2/A3/A1/c3 ;
 wire \V1/V2/A3/A1/M1/c1 ;
 wire \V1/V2/A3/A1/M1/c2 ;
 wire \V1/V2/A3/A1/M1/s1 ;
 wire \V1/V2/A3/A1/M2/c1 ;
 wire \V1/V2/A3/A1/M2/c2 ;
 wire \V1/V2/A3/A1/M2/s1 ;
 wire \V1/V2/A3/A1/M3/c1 ;
 wire \V1/V2/A3/A1/M3/c2 ;
 wire \V1/V2/A3/A1/M3/s1 ;
 wire \V1/V2/A3/A1/M4/c1 ;
 wire \V1/V2/A3/A1/M4/c2 ;
 wire \V1/V2/A3/A1/M4/s1 ;
 wire \V1/V2/A3/A2/c1 ;
 wire \V1/V2/A3/A2/c2 ;
 wire \V1/V2/A3/A2/c3 ;
 wire \V1/V2/A3/A2/M1/c1 ;
 wire \V1/V2/A3/A2/M1/c2 ;
 wire \V1/V2/A3/A2/M1/s1 ;
 wire \V1/V2/A3/A2/M2/c1 ;
 wire \V1/V2/A3/A2/M2/c2 ;
 wire \V1/V2/A3/A2/M2/s1 ;
 wire \V1/V2/A3/A2/M3/c1 ;
 wire \V1/V2/A3/A2/M3/c2 ;
 wire \V1/V2/A3/A2/M3/s1 ;
 wire \V1/V2/A3/A2/M4/c1 ;
 wire \V1/V2/A3/A2/M4/c2 ;
 wire \V1/V2/A3/A2/M4/s1 ;
 wire \V1/V2/V1/c1 ;
 wire \V1/V2/V1/c2 ;
 wire \V1/V2/V1/c3 ;
 wire \V1/V2/V1/overflow ;
 wire \V1/V2/V1/A1/c1 ;
 wire \V1/V2/V1/A1/c2 ;
 wire \V1/V2/V1/A1/c3 ;
 wire \V1/V2/V1/A1/M1/c1 ;
 wire \V1/V2/V1/A1/M1/c2 ;
 wire \V1/V2/V1/A1/M1/s1 ;
 wire \V1/V2/V1/A1/M2/c1 ;
 wire \V1/V2/V1/A1/M2/c2 ;
 wire \V1/V2/V1/A1/M2/s1 ;
 wire \V1/V2/V1/A1/M3/c1 ;
 wire \V1/V2/V1/A1/M3/c2 ;
 wire \V1/V2/V1/A1/M3/s1 ;
 wire \V1/V2/V1/A1/M4/c1 ;
 wire \V1/V2/V1/A1/M4/c2 ;
 wire \V1/V2/V1/A1/M4/s1 ;
 wire \V1/V2/V1/A2/c1 ;
 wire \V1/V2/V1/A2/c2 ;
 wire \V1/V2/V1/A2/c3 ;
 wire \V1/V2/V1/A2/M1/c1 ;
 wire \V1/V2/V1/A2/M1/c2 ;
 wire \V1/V2/V1/A2/M1/s1 ;
 wire \V1/V2/V1/A2/M2/c1 ;
 wire \V1/V2/V1/A2/M2/c2 ;
 wire \V1/V2/V1/A2/M2/s1 ;
 wire \V1/V2/V1/A2/M3/c1 ;
 wire \V1/V2/V1/A2/M3/c2 ;
 wire \V1/V2/V1/A2/M3/s1 ;
 wire \V1/V2/V1/A2/M4/c1 ;
 wire \V1/V2/V1/A2/M4/c2 ;
 wire \V1/V2/V1/A2/M4/s1 ;
 wire \V1/V2/V1/A3/c1 ;
 wire \V1/V2/V1/A3/c2 ;
 wire \V1/V2/V1/A3/c3 ;
 wire \V1/V2/V1/A3/M1/c1 ;
 wire \V1/V2/V1/A3/M1/c2 ;
 wire \V1/V2/V1/A3/M1/s1 ;
 wire \V1/V2/V1/A3/M2/c1 ;
 wire \V1/V2/V1/A3/M2/c2 ;
 wire \V1/V2/V1/A3/M2/s1 ;
 wire \V1/V2/V1/A3/M3/c1 ;
 wire \V1/V2/V1/A3/M3/c2 ;
 wire \V1/V2/V1/A3/M3/s1 ;
 wire \V1/V2/V1/A3/M4/c1 ;
 wire \V1/V2/V1/A3/M4/c2 ;
 wire \V1/V2/V1/A3/M4/s1 ;
 wire \V1/V2/V1/V1/w1 ;
 wire \V1/V2/V1/V1/w2 ;
 wire \V1/V2/V1/V1/w3 ;
 wire \V1/V2/V1/V1/w4 ;
 wire \V1/V2/V1/V2/w1 ;
 wire \V1/V2/V1/V2/w2 ;
 wire \V1/V2/V1/V2/w3 ;
 wire \V1/V2/V1/V2/w4 ;
 wire \V1/V2/V1/V3/w1 ;
 wire \V1/V2/V1/V3/w2 ;
 wire \V1/V2/V1/V3/w3 ;
 wire \V1/V2/V1/V3/w4 ;
 wire \V1/V2/V1/V4/w1 ;
 wire \V1/V2/V1/V4/w2 ;
 wire \V1/V2/V1/V4/w3 ;
 wire \V1/V2/V1/V4/w4 ;
 wire \V1/V2/V2/c1 ;
 wire \V1/V2/V2/c2 ;
 wire \V1/V2/V2/c3 ;
 wire \V1/V2/V2/overflow ;
 wire \V1/V2/V2/A1/c1 ;
 wire \V1/V2/V2/A1/c2 ;
 wire \V1/V2/V2/A1/c3 ;
 wire \V1/V2/V2/A1/M1/c1 ;
 wire \V1/V2/V2/A1/M1/c2 ;
 wire \V1/V2/V2/A1/M1/s1 ;
 wire \V1/V2/V2/A1/M2/c1 ;
 wire \V1/V2/V2/A1/M2/c2 ;
 wire \V1/V2/V2/A1/M2/s1 ;
 wire \V1/V2/V2/A1/M3/c1 ;
 wire \V1/V2/V2/A1/M3/c2 ;
 wire \V1/V2/V2/A1/M3/s1 ;
 wire \V1/V2/V2/A1/M4/c1 ;
 wire \V1/V2/V2/A1/M4/c2 ;
 wire \V1/V2/V2/A1/M4/s1 ;
 wire \V1/V2/V2/A2/c1 ;
 wire \V1/V2/V2/A2/c2 ;
 wire \V1/V2/V2/A2/c3 ;
 wire \V1/V2/V2/A2/M1/c1 ;
 wire \V1/V2/V2/A2/M1/c2 ;
 wire \V1/V2/V2/A2/M1/s1 ;
 wire \V1/V2/V2/A2/M2/c1 ;
 wire \V1/V2/V2/A2/M2/c2 ;
 wire \V1/V2/V2/A2/M2/s1 ;
 wire \V1/V2/V2/A2/M3/c1 ;
 wire \V1/V2/V2/A2/M3/c2 ;
 wire \V1/V2/V2/A2/M3/s1 ;
 wire \V1/V2/V2/A2/M4/c1 ;
 wire \V1/V2/V2/A2/M4/c2 ;
 wire \V1/V2/V2/A2/M4/s1 ;
 wire \V1/V2/V2/A3/c1 ;
 wire \V1/V2/V2/A3/c2 ;
 wire \V1/V2/V2/A3/c3 ;
 wire \V1/V2/V2/A3/M1/c1 ;
 wire \V1/V2/V2/A3/M1/c2 ;
 wire \V1/V2/V2/A3/M1/s1 ;
 wire \V1/V2/V2/A3/M2/c1 ;
 wire \V1/V2/V2/A3/M2/c2 ;
 wire \V1/V2/V2/A3/M2/s1 ;
 wire \V1/V2/V2/A3/M3/c1 ;
 wire \V1/V2/V2/A3/M3/c2 ;
 wire \V1/V2/V2/A3/M3/s1 ;
 wire \V1/V2/V2/A3/M4/c1 ;
 wire \V1/V2/V2/A3/M4/c2 ;
 wire \V1/V2/V2/A3/M4/s1 ;
 wire \V1/V2/V2/V1/w1 ;
 wire \V1/V2/V2/V1/w2 ;
 wire \V1/V2/V2/V1/w3 ;
 wire \V1/V2/V2/V1/w4 ;
 wire \V1/V2/V2/V2/w1 ;
 wire \V1/V2/V2/V2/w2 ;
 wire \V1/V2/V2/V2/w3 ;
 wire \V1/V2/V2/V2/w4 ;
 wire \V1/V2/V2/V3/w1 ;
 wire \V1/V2/V2/V3/w2 ;
 wire \V1/V2/V2/V3/w3 ;
 wire \V1/V2/V2/V3/w4 ;
 wire \V1/V2/V2/V4/w1 ;
 wire \V1/V2/V2/V4/w2 ;
 wire \V1/V2/V2/V4/w3 ;
 wire \V1/V2/V2/V4/w4 ;
 wire \V1/V2/V3/c1 ;
 wire \V1/V2/V3/c2 ;
 wire \V1/V2/V3/c3 ;
 wire \V1/V2/V3/overflow ;
 wire \V1/V2/V3/A1/c1 ;
 wire \V1/V2/V3/A1/c2 ;
 wire \V1/V2/V3/A1/c3 ;
 wire \V1/V2/V3/A1/M1/c1 ;
 wire \V1/V2/V3/A1/M1/c2 ;
 wire \V1/V2/V3/A1/M1/s1 ;
 wire \V1/V2/V3/A1/M2/c1 ;
 wire \V1/V2/V3/A1/M2/c2 ;
 wire \V1/V2/V3/A1/M2/s1 ;
 wire \V1/V2/V3/A1/M3/c1 ;
 wire \V1/V2/V3/A1/M3/c2 ;
 wire \V1/V2/V3/A1/M3/s1 ;
 wire \V1/V2/V3/A1/M4/c1 ;
 wire \V1/V2/V3/A1/M4/c2 ;
 wire \V1/V2/V3/A1/M4/s1 ;
 wire \V1/V2/V3/A2/c1 ;
 wire \V1/V2/V3/A2/c2 ;
 wire \V1/V2/V3/A2/c3 ;
 wire \V1/V2/V3/A2/M1/c1 ;
 wire \V1/V2/V3/A2/M1/c2 ;
 wire \V1/V2/V3/A2/M1/s1 ;
 wire \V1/V2/V3/A2/M2/c1 ;
 wire \V1/V2/V3/A2/M2/c2 ;
 wire \V1/V2/V3/A2/M2/s1 ;
 wire \V1/V2/V3/A2/M3/c1 ;
 wire \V1/V2/V3/A2/M3/c2 ;
 wire \V1/V2/V3/A2/M3/s1 ;
 wire \V1/V2/V3/A2/M4/c1 ;
 wire \V1/V2/V3/A2/M4/c2 ;
 wire \V1/V2/V3/A2/M4/s1 ;
 wire \V1/V2/V3/A3/c1 ;
 wire \V1/V2/V3/A3/c2 ;
 wire \V1/V2/V3/A3/c3 ;
 wire \V1/V2/V3/A3/M1/c1 ;
 wire \V1/V2/V3/A3/M1/c2 ;
 wire \V1/V2/V3/A3/M1/s1 ;
 wire \V1/V2/V3/A3/M2/c1 ;
 wire \V1/V2/V3/A3/M2/c2 ;
 wire \V1/V2/V3/A3/M2/s1 ;
 wire \V1/V2/V3/A3/M3/c1 ;
 wire \V1/V2/V3/A3/M3/c2 ;
 wire \V1/V2/V3/A3/M3/s1 ;
 wire \V1/V2/V3/A3/M4/c1 ;
 wire \V1/V2/V3/A3/M4/c2 ;
 wire \V1/V2/V3/A3/M4/s1 ;
 wire \V1/V2/V3/V1/w1 ;
 wire \V1/V2/V3/V1/w2 ;
 wire \V1/V2/V3/V1/w3 ;
 wire \V1/V2/V3/V1/w4 ;
 wire \V1/V2/V3/V2/w1 ;
 wire \V1/V2/V3/V2/w2 ;
 wire \V1/V2/V3/V2/w3 ;
 wire \V1/V2/V3/V2/w4 ;
 wire \V1/V2/V3/V3/w1 ;
 wire \V1/V2/V3/V3/w2 ;
 wire \V1/V2/V3/V3/w3 ;
 wire \V1/V2/V3/V3/w4 ;
 wire \V1/V2/V3/V4/w1 ;
 wire \V1/V2/V3/V4/w2 ;
 wire \V1/V2/V3/V4/w3 ;
 wire \V1/V2/V3/V4/w4 ;
 wire \V1/V2/V4/c1 ;
 wire \V1/V2/V4/c2 ;
 wire \V1/V2/V4/c3 ;
 wire \V1/V2/V4/overflow ;
 wire \V1/V2/V4/A1/c1 ;
 wire \V1/V2/V4/A1/c2 ;
 wire \V1/V2/V4/A1/c3 ;
 wire \V1/V2/V4/A1/M1/c1 ;
 wire \V1/V2/V4/A1/M1/c2 ;
 wire \V1/V2/V4/A1/M1/s1 ;
 wire \V1/V2/V4/A1/M2/c1 ;
 wire \V1/V2/V4/A1/M2/c2 ;
 wire \V1/V2/V4/A1/M2/s1 ;
 wire \V1/V2/V4/A1/M3/c1 ;
 wire \V1/V2/V4/A1/M3/c2 ;
 wire \V1/V2/V4/A1/M3/s1 ;
 wire \V1/V2/V4/A1/M4/c1 ;
 wire \V1/V2/V4/A1/M4/c2 ;
 wire \V1/V2/V4/A1/M4/s1 ;
 wire \V1/V2/V4/A2/c1 ;
 wire \V1/V2/V4/A2/c2 ;
 wire \V1/V2/V4/A2/c3 ;
 wire \V1/V2/V4/A2/M1/c1 ;
 wire \V1/V2/V4/A2/M1/c2 ;
 wire \V1/V2/V4/A2/M1/s1 ;
 wire \V1/V2/V4/A2/M2/c1 ;
 wire \V1/V2/V4/A2/M2/c2 ;
 wire \V1/V2/V4/A2/M2/s1 ;
 wire \V1/V2/V4/A2/M3/c1 ;
 wire \V1/V2/V4/A2/M3/c2 ;
 wire \V1/V2/V4/A2/M3/s1 ;
 wire \V1/V2/V4/A2/M4/c1 ;
 wire \V1/V2/V4/A2/M4/c2 ;
 wire \V1/V2/V4/A2/M4/s1 ;
 wire \V1/V2/V4/A3/c1 ;
 wire \V1/V2/V4/A3/c2 ;
 wire \V1/V2/V4/A3/c3 ;
 wire \V1/V2/V4/A3/M1/c1 ;
 wire \V1/V2/V4/A3/M1/c2 ;
 wire \V1/V2/V4/A3/M1/s1 ;
 wire \V1/V2/V4/A3/M2/c1 ;
 wire \V1/V2/V4/A3/M2/c2 ;
 wire \V1/V2/V4/A3/M2/s1 ;
 wire \V1/V2/V4/A3/M3/c1 ;
 wire \V1/V2/V4/A3/M3/c2 ;
 wire \V1/V2/V4/A3/M3/s1 ;
 wire \V1/V2/V4/A3/M4/c1 ;
 wire \V1/V2/V4/A3/M4/c2 ;
 wire \V1/V2/V4/A3/M4/s1 ;
 wire \V1/V2/V4/V1/w1 ;
 wire \V1/V2/V4/V1/w2 ;
 wire \V1/V2/V4/V1/w3 ;
 wire \V1/V2/V4/V1/w4 ;
 wire \V1/V2/V4/V2/w1 ;
 wire \V1/V2/V4/V2/w2 ;
 wire \V1/V2/V4/V2/w3 ;
 wire \V1/V2/V4/V2/w4 ;
 wire \V1/V2/V4/V3/w1 ;
 wire \V1/V2/V4/V3/w2 ;
 wire \V1/V2/V4/V3/w3 ;
 wire \V1/V2/V4/V3/w4 ;
 wire \V1/V2/V4/V4/w1 ;
 wire \V1/V2/V4/V4/w2 ;
 wire \V1/V2/V4/V4/w3 ;
 wire \V1/V2/V4/V4/w4 ;
 wire \V1/V3/c1 ;
 wire \V1/V3/c2 ;
 wire \V1/V3/c3 ;
 wire \V1/V3/overflow ;
 wire \V1/V3/A1/c1 ;
 wire \V1/V3/A1/A1/c1 ;
 wire \V1/V3/A1/A1/c2 ;
 wire \V1/V3/A1/A1/c3 ;
 wire \V1/V3/A1/A1/M1/c1 ;
 wire \V1/V3/A1/A1/M1/c2 ;
 wire \V1/V3/A1/A1/M1/s1 ;
 wire \V1/V3/A1/A1/M2/c1 ;
 wire \V1/V3/A1/A1/M2/c2 ;
 wire \V1/V3/A1/A1/M2/s1 ;
 wire \V1/V3/A1/A1/M3/c1 ;
 wire \V1/V3/A1/A1/M3/c2 ;
 wire \V1/V3/A1/A1/M3/s1 ;
 wire \V1/V3/A1/A1/M4/c1 ;
 wire \V1/V3/A1/A1/M4/c2 ;
 wire \V1/V3/A1/A1/M4/s1 ;
 wire \V1/V3/A1/A2/c1 ;
 wire \V1/V3/A1/A2/c2 ;
 wire \V1/V3/A1/A2/c3 ;
 wire \V1/V3/A1/A2/M1/c1 ;
 wire \V1/V3/A1/A2/M1/c2 ;
 wire \V1/V3/A1/A2/M1/s1 ;
 wire \V1/V3/A1/A2/M2/c1 ;
 wire \V1/V3/A1/A2/M2/c2 ;
 wire \V1/V3/A1/A2/M2/s1 ;
 wire \V1/V3/A1/A2/M3/c1 ;
 wire \V1/V3/A1/A2/M3/c2 ;
 wire \V1/V3/A1/A2/M3/s1 ;
 wire \V1/V3/A1/A2/M4/c1 ;
 wire \V1/V3/A1/A2/M4/c2 ;
 wire \V1/V3/A1/A2/M4/s1 ;
 wire \V1/V3/A2/c1 ;
 wire \V1/V3/A2/A1/c1 ;
 wire \V1/V3/A2/A1/c2 ;
 wire \V1/V3/A2/A1/c3 ;
 wire \V1/V3/A2/A1/M1/c1 ;
 wire \V1/V3/A2/A1/M1/c2 ;
 wire \V1/V3/A2/A1/M1/s1 ;
 wire \V1/V3/A2/A1/M2/c1 ;
 wire \V1/V3/A2/A1/M2/c2 ;
 wire \V1/V3/A2/A1/M2/s1 ;
 wire \V1/V3/A2/A1/M3/c1 ;
 wire \V1/V3/A2/A1/M3/c2 ;
 wire \V1/V3/A2/A1/M3/s1 ;
 wire \V1/V3/A2/A1/M4/c1 ;
 wire \V1/V3/A2/A1/M4/c2 ;
 wire \V1/V3/A2/A1/M4/s1 ;
 wire \V1/V3/A2/A2/c1 ;
 wire \V1/V3/A2/A2/c2 ;
 wire \V1/V3/A2/A2/c3 ;
 wire \V1/V3/A2/A2/M1/c1 ;
 wire \V1/V3/A2/A2/M1/c2 ;
 wire \V1/V3/A2/A2/M1/s1 ;
 wire \V1/V3/A2/A2/M2/c1 ;
 wire \V1/V3/A2/A2/M2/c2 ;
 wire \V1/V3/A2/A2/M2/s1 ;
 wire \V1/V3/A2/A2/M3/c1 ;
 wire \V1/V3/A2/A2/M3/c2 ;
 wire \V1/V3/A2/A2/M3/s1 ;
 wire \V1/V3/A2/A2/M4/c1 ;
 wire \V1/V3/A2/A2/M4/c2 ;
 wire \V1/V3/A2/A2/M4/s1 ;
 wire \V1/V3/A3/c1 ;
 wire \V1/V3/A3/A1/c1 ;
 wire \V1/V3/A3/A1/c2 ;
 wire \V1/V3/A3/A1/c3 ;
 wire \V1/V3/A3/A1/M1/c1 ;
 wire \V1/V3/A3/A1/M1/c2 ;
 wire \V1/V3/A3/A1/M1/s1 ;
 wire \V1/V3/A3/A1/M2/c1 ;
 wire \V1/V3/A3/A1/M2/c2 ;
 wire \V1/V3/A3/A1/M2/s1 ;
 wire \V1/V3/A3/A1/M3/c1 ;
 wire \V1/V3/A3/A1/M3/c2 ;
 wire \V1/V3/A3/A1/M3/s1 ;
 wire \V1/V3/A3/A1/M4/c1 ;
 wire \V1/V3/A3/A1/M4/c2 ;
 wire \V1/V3/A3/A1/M4/s1 ;
 wire \V1/V3/A3/A2/c1 ;
 wire \V1/V3/A3/A2/c2 ;
 wire \V1/V3/A3/A2/c3 ;
 wire \V1/V3/A3/A2/M1/c1 ;
 wire \V1/V3/A3/A2/M1/c2 ;
 wire \V1/V3/A3/A2/M1/s1 ;
 wire \V1/V3/A3/A2/M2/c1 ;
 wire \V1/V3/A3/A2/M2/c2 ;
 wire \V1/V3/A3/A2/M2/s1 ;
 wire \V1/V3/A3/A2/M3/c1 ;
 wire \V1/V3/A3/A2/M3/c2 ;
 wire \V1/V3/A3/A2/M3/s1 ;
 wire \V1/V3/A3/A2/M4/c1 ;
 wire \V1/V3/A3/A2/M4/c2 ;
 wire \V1/V3/A3/A2/M4/s1 ;
 wire \V1/V3/V1/c1 ;
 wire \V1/V3/V1/c2 ;
 wire \V1/V3/V1/c3 ;
 wire \V1/V3/V1/overflow ;
 wire \V1/V3/V1/A1/c1 ;
 wire \V1/V3/V1/A1/c2 ;
 wire \V1/V3/V1/A1/c3 ;
 wire \V1/V3/V1/A1/M1/c1 ;
 wire \V1/V3/V1/A1/M1/c2 ;
 wire \V1/V3/V1/A1/M1/s1 ;
 wire \V1/V3/V1/A1/M2/c1 ;
 wire \V1/V3/V1/A1/M2/c2 ;
 wire \V1/V3/V1/A1/M2/s1 ;
 wire \V1/V3/V1/A1/M3/c1 ;
 wire \V1/V3/V1/A1/M3/c2 ;
 wire \V1/V3/V1/A1/M3/s1 ;
 wire \V1/V3/V1/A1/M4/c1 ;
 wire \V1/V3/V1/A1/M4/c2 ;
 wire \V1/V3/V1/A1/M4/s1 ;
 wire \V1/V3/V1/A2/c1 ;
 wire \V1/V3/V1/A2/c2 ;
 wire \V1/V3/V1/A2/c3 ;
 wire \V1/V3/V1/A2/M1/c1 ;
 wire \V1/V3/V1/A2/M1/c2 ;
 wire \V1/V3/V1/A2/M1/s1 ;
 wire \V1/V3/V1/A2/M2/c1 ;
 wire \V1/V3/V1/A2/M2/c2 ;
 wire \V1/V3/V1/A2/M2/s1 ;
 wire \V1/V3/V1/A2/M3/c1 ;
 wire \V1/V3/V1/A2/M3/c2 ;
 wire \V1/V3/V1/A2/M3/s1 ;
 wire \V1/V3/V1/A2/M4/c1 ;
 wire \V1/V3/V1/A2/M4/c2 ;
 wire \V1/V3/V1/A2/M4/s1 ;
 wire \V1/V3/V1/A3/c1 ;
 wire \V1/V3/V1/A3/c2 ;
 wire \V1/V3/V1/A3/c3 ;
 wire \V1/V3/V1/A3/M1/c1 ;
 wire \V1/V3/V1/A3/M1/c2 ;
 wire \V1/V3/V1/A3/M1/s1 ;
 wire \V1/V3/V1/A3/M2/c1 ;
 wire \V1/V3/V1/A3/M2/c2 ;
 wire \V1/V3/V1/A3/M2/s1 ;
 wire \V1/V3/V1/A3/M3/c1 ;
 wire \V1/V3/V1/A3/M3/c2 ;
 wire \V1/V3/V1/A3/M3/s1 ;
 wire \V1/V3/V1/A3/M4/c1 ;
 wire \V1/V3/V1/A3/M4/c2 ;
 wire \V1/V3/V1/A3/M4/s1 ;
 wire \V1/V3/V1/V1/w1 ;
 wire \V1/V3/V1/V1/w2 ;
 wire \V1/V3/V1/V1/w3 ;
 wire \V1/V3/V1/V1/w4 ;
 wire \V1/V3/V1/V2/w1 ;
 wire \V1/V3/V1/V2/w2 ;
 wire \V1/V3/V1/V2/w3 ;
 wire \V1/V3/V1/V2/w4 ;
 wire \V1/V3/V1/V3/w1 ;
 wire \V1/V3/V1/V3/w2 ;
 wire \V1/V3/V1/V3/w3 ;
 wire \V1/V3/V1/V3/w4 ;
 wire \V1/V3/V1/V4/w1 ;
 wire \V1/V3/V1/V4/w2 ;
 wire \V1/V3/V1/V4/w3 ;
 wire \V1/V3/V1/V4/w4 ;
 wire \V1/V3/V2/c1 ;
 wire \V1/V3/V2/c2 ;
 wire \V1/V3/V2/c3 ;
 wire \V1/V3/V2/overflow ;
 wire \V1/V3/V2/A1/c1 ;
 wire \V1/V3/V2/A1/c2 ;
 wire \V1/V3/V2/A1/c3 ;
 wire \V1/V3/V2/A1/M1/c1 ;
 wire \V1/V3/V2/A1/M1/c2 ;
 wire \V1/V3/V2/A1/M1/s1 ;
 wire \V1/V3/V2/A1/M2/c1 ;
 wire \V1/V3/V2/A1/M2/c2 ;
 wire \V1/V3/V2/A1/M2/s1 ;
 wire \V1/V3/V2/A1/M3/c1 ;
 wire \V1/V3/V2/A1/M3/c2 ;
 wire \V1/V3/V2/A1/M3/s1 ;
 wire \V1/V3/V2/A1/M4/c1 ;
 wire \V1/V3/V2/A1/M4/c2 ;
 wire \V1/V3/V2/A1/M4/s1 ;
 wire \V1/V3/V2/A2/c1 ;
 wire \V1/V3/V2/A2/c2 ;
 wire \V1/V3/V2/A2/c3 ;
 wire \V1/V3/V2/A2/M1/c1 ;
 wire \V1/V3/V2/A2/M1/c2 ;
 wire \V1/V3/V2/A2/M1/s1 ;
 wire \V1/V3/V2/A2/M2/c1 ;
 wire \V1/V3/V2/A2/M2/c2 ;
 wire \V1/V3/V2/A2/M2/s1 ;
 wire \V1/V3/V2/A2/M3/c1 ;
 wire \V1/V3/V2/A2/M3/c2 ;
 wire \V1/V3/V2/A2/M3/s1 ;
 wire \V1/V3/V2/A2/M4/c1 ;
 wire \V1/V3/V2/A2/M4/c2 ;
 wire \V1/V3/V2/A2/M4/s1 ;
 wire \V1/V3/V2/A3/c1 ;
 wire \V1/V3/V2/A3/c2 ;
 wire \V1/V3/V2/A3/c3 ;
 wire \V1/V3/V2/A3/M1/c1 ;
 wire \V1/V3/V2/A3/M1/c2 ;
 wire \V1/V3/V2/A3/M1/s1 ;
 wire \V1/V3/V2/A3/M2/c1 ;
 wire \V1/V3/V2/A3/M2/c2 ;
 wire \V1/V3/V2/A3/M2/s1 ;
 wire \V1/V3/V2/A3/M3/c1 ;
 wire \V1/V3/V2/A3/M3/c2 ;
 wire \V1/V3/V2/A3/M3/s1 ;
 wire \V1/V3/V2/A3/M4/c1 ;
 wire \V1/V3/V2/A3/M4/c2 ;
 wire \V1/V3/V2/A3/M4/s1 ;
 wire \V1/V3/V2/V1/w1 ;
 wire \V1/V3/V2/V1/w2 ;
 wire \V1/V3/V2/V1/w3 ;
 wire \V1/V3/V2/V1/w4 ;
 wire \V1/V3/V2/V2/w1 ;
 wire \V1/V3/V2/V2/w2 ;
 wire \V1/V3/V2/V2/w3 ;
 wire \V1/V3/V2/V2/w4 ;
 wire \V1/V3/V2/V3/w1 ;
 wire \V1/V3/V2/V3/w2 ;
 wire \V1/V3/V2/V3/w3 ;
 wire \V1/V3/V2/V3/w4 ;
 wire \V1/V3/V2/V4/w1 ;
 wire \V1/V3/V2/V4/w2 ;
 wire \V1/V3/V2/V4/w3 ;
 wire \V1/V3/V2/V4/w4 ;
 wire \V1/V3/V3/c1 ;
 wire \V1/V3/V3/c2 ;
 wire \V1/V3/V3/c3 ;
 wire \V1/V3/V3/overflow ;
 wire \V1/V3/V3/A1/c1 ;
 wire \V1/V3/V3/A1/c2 ;
 wire \V1/V3/V3/A1/c3 ;
 wire \V1/V3/V3/A1/M1/c1 ;
 wire \V1/V3/V3/A1/M1/c2 ;
 wire \V1/V3/V3/A1/M1/s1 ;
 wire \V1/V3/V3/A1/M2/c1 ;
 wire \V1/V3/V3/A1/M2/c2 ;
 wire \V1/V3/V3/A1/M2/s1 ;
 wire \V1/V3/V3/A1/M3/c1 ;
 wire \V1/V3/V3/A1/M3/c2 ;
 wire \V1/V3/V3/A1/M3/s1 ;
 wire \V1/V3/V3/A1/M4/c1 ;
 wire \V1/V3/V3/A1/M4/c2 ;
 wire \V1/V3/V3/A1/M4/s1 ;
 wire \V1/V3/V3/A2/c1 ;
 wire \V1/V3/V3/A2/c2 ;
 wire \V1/V3/V3/A2/c3 ;
 wire \V1/V3/V3/A2/M1/c1 ;
 wire \V1/V3/V3/A2/M1/c2 ;
 wire \V1/V3/V3/A2/M1/s1 ;
 wire \V1/V3/V3/A2/M2/c1 ;
 wire \V1/V3/V3/A2/M2/c2 ;
 wire \V1/V3/V3/A2/M2/s1 ;
 wire \V1/V3/V3/A2/M3/c1 ;
 wire \V1/V3/V3/A2/M3/c2 ;
 wire \V1/V3/V3/A2/M3/s1 ;
 wire \V1/V3/V3/A2/M4/c1 ;
 wire \V1/V3/V3/A2/M4/c2 ;
 wire \V1/V3/V3/A2/M4/s1 ;
 wire \V1/V3/V3/A3/c1 ;
 wire \V1/V3/V3/A3/c2 ;
 wire \V1/V3/V3/A3/c3 ;
 wire \V1/V3/V3/A3/M1/c1 ;
 wire \V1/V3/V3/A3/M1/c2 ;
 wire \V1/V3/V3/A3/M1/s1 ;
 wire \V1/V3/V3/A3/M2/c1 ;
 wire \V1/V3/V3/A3/M2/c2 ;
 wire \V1/V3/V3/A3/M2/s1 ;
 wire \V1/V3/V3/A3/M3/c1 ;
 wire \V1/V3/V3/A3/M3/c2 ;
 wire \V1/V3/V3/A3/M3/s1 ;
 wire \V1/V3/V3/A3/M4/c1 ;
 wire \V1/V3/V3/A3/M4/c2 ;
 wire \V1/V3/V3/A3/M4/s1 ;
 wire \V1/V3/V3/V1/w1 ;
 wire \V1/V3/V3/V1/w2 ;
 wire \V1/V3/V3/V1/w3 ;
 wire \V1/V3/V3/V1/w4 ;
 wire \V1/V3/V3/V2/w1 ;
 wire \V1/V3/V3/V2/w2 ;
 wire \V1/V3/V3/V2/w3 ;
 wire \V1/V3/V3/V2/w4 ;
 wire \V1/V3/V3/V3/w1 ;
 wire \V1/V3/V3/V3/w2 ;
 wire \V1/V3/V3/V3/w3 ;
 wire \V1/V3/V3/V3/w4 ;
 wire \V1/V3/V3/V4/w1 ;
 wire \V1/V3/V3/V4/w2 ;
 wire \V1/V3/V3/V4/w3 ;
 wire \V1/V3/V3/V4/w4 ;
 wire \V1/V3/V4/c1 ;
 wire \V1/V3/V4/c2 ;
 wire \V1/V3/V4/c3 ;
 wire \V1/V3/V4/overflow ;
 wire \V1/V3/V4/A1/c1 ;
 wire \V1/V3/V4/A1/c2 ;
 wire \V1/V3/V4/A1/c3 ;
 wire \V1/V3/V4/A1/M1/c1 ;
 wire \V1/V3/V4/A1/M1/c2 ;
 wire \V1/V3/V4/A1/M1/s1 ;
 wire \V1/V3/V4/A1/M2/c1 ;
 wire \V1/V3/V4/A1/M2/c2 ;
 wire \V1/V3/V4/A1/M2/s1 ;
 wire \V1/V3/V4/A1/M3/c1 ;
 wire \V1/V3/V4/A1/M3/c2 ;
 wire \V1/V3/V4/A1/M3/s1 ;
 wire \V1/V3/V4/A1/M4/c1 ;
 wire \V1/V3/V4/A1/M4/c2 ;
 wire \V1/V3/V4/A1/M4/s1 ;
 wire \V1/V3/V4/A2/c1 ;
 wire \V1/V3/V4/A2/c2 ;
 wire \V1/V3/V4/A2/c3 ;
 wire \V1/V3/V4/A2/M1/c1 ;
 wire \V1/V3/V4/A2/M1/c2 ;
 wire \V1/V3/V4/A2/M1/s1 ;
 wire \V1/V3/V4/A2/M2/c1 ;
 wire \V1/V3/V4/A2/M2/c2 ;
 wire \V1/V3/V4/A2/M2/s1 ;
 wire \V1/V3/V4/A2/M3/c1 ;
 wire \V1/V3/V4/A2/M3/c2 ;
 wire \V1/V3/V4/A2/M3/s1 ;
 wire \V1/V3/V4/A2/M4/c1 ;
 wire \V1/V3/V4/A2/M4/c2 ;
 wire \V1/V3/V4/A2/M4/s1 ;
 wire \V1/V3/V4/A3/c1 ;
 wire \V1/V3/V4/A3/c2 ;
 wire \V1/V3/V4/A3/c3 ;
 wire \V1/V3/V4/A3/M1/c1 ;
 wire \V1/V3/V4/A3/M1/c2 ;
 wire \V1/V3/V4/A3/M1/s1 ;
 wire \V1/V3/V4/A3/M2/c1 ;
 wire \V1/V3/V4/A3/M2/c2 ;
 wire \V1/V3/V4/A3/M2/s1 ;
 wire \V1/V3/V4/A3/M3/c1 ;
 wire \V1/V3/V4/A3/M3/c2 ;
 wire \V1/V3/V4/A3/M3/s1 ;
 wire \V1/V3/V4/A3/M4/c1 ;
 wire \V1/V3/V4/A3/M4/c2 ;
 wire \V1/V3/V4/A3/M4/s1 ;
 wire \V1/V3/V4/V1/w1 ;
 wire \V1/V3/V4/V1/w2 ;
 wire \V1/V3/V4/V1/w3 ;
 wire \V1/V3/V4/V1/w4 ;
 wire \V1/V3/V4/V2/w1 ;
 wire \V1/V3/V4/V2/w2 ;
 wire \V1/V3/V4/V2/w3 ;
 wire \V1/V3/V4/V2/w4 ;
 wire \V1/V3/V4/V3/w1 ;
 wire \V1/V3/V4/V3/w2 ;
 wire \V1/V3/V4/V3/w3 ;
 wire \V1/V3/V4/V3/w4 ;
 wire \V1/V3/V4/V4/w1 ;
 wire \V1/V3/V4/V4/w2 ;
 wire \V1/V3/V4/V4/w3 ;
 wire \V1/V3/V4/V4/w4 ;
 wire \V1/V4/c1 ;
 wire \V1/V4/c2 ;
 wire \V1/V4/c3 ;
 wire \V1/V4/overflow ;
 wire \V1/V4/A1/c1 ;
 wire \V1/V4/A1/A1/c1 ;
 wire \V1/V4/A1/A1/c2 ;
 wire \V1/V4/A1/A1/c3 ;
 wire \V1/V4/A1/A1/M1/c1 ;
 wire \V1/V4/A1/A1/M1/c2 ;
 wire \V1/V4/A1/A1/M1/s1 ;
 wire \V1/V4/A1/A1/M2/c1 ;
 wire \V1/V4/A1/A1/M2/c2 ;
 wire \V1/V4/A1/A1/M2/s1 ;
 wire \V1/V4/A1/A1/M3/c1 ;
 wire \V1/V4/A1/A1/M3/c2 ;
 wire \V1/V4/A1/A1/M3/s1 ;
 wire \V1/V4/A1/A1/M4/c1 ;
 wire \V1/V4/A1/A1/M4/c2 ;
 wire \V1/V4/A1/A1/M4/s1 ;
 wire \V1/V4/A1/A2/c1 ;
 wire \V1/V4/A1/A2/c2 ;
 wire \V1/V4/A1/A2/c3 ;
 wire \V1/V4/A1/A2/M1/c1 ;
 wire \V1/V4/A1/A2/M1/c2 ;
 wire \V1/V4/A1/A2/M1/s1 ;
 wire \V1/V4/A1/A2/M2/c1 ;
 wire \V1/V4/A1/A2/M2/c2 ;
 wire \V1/V4/A1/A2/M2/s1 ;
 wire \V1/V4/A1/A2/M3/c1 ;
 wire \V1/V4/A1/A2/M3/c2 ;
 wire \V1/V4/A1/A2/M3/s1 ;
 wire \V1/V4/A1/A2/M4/c1 ;
 wire \V1/V4/A1/A2/M4/c2 ;
 wire \V1/V4/A1/A2/M4/s1 ;
 wire \V1/V4/A2/c1 ;
 wire \V1/V4/A2/A1/c1 ;
 wire \V1/V4/A2/A1/c2 ;
 wire \V1/V4/A2/A1/c3 ;
 wire \V1/V4/A2/A1/M1/c1 ;
 wire \V1/V4/A2/A1/M1/c2 ;
 wire \V1/V4/A2/A1/M1/s1 ;
 wire \V1/V4/A2/A1/M2/c1 ;
 wire \V1/V4/A2/A1/M2/c2 ;
 wire \V1/V4/A2/A1/M2/s1 ;
 wire \V1/V4/A2/A1/M3/c1 ;
 wire \V1/V4/A2/A1/M3/c2 ;
 wire \V1/V4/A2/A1/M3/s1 ;
 wire \V1/V4/A2/A1/M4/c1 ;
 wire \V1/V4/A2/A1/M4/c2 ;
 wire \V1/V4/A2/A1/M4/s1 ;
 wire \V1/V4/A2/A2/c1 ;
 wire \V1/V4/A2/A2/c2 ;
 wire \V1/V4/A2/A2/c3 ;
 wire \V1/V4/A2/A2/M1/c1 ;
 wire \V1/V4/A2/A2/M1/c2 ;
 wire \V1/V4/A2/A2/M1/s1 ;
 wire \V1/V4/A2/A2/M2/c1 ;
 wire \V1/V4/A2/A2/M2/c2 ;
 wire \V1/V4/A2/A2/M2/s1 ;
 wire \V1/V4/A2/A2/M3/c1 ;
 wire \V1/V4/A2/A2/M3/c2 ;
 wire \V1/V4/A2/A2/M3/s1 ;
 wire \V1/V4/A2/A2/M4/c1 ;
 wire \V1/V4/A2/A2/M4/c2 ;
 wire \V1/V4/A2/A2/M4/s1 ;
 wire \V1/V4/A3/c1 ;
 wire \V1/V4/A3/A1/c1 ;
 wire \V1/V4/A3/A1/c2 ;
 wire \V1/V4/A3/A1/c3 ;
 wire \V1/V4/A3/A1/M1/c1 ;
 wire \V1/V4/A3/A1/M1/c2 ;
 wire \V1/V4/A3/A1/M1/s1 ;
 wire \V1/V4/A3/A1/M2/c1 ;
 wire \V1/V4/A3/A1/M2/c2 ;
 wire \V1/V4/A3/A1/M2/s1 ;
 wire \V1/V4/A3/A1/M3/c1 ;
 wire \V1/V4/A3/A1/M3/c2 ;
 wire \V1/V4/A3/A1/M3/s1 ;
 wire \V1/V4/A3/A1/M4/c1 ;
 wire \V1/V4/A3/A1/M4/c2 ;
 wire \V1/V4/A3/A1/M4/s1 ;
 wire \V1/V4/A3/A2/c1 ;
 wire \V1/V4/A3/A2/c2 ;
 wire \V1/V4/A3/A2/c3 ;
 wire \V1/V4/A3/A2/M1/c1 ;
 wire \V1/V4/A3/A2/M1/c2 ;
 wire \V1/V4/A3/A2/M1/s1 ;
 wire \V1/V4/A3/A2/M2/c1 ;
 wire \V1/V4/A3/A2/M2/c2 ;
 wire \V1/V4/A3/A2/M2/s1 ;
 wire \V1/V4/A3/A2/M3/c1 ;
 wire \V1/V4/A3/A2/M3/c2 ;
 wire \V1/V4/A3/A2/M3/s1 ;
 wire \V1/V4/A3/A2/M4/c1 ;
 wire \V1/V4/A3/A2/M4/c2 ;
 wire \V1/V4/A3/A2/M4/s1 ;
 wire \V1/V4/V1/c1 ;
 wire \V1/V4/V1/c2 ;
 wire \V1/V4/V1/c3 ;
 wire \V1/V4/V1/overflow ;
 wire \V1/V4/V1/A1/c1 ;
 wire \V1/V4/V1/A1/c2 ;
 wire \V1/V4/V1/A1/c3 ;
 wire \V1/V4/V1/A1/M1/c1 ;
 wire \V1/V4/V1/A1/M1/c2 ;
 wire \V1/V4/V1/A1/M1/s1 ;
 wire \V1/V4/V1/A1/M2/c1 ;
 wire \V1/V4/V1/A1/M2/c2 ;
 wire \V1/V4/V1/A1/M2/s1 ;
 wire \V1/V4/V1/A1/M3/c1 ;
 wire \V1/V4/V1/A1/M3/c2 ;
 wire \V1/V4/V1/A1/M3/s1 ;
 wire \V1/V4/V1/A1/M4/c1 ;
 wire \V1/V4/V1/A1/M4/c2 ;
 wire \V1/V4/V1/A1/M4/s1 ;
 wire \V1/V4/V1/A2/c1 ;
 wire \V1/V4/V1/A2/c2 ;
 wire \V1/V4/V1/A2/c3 ;
 wire \V1/V4/V1/A2/M1/c1 ;
 wire \V1/V4/V1/A2/M1/c2 ;
 wire \V1/V4/V1/A2/M1/s1 ;
 wire \V1/V4/V1/A2/M2/c1 ;
 wire \V1/V4/V1/A2/M2/c2 ;
 wire \V1/V4/V1/A2/M2/s1 ;
 wire \V1/V4/V1/A2/M3/c1 ;
 wire \V1/V4/V1/A2/M3/c2 ;
 wire \V1/V4/V1/A2/M3/s1 ;
 wire \V1/V4/V1/A2/M4/c1 ;
 wire \V1/V4/V1/A2/M4/c2 ;
 wire \V1/V4/V1/A2/M4/s1 ;
 wire \V1/V4/V1/A3/c1 ;
 wire \V1/V4/V1/A3/c2 ;
 wire \V1/V4/V1/A3/c3 ;
 wire \V1/V4/V1/A3/M1/c1 ;
 wire \V1/V4/V1/A3/M1/c2 ;
 wire \V1/V4/V1/A3/M1/s1 ;
 wire \V1/V4/V1/A3/M2/c1 ;
 wire \V1/V4/V1/A3/M2/c2 ;
 wire \V1/V4/V1/A3/M2/s1 ;
 wire \V1/V4/V1/A3/M3/c1 ;
 wire \V1/V4/V1/A3/M3/c2 ;
 wire \V1/V4/V1/A3/M3/s1 ;
 wire \V1/V4/V1/A3/M4/c1 ;
 wire \V1/V4/V1/A3/M4/c2 ;
 wire \V1/V4/V1/A3/M4/s1 ;
 wire \V1/V4/V1/V1/w1 ;
 wire \V1/V4/V1/V1/w2 ;
 wire \V1/V4/V1/V1/w3 ;
 wire \V1/V4/V1/V1/w4 ;
 wire \V1/V4/V1/V2/w1 ;
 wire \V1/V4/V1/V2/w2 ;
 wire \V1/V4/V1/V2/w3 ;
 wire \V1/V4/V1/V2/w4 ;
 wire \V1/V4/V1/V3/w1 ;
 wire \V1/V4/V1/V3/w2 ;
 wire \V1/V4/V1/V3/w3 ;
 wire \V1/V4/V1/V3/w4 ;
 wire \V1/V4/V1/V4/w1 ;
 wire \V1/V4/V1/V4/w2 ;
 wire \V1/V4/V1/V4/w3 ;
 wire \V1/V4/V1/V4/w4 ;
 wire \V1/V4/V2/c1 ;
 wire \V1/V4/V2/c2 ;
 wire \V1/V4/V2/c3 ;
 wire \V1/V4/V2/overflow ;
 wire \V1/V4/V2/A1/c1 ;
 wire \V1/V4/V2/A1/c2 ;
 wire \V1/V4/V2/A1/c3 ;
 wire \V1/V4/V2/A1/M1/c1 ;
 wire \V1/V4/V2/A1/M1/c2 ;
 wire \V1/V4/V2/A1/M1/s1 ;
 wire \V1/V4/V2/A1/M2/c1 ;
 wire \V1/V4/V2/A1/M2/c2 ;
 wire \V1/V4/V2/A1/M2/s1 ;
 wire \V1/V4/V2/A1/M3/c1 ;
 wire \V1/V4/V2/A1/M3/c2 ;
 wire \V1/V4/V2/A1/M3/s1 ;
 wire \V1/V4/V2/A1/M4/c1 ;
 wire \V1/V4/V2/A1/M4/c2 ;
 wire \V1/V4/V2/A1/M4/s1 ;
 wire \V1/V4/V2/A2/c1 ;
 wire \V1/V4/V2/A2/c2 ;
 wire \V1/V4/V2/A2/c3 ;
 wire \V1/V4/V2/A2/M1/c1 ;
 wire \V1/V4/V2/A2/M1/c2 ;
 wire \V1/V4/V2/A2/M1/s1 ;
 wire \V1/V4/V2/A2/M2/c1 ;
 wire \V1/V4/V2/A2/M2/c2 ;
 wire \V1/V4/V2/A2/M2/s1 ;
 wire \V1/V4/V2/A2/M3/c1 ;
 wire \V1/V4/V2/A2/M3/c2 ;
 wire \V1/V4/V2/A2/M3/s1 ;
 wire \V1/V4/V2/A2/M4/c1 ;
 wire \V1/V4/V2/A2/M4/c2 ;
 wire \V1/V4/V2/A2/M4/s1 ;
 wire \V1/V4/V2/A3/c1 ;
 wire \V1/V4/V2/A3/c2 ;
 wire \V1/V4/V2/A3/c3 ;
 wire \V1/V4/V2/A3/M1/c1 ;
 wire \V1/V4/V2/A3/M1/c2 ;
 wire \V1/V4/V2/A3/M1/s1 ;
 wire \V1/V4/V2/A3/M2/c1 ;
 wire \V1/V4/V2/A3/M2/c2 ;
 wire \V1/V4/V2/A3/M2/s1 ;
 wire \V1/V4/V2/A3/M3/c1 ;
 wire \V1/V4/V2/A3/M3/c2 ;
 wire \V1/V4/V2/A3/M3/s1 ;
 wire \V1/V4/V2/A3/M4/c1 ;
 wire \V1/V4/V2/A3/M4/c2 ;
 wire \V1/V4/V2/A3/M4/s1 ;
 wire \V1/V4/V2/V1/w1 ;
 wire \V1/V4/V2/V1/w2 ;
 wire \V1/V4/V2/V1/w3 ;
 wire \V1/V4/V2/V1/w4 ;
 wire \V1/V4/V2/V2/w1 ;
 wire \V1/V4/V2/V2/w2 ;
 wire \V1/V4/V2/V2/w3 ;
 wire \V1/V4/V2/V2/w4 ;
 wire \V1/V4/V2/V3/w1 ;
 wire \V1/V4/V2/V3/w2 ;
 wire \V1/V4/V2/V3/w3 ;
 wire \V1/V4/V2/V3/w4 ;
 wire \V1/V4/V2/V4/w1 ;
 wire \V1/V4/V2/V4/w2 ;
 wire \V1/V4/V2/V4/w3 ;
 wire \V1/V4/V2/V4/w4 ;
 wire \V1/V4/V3/c1 ;
 wire \V1/V4/V3/c2 ;
 wire \V1/V4/V3/c3 ;
 wire \V1/V4/V3/overflow ;
 wire \V1/V4/V3/A1/c1 ;
 wire \V1/V4/V3/A1/c2 ;
 wire \V1/V4/V3/A1/c3 ;
 wire \V1/V4/V3/A1/M1/c1 ;
 wire \V1/V4/V3/A1/M1/c2 ;
 wire \V1/V4/V3/A1/M1/s1 ;
 wire \V1/V4/V3/A1/M2/c1 ;
 wire \V1/V4/V3/A1/M2/c2 ;
 wire \V1/V4/V3/A1/M2/s1 ;
 wire \V1/V4/V3/A1/M3/c1 ;
 wire \V1/V4/V3/A1/M3/c2 ;
 wire \V1/V4/V3/A1/M3/s1 ;
 wire \V1/V4/V3/A1/M4/c1 ;
 wire \V1/V4/V3/A1/M4/c2 ;
 wire \V1/V4/V3/A1/M4/s1 ;
 wire \V1/V4/V3/A2/c1 ;
 wire \V1/V4/V3/A2/c2 ;
 wire \V1/V4/V3/A2/c3 ;
 wire \V1/V4/V3/A2/M1/c1 ;
 wire \V1/V4/V3/A2/M1/c2 ;
 wire \V1/V4/V3/A2/M1/s1 ;
 wire \V1/V4/V3/A2/M2/c1 ;
 wire \V1/V4/V3/A2/M2/c2 ;
 wire \V1/V4/V3/A2/M2/s1 ;
 wire \V1/V4/V3/A2/M3/c1 ;
 wire \V1/V4/V3/A2/M3/c2 ;
 wire \V1/V4/V3/A2/M3/s1 ;
 wire \V1/V4/V3/A2/M4/c1 ;
 wire \V1/V4/V3/A2/M4/c2 ;
 wire \V1/V4/V3/A2/M4/s1 ;
 wire \V1/V4/V3/A3/c1 ;
 wire \V1/V4/V3/A3/c2 ;
 wire \V1/V4/V3/A3/c3 ;
 wire \V1/V4/V3/A3/M1/c1 ;
 wire \V1/V4/V3/A3/M1/c2 ;
 wire \V1/V4/V3/A3/M1/s1 ;
 wire \V1/V4/V3/A3/M2/c1 ;
 wire \V1/V4/V3/A3/M2/c2 ;
 wire \V1/V4/V3/A3/M2/s1 ;
 wire \V1/V4/V3/A3/M3/c1 ;
 wire \V1/V4/V3/A3/M3/c2 ;
 wire \V1/V4/V3/A3/M3/s1 ;
 wire \V1/V4/V3/A3/M4/c1 ;
 wire \V1/V4/V3/A3/M4/c2 ;
 wire \V1/V4/V3/A3/M4/s1 ;
 wire \V1/V4/V3/V1/w1 ;
 wire \V1/V4/V3/V1/w2 ;
 wire \V1/V4/V3/V1/w3 ;
 wire \V1/V4/V3/V1/w4 ;
 wire \V1/V4/V3/V2/w1 ;
 wire \V1/V4/V3/V2/w2 ;
 wire \V1/V4/V3/V2/w3 ;
 wire \V1/V4/V3/V2/w4 ;
 wire \V1/V4/V3/V3/w1 ;
 wire \V1/V4/V3/V3/w2 ;
 wire \V1/V4/V3/V3/w3 ;
 wire \V1/V4/V3/V3/w4 ;
 wire \V1/V4/V3/V4/w1 ;
 wire \V1/V4/V3/V4/w2 ;
 wire \V1/V4/V3/V4/w3 ;
 wire \V1/V4/V3/V4/w4 ;
 wire \V1/V4/V4/c1 ;
 wire \V1/V4/V4/c2 ;
 wire \V1/V4/V4/c3 ;
 wire \V1/V4/V4/overflow ;
 wire \V1/V4/V4/A1/c1 ;
 wire \V1/V4/V4/A1/c2 ;
 wire \V1/V4/V4/A1/c3 ;
 wire \V1/V4/V4/A1/M1/c1 ;
 wire \V1/V4/V4/A1/M1/c2 ;
 wire \V1/V4/V4/A1/M1/s1 ;
 wire \V1/V4/V4/A1/M2/c1 ;
 wire \V1/V4/V4/A1/M2/c2 ;
 wire \V1/V4/V4/A1/M2/s1 ;
 wire \V1/V4/V4/A1/M3/c1 ;
 wire \V1/V4/V4/A1/M3/c2 ;
 wire \V1/V4/V4/A1/M3/s1 ;
 wire \V1/V4/V4/A1/M4/c1 ;
 wire \V1/V4/V4/A1/M4/c2 ;
 wire \V1/V4/V4/A1/M4/s1 ;
 wire \V1/V4/V4/A2/c1 ;
 wire \V1/V4/V4/A2/c2 ;
 wire \V1/V4/V4/A2/c3 ;
 wire \V1/V4/V4/A2/M1/c1 ;
 wire \V1/V4/V4/A2/M1/c2 ;
 wire \V1/V4/V4/A2/M1/s1 ;
 wire \V1/V4/V4/A2/M2/c1 ;
 wire \V1/V4/V4/A2/M2/c2 ;
 wire \V1/V4/V4/A2/M2/s1 ;
 wire \V1/V4/V4/A2/M3/c1 ;
 wire \V1/V4/V4/A2/M3/c2 ;
 wire \V1/V4/V4/A2/M3/s1 ;
 wire \V1/V4/V4/A2/M4/c1 ;
 wire \V1/V4/V4/A2/M4/c2 ;
 wire \V1/V4/V4/A2/M4/s1 ;
 wire \V1/V4/V4/A3/c1 ;
 wire \V1/V4/V4/A3/c2 ;
 wire \V1/V4/V4/A3/c3 ;
 wire \V1/V4/V4/A3/M1/c1 ;
 wire \V1/V4/V4/A3/M1/c2 ;
 wire \V1/V4/V4/A3/M1/s1 ;
 wire \V1/V4/V4/A3/M2/c1 ;
 wire \V1/V4/V4/A3/M2/c2 ;
 wire \V1/V4/V4/A3/M2/s1 ;
 wire \V1/V4/V4/A3/M3/c1 ;
 wire \V1/V4/V4/A3/M3/c2 ;
 wire \V1/V4/V4/A3/M3/s1 ;
 wire \V1/V4/V4/A3/M4/c1 ;
 wire \V1/V4/V4/A3/M4/c2 ;
 wire \V1/V4/V4/A3/M4/s1 ;
 wire \V1/V4/V4/V1/w1 ;
 wire \V1/V4/V4/V1/w2 ;
 wire \V1/V4/V4/V1/w3 ;
 wire \V1/V4/V4/V1/w4 ;
 wire \V1/V4/V4/V2/w1 ;
 wire \V1/V4/V4/V2/w2 ;
 wire \V1/V4/V4/V2/w3 ;
 wire \V1/V4/V4/V2/w4 ;
 wire \V1/V4/V4/V3/w1 ;
 wire \V1/V4/V4/V3/w2 ;
 wire \V1/V4/V4/V3/w3 ;
 wire \V1/V4/V4/V3/w4 ;
 wire \V1/V4/V4/V4/w1 ;
 wire \V1/V4/V4/V4/w2 ;
 wire \V1/V4/V4/V4/w3 ;
 wire \V1/V4/V4/V4/w4 ;
 wire \V2/c1 ;
 wire \V2/c2 ;
 wire \V2/c3 ;
 wire \V2/overflow ;
 wire \V2/A1/c1 ;
 wire \V2/A1/A1/c1 ;
 wire \V2/A1/A1/A1/c1 ;
 wire \V2/A1/A1/A1/c2 ;
 wire \V2/A1/A1/A1/c3 ;
 wire \V2/A1/A1/A1/M1/c1 ;
 wire \V2/A1/A1/A1/M1/c2 ;
 wire \V2/A1/A1/A1/M1/s1 ;
 wire \V2/A1/A1/A1/M2/c1 ;
 wire \V2/A1/A1/A1/M2/c2 ;
 wire \V2/A1/A1/A1/M2/s1 ;
 wire \V2/A1/A1/A1/M3/c1 ;
 wire \V2/A1/A1/A1/M3/c2 ;
 wire \V2/A1/A1/A1/M3/s1 ;
 wire \V2/A1/A1/A1/M4/c1 ;
 wire \V2/A1/A1/A1/M4/c2 ;
 wire \V2/A1/A1/A1/M4/s1 ;
 wire \V2/A1/A1/A2/c1 ;
 wire \V2/A1/A1/A2/c2 ;
 wire \V2/A1/A1/A2/c3 ;
 wire \V2/A1/A1/A2/M1/c1 ;
 wire \V2/A1/A1/A2/M1/c2 ;
 wire \V2/A1/A1/A2/M1/s1 ;
 wire \V2/A1/A1/A2/M2/c1 ;
 wire \V2/A1/A1/A2/M2/c2 ;
 wire \V2/A1/A1/A2/M2/s1 ;
 wire \V2/A1/A1/A2/M3/c1 ;
 wire \V2/A1/A1/A2/M3/c2 ;
 wire \V2/A1/A1/A2/M3/s1 ;
 wire \V2/A1/A1/A2/M4/c1 ;
 wire \V2/A1/A1/A2/M4/c2 ;
 wire \V2/A1/A1/A2/M4/s1 ;
 wire \V2/A1/A2/c1 ;
 wire \V2/A1/A2/A1/c1 ;
 wire \V2/A1/A2/A1/c2 ;
 wire \V2/A1/A2/A1/c3 ;
 wire \V2/A1/A2/A1/M1/c1 ;
 wire \V2/A1/A2/A1/M1/c2 ;
 wire \V2/A1/A2/A1/M1/s1 ;
 wire \V2/A1/A2/A1/M2/c1 ;
 wire \V2/A1/A2/A1/M2/c2 ;
 wire \V2/A1/A2/A1/M2/s1 ;
 wire \V2/A1/A2/A1/M3/c1 ;
 wire \V2/A1/A2/A1/M3/c2 ;
 wire \V2/A1/A2/A1/M3/s1 ;
 wire \V2/A1/A2/A1/M4/c1 ;
 wire \V2/A1/A2/A1/M4/c2 ;
 wire \V2/A1/A2/A1/M4/s1 ;
 wire \V2/A1/A2/A2/c1 ;
 wire \V2/A1/A2/A2/c2 ;
 wire \V2/A1/A2/A2/c3 ;
 wire \V2/A1/A2/A2/M1/c1 ;
 wire \V2/A1/A2/A2/M1/c2 ;
 wire \V2/A1/A2/A2/M1/s1 ;
 wire \V2/A1/A2/A2/M2/c1 ;
 wire \V2/A1/A2/A2/M2/c2 ;
 wire \V2/A1/A2/A2/M2/s1 ;
 wire \V2/A1/A2/A2/M3/c1 ;
 wire \V2/A1/A2/A2/M3/c2 ;
 wire \V2/A1/A2/A2/M3/s1 ;
 wire \V2/A1/A2/A2/M4/c1 ;
 wire \V2/A1/A2/A2/M4/c2 ;
 wire \V2/A1/A2/A2/M4/s1 ;
 wire \V2/A2/c1 ;
 wire \V2/A2/A1/c1 ;
 wire \V2/A2/A1/A1/c1 ;
 wire \V2/A2/A1/A1/c2 ;
 wire \V2/A2/A1/A1/c3 ;
 wire \V2/A2/A1/A1/M1/c1 ;
 wire \V2/A2/A1/A1/M1/c2 ;
 wire \V2/A2/A1/A1/M1/s1 ;
 wire \V2/A2/A1/A1/M2/c1 ;
 wire \V2/A2/A1/A1/M2/c2 ;
 wire \V2/A2/A1/A1/M2/s1 ;
 wire \V2/A2/A1/A1/M3/c1 ;
 wire \V2/A2/A1/A1/M3/c2 ;
 wire \V2/A2/A1/A1/M3/s1 ;
 wire \V2/A2/A1/A1/M4/c1 ;
 wire \V2/A2/A1/A1/M4/c2 ;
 wire \V2/A2/A1/A1/M4/s1 ;
 wire \V2/A2/A1/A2/c1 ;
 wire \V2/A2/A1/A2/c2 ;
 wire \V2/A2/A1/A2/c3 ;
 wire \V2/A2/A1/A2/M1/c1 ;
 wire \V2/A2/A1/A2/M1/c2 ;
 wire \V2/A2/A1/A2/M1/s1 ;
 wire \V2/A2/A1/A2/M2/c1 ;
 wire \V2/A2/A1/A2/M2/c2 ;
 wire \V2/A2/A1/A2/M2/s1 ;
 wire \V2/A2/A1/A2/M3/c1 ;
 wire \V2/A2/A1/A2/M3/c2 ;
 wire \V2/A2/A1/A2/M3/s1 ;
 wire \V2/A2/A1/A2/M4/c1 ;
 wire \V2/A2/A1/A2/M4/c2 ;
 wire \V2/A2/A1/A2/M4/s1 ;
 wire \V2/A2/A2/c1 ;
 wire \V2/A2/A2/A1/c1 ;
 wire \V2/A2/A2/A1/c2 ;
 wire \V2/A2/A2/A1/c3 ;
 wire \V2/A2/A2/A1/M1/c1 ;
 wire \V2/A2/A2/A1/M1/c2 ;
 wire \V2/A2/A2/A1/M1/s1 ;
 wire \V2/A2/A2/A1/M2/c1 ;
 wire \V2/A2/A2/A1/M2/c2 ;
 wire \V2/A2/A2/A1/M2/s1 ;
 wire \V2/A2/A2/A1/M3/c1 ;
 wire \V2/A2/A2/A1/M3/c2 ;
 wire \V2/A2/A2/A1/M3/s1 ;
 wire \V2/A2/A2/A1/M4/c1 ;
 wire \V2/A2/A2/A1/M4/c2 ;
 wire \V2/A2/A2/A1/M4/s1 ;
 wire \V2/A2/A2/A2/c1 ;
 wire \V2/A2/A2/A2/c2 ;
 wire \V2/A2/A2/A2/c3 ;
 wire \V2/A2/A2/A2/M1/c1 ;
 wire \V2/A2/A2/A2/M1/c2 ;
 wire \V2/A2/A2/A2/M1/s1 ;
 wire \V2/A2/A2/A2/M2/c1 ;
 wire \V2/A2/A2/A2/M2/c2 ;
 wire \V2/A2/A2/A2/M2/s1 ;
 wire \V2/A2/A2/A2/M3/c1 ;
 wire \V2/A2/A2/A2/M3/c2 ;
 wire \V2/A2/A2/A2/M3/s1 ;
 wire \V2/A2/A2/A2/M4/c1 ;
 wire \V2/A2/A2/A2/M4/c2 ;
 wire \V2/A2/A2/A2/M4/s1 ;
 wire \V2/A3/c1 ;
 wire \V2/A3/A1/c1 ;
 wire \V2/A3/A1/A1/c1 ;
 wire \V2/A3/A1/A1/c2 ;
 wire \V2/A3/A1/A1/c3 ;
 wire \V2/A3/A1/A1/M1/c1 ;
 wire \V2/A3/A1/A1/M1/c2 ;
 wire \V2/A3/A1/A1/M1/s1 ;
 wire \V2/A3/A1/A1/M2/c1 ;
 wire \V2/A3/A1/A1/M2/c2 ;
 wire \V2/A3/A1/A1/M2/s1 ;
 wire \V2/A3/A1/A1/M3/c1 ;
 wire \V2/A3/A1/A1/M3/c2 ;
 wire \V2/A3/A1/A1/M3/s1 ;
 wire \V2/A3/A1/A1/M4/c1 ;
 wire \V2/A3/A1/A1/M4/c2 ;
 wire \V2/A3/A1/A1/M4/s1 ;
 wire \V2/A3/A1/A2/c1 ;
 wire \V2/A3/A1/A2/c2 ;
 wire \V2/A3/A1/A2/c3 ;
 wire \V2/A3/A1/A2/M1/c1 ;
 wire \V2/A3/A1/A2/M1/c2 ;
 wire \V2/A3/A1/A2/M1/s1 ;
 wire \V2/A3/A1/A2/M2/c1 ;
 wire \V2/A3/A1/A2/M2/c2 ;
 wire \V2/A3/A1/A2/M2/s1 ;
 wire \V2/A3/A1/A2/M3/c1 ;
 wire \V2/A3/A1/A2/M3/c2 ;
 wire \V2/A3/A1/A2/M3/s1 ;
 wire \V2/A3/A1/A2/M4/c1 ;
 wire \V2/A3/A1/A2/M4/c2 ;
 wire \V2/A3/A1/A2/M4/s1 ;
 wire \V2/A3/A2/c1 ;
 wire \V2/A3/A2/A1/c1 ;
 wire \V2/A3/A2/A1/c2 ;
 wire \V2/A3/A2/A1/c3 ;
 wire \V2/A3/A2/A1/M1/c1 ;
 wire \V2/A3/A2/A1/M1/c2 ;
 wire \V2/A3/A2/A1/M1/s1 ;
 wire \V2/A3/A2/A1/M2/c1 ;
 wire \V2/A3/A2/A1/M2/c2 ;
 wire \V2/A3/A2/A1/M2/s1 ;
 wire \V2/A3/A2/A1/M3/c1 ;
 wire \V2/A3/A2/A1/M3/c2 ;
 wire \V2/A3/A2/A1/M3/s1 ;
 wire \V2/A3/A2/A1/M4/c1 ;
 wire \V2/A3/A2/A1/M4/c2 ;
 wire \V2/A3/A2/A1/M4/s1 ;
 wire \V2/A3/A2/A2/c1 ;
 wire \V2/A3/A2/A2/c2 ;
 wire \V2/A3/A2/A2/c3 ;
 wire \V2/A3/A2/A2/M1/c1 ;
 wire \V2/A3/A2/A2/M1/c2 ;
 wire \V2/A3/A2/A2/M1/s1 ;
 wire \V2/A3/A2/A2/M2/c1 ;
 wire \V2/A3/A2/A2/M2/c2 ;
 wire \V2/A3/A2/A2/M2/s1 ;
 wire \V2/A3/A2/A2/M3/c1 ;
 wire \V2/A3/A2/A2/M3/c2 ;
 wire \V2/A3/A2/A2/M3/s1 ;
 wire \V2/A3/A2/A2/M4/c1 ;
 wire \V2/A3/A2/A2/M4/c2 ;
 wire \V2/A3/A2/A2/M4/s1 ;
 wire \V2/V1/c1 ;
 wire \V2/V1/c2 ;
 wire \V2/V1/c3 ;
 wire \V2/V1/overflow ;
 wire \V2/V1/A1/c1 ;
 wire \V2/V1/A1/A1/c1 ;
 wire \V2/V1/A1/A1/c2 ;
 wire \V2/V1/A1/A1/c3 ;
 wire \V2/V1/A1/A1/M1/c1 ;
 wire \V2/V1/A1/A1/M1/c2 ;
 wire \V2/V1/A1/A1/M1/s1 ;
 wire \V2/V1/A1/A1/M2/c1 ;
 wire \V2/V1/A1/A1/M2/c2 ;
 wire \V2/V1/A1/A1/M2/s1 ;
 wire \V2/V1/A1/A1/M3/c1 ;
 wire \V2/V1/A1/A1/M3/c2 ;
 wire \V2/V1/A1/A1/M3/s1 ;
 wire \V2/V1/A1/A1/M4/c1 ;
 wire \V2/V1/A1/A1/M4/c2 ;
 wire \V2/V1/A1/A1/M4/s1 ;
 wire \V2/V1/A1/A2/c1 ;
 wire \V2/V1/A1/A2/c2 ;
 wire \V2/V1/A1/A2/c3 ;
 wire \V2/V1/A1/A2/M1/c1 ;
 wire \V2/V1/A1/A2/M1/c2 ;
 wire \V2/V1/A1/A2/M1/s1 ;
 wire \V2/V1/A1/A2/M2/c1 ;
 wire \V2/V1/A1/A2/M2/c2 ;
 wire \V2/V1/A1/A2/M2/s1 ;
 wire \V2/V1/A1/A2/M3/c1 ;
 wire \V2/V1/A1/A2/M3/c2 ;
 wire \V2/V1/A1/A2/M3/s1 ;
 wire \V2/V1/A1/A2/M4/c1 ;
 wire \V2/V1/A1/A2/M4/c2 ;
 wire \V2/V1/A1/A2/M4/s1 ;
 wire \V2/V1/A2/c1 ;
 wire \V2/V1/A2/A1/c1 ;
 wire \V2/V1/A2/A1/c2 ;
 wire \V2/V1/A2/A1/c3 ;
 wire \V2/V1/A2/A1/M1/c1 ;
 wire \V2/V1/A2/A1/M1/c2 ;
 wire \V2/V1/A2/A1/M1/s1 ;
 wire \V2/V1/A2/A1/M2/c1 ;
 wire \V2/V1/A2/A1/M2/c2 ;
 wire \V2/V1/A2/A1/M2/s1 ;
 wire \V2/V1/A2/A1/M3/c1 ;
 wire \V2/V1/A2/A1/M3/c2 ;
 wire \V2/V1/A2/A1/M3/s1 ;
 wire \V2/V1/A2/A1/M4/c1 ;
 wire \V2/V1/A2/A1/M4/c2 ;
 wire \V2/V1/A2/A1/M4/s1 ;
 wire \V2/V1/A2/A2/c1 ;
 wire \V2/V1/A2/A2/c2 ;
 wire \V2/V1/A2/A2/c3 ;
 wire \V2/V1/A2/A2/M1/c1 ;
 wire \V2/V1/A2/A2/M1/c2 ;
 wire \V2/V1/A2/A2/M1/s1 ;
 wire \V2/V1/A2/A2/M2/c1 ;
 wire \V2/V1/A2/A2/M2/c2 ;
 wire \V2/V1/A2/A2/M2/s1 ;
 wire \V2/V1/A2/A2/M3/c1 ;
 wire \V2/V1/A2/A2/M3/c2 ;
 wire \V2/V1/A2/A2/M3/s1 ;
 wire \V2/V1/A2/A2/M4/c1 ;
 wire \V2/V1/A2/A2/M4/c2 ;
 wire \V2/V1/A2/A2/M4/s1 ;
 wire \V2/V1/A3/c1 ;
 wire \V2/V1/A3/A1/c1 ;
 wire \V2/V1/A3/A1/c2 ;
 wire \V2/V1/A3/A1/c3 ;
 wire \V2/V1/A3/A1/M1/c1 ;
 wire \V2/V1/A3/A1/M1/c2 ;
 wire \V2/V1/A3/A1/M1/s1 ;
 wire \V2/V1/A3/A1/M2/c1 ;
 wire \V2/V1/A3/A1/M2/c2 ;
 wire \V2/V1/A3/A1/M2/s1 ;
 wire \V2/V1/A3/A1/M3/c1 ;
 wire \V2/V1/A3/A1/M3/c2 ;
 wire \V2/V1/A3/A1/M3/s1 ;
 wire \V2/V1/A3/A1/M4/c1 ;
 wire \V2/V1/A3/A1/M4/c2 ;
 wire \V2/V1/A3/A1/M4/s1 ;
 wire \V2/V1/A3/A2/c1 ;
 wire \V2/V1/A3/A2/c2 ;
 wire \V2/V1/A3/A2/c3 ;
 wire \V2/V1/A3/A2/M1/c1 ;
 wire \V2/V1/A3/A2/M1/c2 ;
 wire \V2/V1/A3/A2/M1/s1 ;
 wire \V2/V1/A3/A2/M2/c1 ;
 wire \V2/V1/A3/A2/M2/c2 ;
 wire \V2/V1/A3/A2/M2/s1 ;
 wire \V2/V1/A3/A2/M3/c1 ;
 wire \V2/V1/A3/A2/M3/c2 ;
 wire \V2/V1/A3/A2/M3/s1 ;
 wire \V2/V1/A3/A2/M4/c1 ;
 wire \V2/V1/A3/A2/M4/c2 ;
 wire \V2/V1/A3/A2/M4/s1 ;
 wire \V2/V1/V1/c1 ;
 wire \V2/V1/V1/c2 ;
 wire \V2/V1/V1/c3 ;
 wire \V2/V1/V1/overflow ;
 wire \V2/V1/V1/A1/c1 ;
 wire \V2/V1/V1/A1/c2 ;
 wire \V2/V1/V1/A1/c3 ;
 wire \V2/V1/V1/A1/M1/c1 ;
 wire \V2/V1/V1/A1/M1/c2 ;
 wire \V2/V1/V1/A1/M1/s1 ;
 wire \V2/V1/V1/A1/M2/c1 ;
 wire \V2/V1/V1/A1/M2/c2 ;
 wire \V2/V1/V1/A1/M2/s1 ;
 wire \V2/V1/V1/A1/M3/c1 ;
 wire \V2/V1/V1/A1/M3/c2 ;
 wire \V2/V1/V1/A1/M3/s1 ;
 wire \V2/V1/V1/A1/M4/c1 ;
 wire \V2/V1/V1/A1/M4/c2 ;
 wire \V2/V1/V1/A1/M4/s1 ;
 wire \V2/V1/V1/A2/c1 ;
 wire \V2/V1/V1/A2/c2 ;
 wire \V2/V1/V1/A2/c3 ;
 wire \V2/V1/V1/A2/M1/c1 ;
 wire \V2/V1/V1/A2/M1/c2 ;
 wire \V2/V1/V1/A2/M1/s1 ;
 wire \V2/V1/V1/A2/M2/c1 ;
 wire \V2/V1/V1/A2/M2/c2 ;
 wire \V2/V1/V1/A2/M2/s1 ;
 wire \V2/V1/V1/A2/M3/c1 ;
 wire \V2/V1/V1/A2/M3/c2 ;
 wire \V2/V1/V1/A2/M3/s1 ;
 wire \V2/V1/V1/A2/M4/c1 ;
 wire \V2/V1/V1/A2/M4/c2 ;
 wire \V2/V1/V1/A2/M4/s1 ;
 wire \V2/V1/V1/A3/c1 ;
 wire \V2/V1/V1/A3/c2 ;
 wire \V2/V1/V1/A3/c3 ;
 wire \V2/V1/V1/A3/M1/c1 ;
 wire \V2/V1/V1/A3/M1/c2 ;
 wire \V2/V1/V1/A3/M1/s1 ;
 wire \V2/V1/V1/A3/M2/c1 ;
 wire \V2/V1/V1/A3/M2/c2 ;
 wire \V2/V1/V1/A3/M2/s1 ;
 wire \V2/V1/V1/A3/M3/c1 ;
 wire \V2/V1/V1/A3/M3/c2 ;
 wire \V2/V1/V1/A3/M3/s1 ;
 wire \V2/V1/V1/A3/M4/c1 ;
 wire \V2/V1/V1/A3/M4/c2 ;
 wire \V2/V1/V1/A3/M4/s1 ;
 wire \V2/V1/V1/V1/w1 ;
 wire \V2/V1/V1/V1/w2 ;
 wire \V2/V1/V1/V1/w3 ;
 wire \V2/V1/V1/V1/w4 ;
 wire \V2/V1/V1/V2/w1 ;
 wire \V2/V1/V1/V2/w2 ;
 wire \V2/V1/V1/V2/w3 ;
 wire \V2/V1/V1/V2/w4 ;
 wire \V2/V1/V1/V3/w1 ;
 wire \V2/V1/V1/V3/w2 ;
 wire \V2/V1/V1/V3/w3 ;
 wire \V2/V1/V1/V3/w4 ;
 wire \V2/V1/V1/V4/w1 ;
 wire \V2/V1/V1/V4/w2 ;
 wire \V2/V1/V1/V4/w3 ;
 wire \V2/V1/V1/V4/w4 ;
 wire \V2/V1/V2/c1 ;
 wire \V2/V1/V2/c2 ;
 wire \V2/V1/V2/c3 ;
 wire \V2/V1/V2/overflow ;
 wire \V2/V1/V2/A1/c1 ;
 wire \V2/V1/V2/A1/c2 ;
 wire \V2/V1/V2/A1/c3 ;
 wire \V2/V1/V2/A1/M1/c1 ;
 wire \V2/V1/V2/A1/M1/c2 ;
 wire \V2/V1/V2/A1/M1/s1 ;
 wire \V2/V1/V2/A1/M2/c1 ;
 wire \V2/V1/V2/A1/M2/c2 ;
 wire \V2/V1/V2/A1/M2/s1 ;
 wire \V2/V1/V2/A1/M3/c1 ;
 wire \V2/V1/V2/A1/M3/c2 ;
 wire \V2/V1/V2/A1/M3/s1 ;
 wire \V2/V1/V2/A1/M4/c1 ;
 wire \V2/V1/V2/A1/M4/c2 ;
 wire \V2/V1/V2/A1/M4/s1 ;
 wire \V2/V1/V2/A2/c1 ;
 wire \V2/V1/V2/A2/c2 ;
 wire \V2/V1/V2/A2/c3 ;
 wire \V2/V1/V2/A2/M1/c1 ;
 wire \V2/V1/V2/A2/M1/c2 ;
 wire \V2/V1/V2/A2/M1/s1 ;
 wire \V2/V1/V2/A2/M2/c1 ;
 wire \V2/V1/V2/A2/M2/c2 ;
 wire \V2/V1/V2/A2/M2/s1 ;
 wire \V2/V1/V2/A2/M3/c1 ;
 wire \V2/V1/V2/A2/M3/c2 ;
 wire \V2/V1/V2/A2/M3/s1 ;
 wire \V2/V1/V2/A2/M4/c1 ;
 wire \V2/V1/V2/A2/M4/c2 ;
 wire \V2/V1/V2/A2/M4/s1 ;
 wire \V2/V1/V2/A3/c1 ;
 wire \V2/V1/V2/A3/c2 ;
 wire \V2/V1/V2/A3/c3 ;
 wire \V2/V1/V2/A3/M1/c1 ;
 wire \V2/V1/V2/A3/M1/c2 ;
 wire \V2/V1/V2/A3/M1/s1 ;
 wire \V2/V1/V2/A3/M2/c1 ;
 wire \V2/V1/V2/A3/M2/c2 ;
 wire \V2/V1/V2/A3/M2/s1 ;
 wire \V2/V1/V2/A3/M3/c1 ;
 wire \V2/V1/V2/A3/M3/c2 ;
 wire \V2/V1/V2/A3/M3/s1 ;
 wire \V2/V1/V2/A3/M4/c1 ;
 wire \V2/V1/V2/A3/M4/c2 ;
 wire \V2/V1/V2/A3/M4/s1 ;
 wire \V2/V1/V2/V1/w1 ;
 wire \V2/V1/V2/V1/w2 ;
 wire \V2/V1/V2/V1/w3 ;
 wire \V2/V1/V2/V1/w4 ;
 wire \V2/V1/V2/V2/w1 ;
 wire \V2/V1/V2/V2/w2 ;
 wire \V2/V1/V2/V2/w3 ;
 wire \V2/V1/V2/V2/w4 ;
 wire \V2/V1/V2/V3/w1 ;
 wire \V2/V1/V2/V3/w2 ;
 wire \V2/V1/V2/V3/w3 ;
 wire \V2/V1/V2/V3/w4 ;
 wire \V2/V1/V2/V4/w1 ;
 wire \V2/V1/V2/V4/w2 ;
 wire \V2/V1/V2/V4/w3 ;
 wire \V2/V1/V2/V4/w4 ;
 wire \V2/V1/V3/c1 ;
 wire \V2/V1/V3/c2 ;
 wire \V2/V1/V3/c3 ;
 wire \V2/V1/V3/overflow ;
 wire \V2/V1/V3/A1/c1 ;
 wire \V2/V1/V3/A1/c2 ;
 wire \V2/V1/V3/A1/c3 ;
 wire \V2/V1/V3/A1/M1/c1 ;
 wire \V2/V1/V3/A1/M1/c2 ;
 wire \V2/V1/V3/A1/M1/s1 ;
 wire \V2/V1/V3/A1/M2/c1 ;
 wire \V2/V1/V3/A1/M2/c2 ;
 wire \V2/V1/V3/A1/M2/s1 ;
 wire \V2/V1/V3/A1/M3/c1 ;
 wire \V2/V1/V3/A1/M3/c2 ;
 wire \V2/V1/V3/A1/M3/s1 ;
 wire \V2/V1/V3/A1/M4/c1 ;
 wire \V2/V1/V3/A1/M4/c2 ;
 wire \V2/V1/V3/A1/M4/s1 ;
 wire \V2/V1/V3/A2/c1 ;
 wire \V2/V1/V3/A2/c2 ;
 wire \V2/V1/V3/A2/c3 ;
 wire \V2/V1/V3/A2/M1/c1 ;
 wire \V2/V1/V3/A2/M1/c2 ;
 wire \V2/V1/V3/A2/M1/s1 ;
 wire \V2/V1/V3/A2/M2/c1 ;
 wire \V2/V1/V3/A2/M2/c2 ;
 wire \V2/V1/V3/A2/M2/s1 ;
 wire \V2/V1/V3/A2/M3/c1 ;
 wire \V2/V1/V3/A2/M3/c2 ;
 wire \V2/V1/V3/A2/M3/s1 ;
 wire \V2/V1/V3/A2/M4/c1 ;
 wire \V2/V1/V3/A2/M4/c2 ;
 wire \V2/V1/V3/A2/M4/s1 ;
 wire \V2/V1/V3/A3/c1 ;
 wire \V2/V1/V3/A3/c2 ;
 wire \V2/V1/V3/A3/c3 ;
 wire \V2/V1/V3/A3/M1/c1 ;
 wire \V2/V1/V3/A3/M1/c2 ;
 wire \V2/V1/V3/A3/M1/s1 ;
 wire \V2/V1/V3/A3/M2/c1 ;
 wire \V2/V1/V3/A3/M2/c2 ;
 wire \V2/V1/V3/A3/M2/s1 ;
 wire \V2/V1/V3/A3/M3/c1 ;
 wire \V2/V1/V3/A3/M3/c2 ;
 wire \V2/V1/V3/A3/M3/s1 ;
 wire \V2/V1/V3/A3/M4/c1 ;
 wire \V2/V1/V3/A3/M4/c2 ;
 wire \V2/V1/V3/A3/M4/s1 ;
 wire \V2/V1/V3/V1/w1 ;
 wire \V2/V1/V3/V1/w2 ;
 wire \V2/V1/V3/V1/w3 ;
 wire \V2/V1/V3/V1/w4 ;
 wire \V2/V1/V3/V2/w1 ;
 wire \V2/V1/V3/V2/w2 ;
 wire \V2/V1/V3/V2/w3 ;
 wire \V2/V1/V3/V2/w4 ;
 wire \V2/V1/V3/V3/w1 ;
 wire \V2/V1/V3/V3/w2 ;
 wire \V2/V1/V3/V3/w3 ;
 wire \V2/V1/V3/V3/w4 ;
 wire \V2/V1/V3/V4/w1 ;
 wire \V2/V1/V3/V4/w2 ;
 wire \V2/V1/V3/V4/w3 ;
 wire \V2/V1/V3/V4/w4 ;
 wire \V2/V1/V4/c1 ;
 wire \V2/V1/V4/c2 ;
 wire \V2/V1/V4/c3 ;
 wire \V2/V1/V4/overflow ;
 wire \V2/V1/V4/A1/c1 ;
 wire \V2/V1/V4/A1/c2 ;
 wire \V2/V1/V4/A1/c3 ;
 wire \V2/V1/V4/A1/M1/c1 ;
 wire \V2/V1/V4/A1/M1/c2 ;
 wire \V2/V1/V4/A1/M1/s1 ;
 wire \V2/V1/V4/A1/M2/c1 ;
 wire \V2/V1/V4/A1/M2/c2 ;
 wire \V2/V1/V4/A1/M2/s1 ;
 wire \V2/V1/V4/A1/M3/c1 ;
 wire \V2/V1/V4/A1/M3/c2 ;
 wire \V2/V1/V4/A1/M3/s1 ;
 wire \V2/V1/V4/A1/M4/c1 ;
 wire \V2/V1/V4/A1/M4/c2 ;
 wire \V2/V1/V4/A1/M4/s1 ;
 wire \V2/V1/V4/A2/c1 ;
 wire \V2/V1/V4/A2/c2 ;
 wire \V2/V1/V4/A2/c3 ;
 wire \V2/V1/V4/A2/M1/c1 ;
 wire \V2/V1/V4/A2/M1/c2 ;
 wire \V2/V1/V4/A2/M1/s1 ;
 wire \V2/V1/V4/A2/M2/c1 ;
 wire \V2/V1/V4/A2/M2/c2 ;
 wire \V2/V1/V4/A2/M2/s1 ;
 wire \V2/V1/V4/A2/M3/c1 ;
 wire \V2/V1/V4/A2/M3/c2 ;
 wire \V2/V1/V4/A2/M3/s1 ;
 wire \V2/V1/V4/A2/M4/c1 ;
 wire \V2/V1/V4/A2/M4/c2 ;
 wire \V2/V1/V4/A2/M4/s1 ;
 wire \V2/V1/V4/A3/c1 ;
 wire \V2/V1/V4/A3/c2 ;
 wire \V2/V1/V4/A3/c3 ;
 wire \V2/V1/V4/A3/M1/c1 ;
 wire \V2/V1/V4/A3/M1/c2 ;
 wire \V2/V1/V4/A3/M1/s1 ;
 wire \V2/V1/V4/A3/M2/c1 ;
 wire \V2/V1/V4/A3/M2/c2 ;
 wire \V2/V1/V4/A3/M2/s1 ;
 wire \V2/V1/V4/A3/M3/c1 ;
 wire \V2/V1/V4/A3/M3/c2 ;
 wire \V2/V1/V4/A3/M3/s1 ;
 wire \V2/V1/V4/A3/M4/c1 ;
 wire \V2/V1/V4/A3/M4/c2 ;
 wire \V2/V1/V4/A3/M4/s1 ;
 wire \V2/V1/V4/V1/w1 ;
 wire \V2/V1/V4/V1/w2 ;
 wire \V2/V1/V4/V1/w3 ;
 wire \V2/V1/V4/V1/w4 ;
 wire \V2/V1/V4/V2/w1 ;
 wire \V2/V1/V4/V2/w2 ;
 wire \V2/V1/V4/V2/w3 ;
 wire \V2/V1/V4/V2/w4 ;
 wire \V2/V1/V4/V3/w1 ;
 wire \V2/V1/V4/V3/w2 ;
 wire \V2/V1/V4/V3/w3 ;
 wire \V2/V1/V4/V3/w4 ;
 wire \V2/V1/V4/V4/w1 ;
 wire \V2/V1/V4/V4/w2 ;
 wire \V2/V1/V4/V4/w3 ;
 wire \V2/V1/V4/V4/w4 ;
 wire \V2/V2/c1 ;
 wire \V2/V2/c2 ;
 wire \V2/V2/c3 ;
 wire \V2/V2/overflow ;
 wire \V2/V2/A1/c1 ;
 wire \V2/V2/A1/A1/c1 ;
 wire \V2/V2/A1/A1/c2 ;
 wire \V2/V2/A1/A1/c3 ;
 wire \V2/V2/A1/A1/M1/c1 ;
 wire \V2/V2/A1/A1/M1/c2 ;
 wire \V2/V2/A1/A1/M1/s1 ;
 wire \V2/V2/A1/A1/M2/c1 ;
 wire \V2/V2/A1/A1/M2/c2 ;
 wire \V2/V2/A1/A1/M2/s1 ;
 wire \V2/V2/A1/A1/M3/c1 ;
 wire \V2/V2/A1/A1/M3/c2 ;
 wire \V2/V2/A1/A1/M3/s1 ;
 wire \V2/V2/A1/A1/M4/c1 ;
 wire \V2/V2/A1/A1/M4/c2 ;
 wire \V2/V2/A1/A1/M4/s1 ;
 wire \V2/V2/A1/A2/c1 ;
 wire \V2/V2/A1/A2/c2 ;
 wire \V2/V2/A1/A2/c3 ;
 wire \V2/V2/A1/A2/M1/c1 ;
 wire \V2/V2/A1/A2/M1/c2 ;
 wire \V2/V2/A1/A2/M1/s1 ;
 wire \V2/V2/A1/A2/M2/c1 ;
 wire \V2/V2/A1/A2/M2/c2 ;
 wire \V2/V2/A1/A2/M2/s1 ;
 wire \V2/V2/A1/A2/M3/c1 ;
 wire \V2/V2/A1/A2/M3/c2 ;
 wire \V2/V2/A1/A2/M3/s1 ;
 wire \V2/V2/A1/A2/M4/c1 ;
 wire \V2/V2/A1/A2/M4/c2 ;
 wire \V2/V2/A1/A2/M4/s1 ;
 wire \V2/V2/A2/c1 ;
 wire \V2/V2/A2/A1/c1 ;
 wire \V2/V2/A2/A1/c2 ;
 wire \V2/V2/A2/A1/c3 ;
 wire \V2/V2/A2/A1/M1/c1 ;
 wire \V2/V2/A2/A1/M1/c2 ;
 wire \V2/V2/A2/A1/M1/s1 ;
 wire \V2/V2/A2/A1/M2/c1 ;
 wire \V2/V2/A2/A1/M2/c2 ;
 wire \V2/V2/A2/A1/M2/s1 ;
 wire \V2/V2/A2/A1/M3/c1 ;
 wire \V2/V2/A2/A1/M3/c2 ;
 wire \V2/V2/A2/A1/M3/s1 ;
 wire \V2/V2/A2/A1/M4/c1 ;
 wire \V2/V2/A2/A1/M4/c2 ;
 wire \V2/V2/A2/A1/M4/s1 ;
 wire \V2/V2/A2/A2/c1 ;
 wire \V2/V2/A2/A2/c2 ;
 wire \V2/V2/A2/A2/c3 ;
 wire \V2/V2/A2/A2/M1/c1 ;
 wire \V2/V2/A2/A2/M1/c2 ;
 wire \V2/V2/A2/A2/M1/s1 ;
 wire \V2/V2/A2/A2/M2/c1 ;
 wire \V2/V2/A2/A2/M2/c2 ;
 wire \V2/V2/A2/A2/M2/s1 ;
 wire \V2/V2/A2/A2/M3/c1 ;
 wire \V2/V2/A2/A2/M3/c2 ;
 wire \V2/V2/A2/A2/M3/s1 ;
 wire \V2/V2/A2/A2/M4/c1 ;
 wire \V2/V2/A2/A2/M4/c2 ;
 wire \V2/V2/A2/A2/M4/s1 ;
 wire \V2/V2/A3/c1 ;
 wire \V2/V2/A3/A1/c1 ;
 wire \V2/V2/A3/A1/c2 ;
 wire \V2/V2/A3/A1/c3 ;
 wire \V2/V2/A3/A1/M1/c1 ;
 wire \V2/V2/A3/A1/M1/c2 ;
 wire \V2/V2/A3/A1/M1/s1 ;
 wire \V2/V2/A3/A1/M2/c1 ;
 wire \V2/V2/A3/A1/M2/c2 ;
 wire \V2/V2/A3/A1/M2/s1 ;
 wire \V2/V2/A3/A1/M3/c1 ;
 wire \V2/V2/A3/A1/M3/c2 ;
 wire \V2/V2/A3/A1/M3/s1 ;
 wire \V2/V2/A3/A1/M4/c1 ;
 wire \V2/V2/A3/A1/M4/c2 ;
 wire \V2/V2/A3/A1/M4/s1 ;
 wire \V2/V2/A3/A2/c1 ;
 wire \V2/V2/A3/A2/c2 ;
 wire \V2/V2/A3/A2/c3 ;
 wire \V2/V2/A3/A2/M1/c1 ;
 wire \V2/V2/A3/A2/M1/c2 ;
 wire \V2/V2/A3/A2/M1/s1 ;
 wire \V2/V2/A3/A2/M2/c1 ;
 wire \V2/V2/A3/A2/M2/c2 ;
 wire \V2/V2/A3/A2/M2/s1 ;
 wire \V2/V2/A3/A2/M3/c1 ;
 wire \V2/V2/A3/A2/M3/c2 ;
 wire \V2/V2/A3/A2/M3/s1 ;
 wire \V2/V2/A3/A2/M4/c1 ;
 wire \V2/V2/A3/A2/M4/c2 ;
 wire \V2/V2/A3/A2/M4/s1 ;
 wire \V2/V2/V1/c1 ;
 wire \V2/V2/V1/c2 ;
 wire \V2/V2/V1/c3 ;
 wire \V2/V2/V1/overflow ;
 wire \V2/V2/V1/A1/c1 ;
 wire \V2/V2/V1/A1/c2 ;
 wire \V2/V2/V1/A1/c3 ;
 wire \V2/V2/V1/A1/M1/c1 ;
 wire \V2/V2/V1/A1/M1/c2 ;
 wire \V2/V2/V1/A1/M1/s1 ;
 wire \V2/V2/V1/A1/M2/c1 ;
 wire \V2/V2/V1/A1/M2/c2 ;
 wire \V2/V2/V1/A1/M2/s1 ;
 wire \V2/V2/V1/A1/M3/c1 ;
 wire \V2/V2/V1/A1/M3/c2 ;
 wire \V2/V2/V1/A1/M3/s1 ;
 wire \V2/V2/V1/A1/M4/c1 ;
 wire \V2/V2/V1/A1/M4/c2 ;
 wire \V2/V2/V1/A1/M4/s1 ;
 wire \V2/V2/V1/A2/c1 ;
 wire \V2/V2/V1/A2/c2 ;
 wire \V2/V2/V1/A2/c3 ;
 wire \V2/V2/V1/A2/M1/c1 ;
 wire \V2/V2/V1/A2/M1/c2 ;
 wire \V2/V2/V1/A2/M1/s1 ;
 wire \V2/V2/V1/A2/M2/c1 ;
 wire \V2/V2/V1/A2/M2/c2 ;
 wire \V2/V2/V1/A2/M2/s1 ;
 wire \V2/V2/V1/A2/M3/c1 ;
 wire \V2/V2/V1/A2/M3/c2 ;
 wire \V2/V2/V1/A2/M3/s1 ;
 wire \V2/V2/V1/A2/M4/c1 ;
 wire \V2/V2/V1/A2/M4/c2 ;
 wire \V2/V2/V1/A2/M4/s1 ;
 wire \V2/V2/V1/A3/c1 ;
 wire \V2/V2/V1/A3/c2 ;
 wire \V2/V2/V1/A3/c3 ;
 wire \V2/V2/V1/A3/M1/c1 ;
 wire \V2/V2/V1/A3/M1/c2 ;
 wire \V2/V2/V1/A3/M1/s1 ;
 wire \V2/V2/V1/A3/M2/c1 ;
 wire \V2/V2/V1/A3/M2/c2 ;
 wire \V2/V2/V1/A3/M2/s1 ;
 wire \V2/V2/V1/A3/M3/c1 ;
 wire \V2/V2/V1/A3/M3/c2 ;
 wire \V2/V2/V1/A3/M3/s1 ;
 wire \V2/V2/V1/A3/M4/c1 ;
 wire \V2/V2/V1/A3/M4/c2 ;
 wire \V2/V2/V1/A3/M4/s1 ;
 wire \V2/V2/V1/V1/w1 ;
 wire \V2/V2/V1/V1/w2 ;
 wire \V2/V2/V1/V1/w3 ;
 wire \V2/V2/V1/V1/w4 ;
 wire \V2/V2/V1/V2/w1 ;
 wire \V2/V2/V1/V2/w2 ;
 wire \V2/V2/V1/V2/w3 ;
 wire \V2/V2/V1/V2/w4 ;
 wire \V2/V2/V1/V3/w1 ;
 wire \V2/V2/V1/V3/w2 ;
 wire \V2/V2/V1/V3/w3 ;
 wire \V2/V2/V1/V3/w4 ;
 wire \V2/V2/V1/V4/w1 ;
 wire \V2/V2/V1/V4/w2 ;
 wire \V2/V2/V1/V4/w3 ;
 wire \V2/V2/V1/V4/w4 ;
 wire \V2/V2/V2/c1 ;
 wire \V2/V2/V2/c2 ;
 wire \V2/V2/V2/c3 ;
 wire \V2/V2/V2/overflow ;
 wire \V2/V2/V2/A1/c1 ;
 wire \V2/V2/V2/A1/c2 ;
 wire \V2/V2/V2/A1/c3 ;
 wire \V2/V2/V2/A1/M1/c1 ;
 wire \V2/V2/V2/A1/M1/c2 ;
 wire \V2/V2/V2/A1/M1/s1 ;
 wire \V2/V2/V2/A1/M2/c1 ;
 wire \V2/V2/V2/A1/M2/c2 ;
 wire \V2/V2/V2/A1/M2/s1 ;
 wire \V2/V2/V2/A1/M3/c1 ;
 wire \V2/V2/V2/A1/M3/c2 ;
 wire \V2/V2/V2/A1/M3/s1 ;
 wire \V2/V2/V2/A1/M4/c1 ;
 wire \V2/V2/V2/A1/M4/c2 ;
 wire \V2/V2/V2/A1/M4/s1 ;
 wire \V2/V2/V2/A2/c1 ;
 wire \V2/V2/V2/A2/c2 ;
 wire \V2/V2/V2/A2/c3 ;
 wire \V2/V2/V2/A2/M1/c1 ;
 wire \V2/V2/V2/A2/M1/c2 ;
 wire \V2/V2/V2/A2/M1/s1 ;
 wire \V2/V2/V2/A2/M2/c1 ;
 wire \V2/V2/V2/A2/M2/c2 ;
 wire \V2/V2/V2/A2/M2/s1 ;
 wire \V2/V2/V2/A2/M3/c1 ;
 wire \V2/V2/V2/A2/M3/c2 ;
 wire \V2/V2/V2/A2/M3/s1 ;
 wire \V2/V2/V2/A2/M4/c1 ;
 wire \V2/V2/V2/A2/M4/c2 ;
 wire \V2/V2/V2/A2/M4/s1 ;
 wire \V2/V2/V2/A3/c1 ;
 wire \V2/V2/V2/A3/c2 ;
 wire \V2/V2/V2/A3/c3 ;
 wire \V2/V2/V2/A3/M1/c1 ;
 wire \V2/V2/V2/A3/M1/c2 ;
 wire \V2/V2/V2/A3/M1/s1 ;
 wire \V2/V2/V2/A3/M2/c1 ;
 wire \V2/V2/V2/A3/M2/c2 ;
 wire \V2/V2/V2/A3/M2/s1 ;
 wire \V2/V2/V2/A3/M3/c1 ;
 wire \V2/V2/V2/A3/M3/c2 ;
 wire \V2/V2/V2/A3/M3/s1 ;
 wire \V2/V2/V2/A3/M4/c1 ;
 wire \V2/V2/V2/A3/M4/c2 ;
 wire \V2/V2/V2/A3/M4/s1 ;
 wire \V2/V2/V2/V1/w1 ;
 wire \V2/V2/V2/V1/w2 ;
 wire \V2/V2/V2/V1/w3 ;
 wire \V2/V2/V2/V1/w4 ;
 wire \V2/V2/V2/V2/w1 ;
 wire \V2/V2/V2/V2/w2 ;
 wire \V2/V2/V2/V2/w3 ;
 wire \V2/V2/V2/V2/w4 ;
 wire \V2/V2/V2/V3/w1 ;
 wire \V2/V2/V2/V3/w2 ;
 wire \V2/V2/V2/V3/w3 ;
 wire \V2/V2/V2/V3/w4 ;
 wire \V2/V2/V2/V4/w1 ;
 wire \V2/V2/V2/V4/w2 ;
 wire \V2/V2/V2/V4/w3 ;
 wire \V2/V2/V2/V4/w4 ;
 wire \V2/V2/V3/c1 ;
 wire \V2/V2/V3/c2 ;
 wire \V2/V2/V3/c3 ;
 wire \V2/V2/V3/overflow ;
 wire \V2/V2/V3/A1/c1 ;
 wire \V2/V2/V3/A1/c2 ;
 wire \V2/V2/V3/A1/c3 ;
 wire \V2/V2/V3/A1/M1/c1 ;
 wire \V2/V2/V3/A1/M1/c2 ;
 wire \V2/V2/V3/A1/M1/s1 ;
 wire \V2/V2/V3/A1/M2/c1 ;
 wire \V2/V2/V3/A1/M2/c2 ;
 wire \V2/V2/V3/A1/M2/s1 ;
 wire \V2/V2/V3/A1/M3/c1 ;
 wire \V2/V2/V3/A1/M3/c2 ;
 wire \V2/V2/V3/A1/M3/s1 ;
 wire \V2/V2/V3/A1/M4/c1 ;
 wire \V2/V2/V3/A1/M4/c2 ;
 wire \V2/V2/V3/A1/M4/s1 ;
 wire \V2/V2/V3/A2/c1 ;
 wire \V2/V2/V3/A2/c2 ;
 wire \V2/V2/V3/A2/c3 ;
 wire \V2/V2/V3/A2/M1/c1 ;
 wire \V2/V2/V3/A2/M1/c2 ;
 wire \V2/V2/V3/A2/M1/s1 ;
 wire \V2/V2/V3/A2/M2/c1 ;
 wire \V2/V2/V3/A2/M2/c2 ;
 wire \V2/V2/V3/A2/M2/s1 ;
 wire \V2/V2/V3/A2/M3/c1 ;
 wire \V2/V2/V3/A2/M3/c2 ;
 wire \V2/V2/V3/A2/M3/s1 ;
 wire \V2/V2/V3/A2/M4/c1 ;
 wire \V2/V2/V3/A2/M4/c2 ;
 wire \V2/V2/V3/A2/M4/s1 ;
 wire \V2/V2/V3/A3/c1 ;
 wire \V2/V2/V3/A3/c2 ;
 wire \V2/V2/V3/A3/c3 ;
 wire \V2/V2/V3/A3/M1/c1 ;
 wire \V2/V2/V3/A3/M1/c2 ;
 wire \V2/V2/V3/A3/M1/s1 ;
 wire \V2/V2/V3/A3/M2/c1 ;
 wire \V2/V2/V3/A3/M2/c2 ;
 wire \V2/V2/V3/A3/M2/s1 ;
 wire \V2/V2/V3/A3/M3/c1 ;
 wire \V2/V2/V3/A3/M3/c2 ;
 wire \V2/V2/V3/A3/M3/s1 ;
 wire \V2/V2/V3/A3/M4/c1 ;
 wire \V2/V2/V3/A3/M4/c2 ;
 wire \V2/V2/V3/A3/M4/s1 ;
 wire \V2/V2/V3/V1/w1 ;
 wire \V2/V2/V3/V1/w2 ;
 wire \V2/V2/V3/V1/w3 ;
 wire \V2/V2/V3/V1/w4 ;
 wire \V2/V2/V3/V2/w1 ;
 wire \V2/V2/V3/V2/w2 ;
 wire \V2/V2/V3/V2/w3 ;
 wire \V2/V2/V3/V2/w4 ;
 wire \V2/V2/V3/V3/w1 ;
 wire \V2/V2/V3/V3/w2 ;
 wire \V2/V2/V3/V3/w3 ;
 wire \V2/V2/V3/V3/w4 ;
 wire \V2/V2/V3/V4/w1 ;
 wire \V2/V2/V3/V4/w2 ;
 wire \V2/V2/V3/V4/w3 ;
 wire \V2/V2/V3/V4/w4 ;
 wire \V2/V2/V4/c1 ;
 wire \V2/V2/V4/c2 ;
 wire \V2/V2/V4/c3 ;
 wire \V2/V2/V4/overflow ;
 wire \V2/V2/V4/A1/c1 ;
 wire \V2/V2/V4/A1/c2 ;
 wire \V2/V2/V4/A1/c3 ;
 wire \V2/V2/V4/A1/M1/c1 ;
 wire \V2/V2/V4/A1/M1/c2 ;
 wire \V2/V2/V4/A1/M1/s1 ;
 wire \V2/V2/V4/A1/M2/c1 ;
 wire \V2/V2/V4/A1/M2/c2 ;
 wire \V2/V2/V4/A1/M2/s1 ;
 wire \V2/V2/V4/A1/M3/c1 ;
 wire \V2/V2/V4/A1/M3/c2 ;
 wire \V2/V2/V4/A1/M3/s1 ;
 wire \V2/V2/V4/A1/M4/c1 ;
 wire \V2/V2/V4/A1/M4/c2 ;
 wire \V2/V2/V4/A1/M4/s1 ;
 wire \V2/V2/V4/A2/c1 ;
 wire \V2/V2/V4/A2/c2 ;
 wire \V2/V2/V4/A2/c3 ;
 wire \V2/V2/V4/A2/M1/c1 ;
 wire \V2/V2/V4/A2/M1/c2 ;
 wire \V2/V2/V4/A2/M1/s1 ;
 wire \V2/V2/V4/A2/M2/c1 ;
 wire \V2/V2/V4/A2/M2/c2 ;
 wire \V2/V2/V4/A2/M2/s1 ;
 wire \V2/V2/V4/A2/M3/c1 ;
 wire \V2/V2/V4/A2/M3/c2 ;
 wire \V2/V2/V4/A2/M3/s1 ;
 wire \V2/V2/V4/A2/M4/c1 ;
 wire \V2/V2/V4/A2/M4/c2 ;
 wire \V2/V2/V4/A2/M4/s1 ;
 wire \V2/V2/V4/A3/c1 ;
 wire \V2/V2/V4/A3/c2 ;
 wire \V2/V2/V4/A3/c3 ;
 wire \V2/V2/V4/A3/M1/c1 ;
 wire \V2/V2/V4/A3/M1/c2 ;
 wire \V2/V2/V4/A3/M1/s1 ;
 wire \V2/V2/V4/A3/M2/c1 ;
 wire \V2/V2/V4/A3/M2/c2 ;
 wire \V2/V2/V4/A3/M2/s1 ;
 wire \V2/V2/V4/A3/M3/c1 ;
 wire \V2/V2/V4/A3/M3/c2 ;
 wire \V2/V2/V4/A3/M3/s1 ;
 wire \V2/V2/V4/A3/M4/c1 ;
 wire \V2/V2/V4/A3/M4/c2 ;
 wire \V2/V2/V4/A3/M4/s1 ;
 wire \V2/V2/V4/V1/w1 ;
 wire \V2/V2/V4/V1/w2 ;
 wire \V2/V2/V4/V1/w3 ;
 wire \V2/V2/V4/V1/w4 ;
 wire \V2/V2/V4/V2/w1 ;
 wire \V2/V2/V4/V2/w2 ;
 wire \V2/V2/V4/V2/w3 ;
 wire \V2/V2/V4/V2/w4 ;
 wire \V2/V2/V4/V3/w1 ;
 wire \V2/V2/V4/V3/w2 ;
 wire \V2/V2/V4/V3/w3 ;
 wire \V2/V2/V4/V3/w4 ;
 wire \V2/V2/V4/V4/w1 ;
 wire \V2/V2/V4/V4/w2 ;
 wire \V2/V2/V4/V4/w3 ;
 wire \V2/V2/V4/V4/w4 ;
 wire \V2/V3/c1 ;
 wire \V2/V3/c2 ;
 wire \V2/V3/c3 ;
 wire \V2/V3/overflow ;
 wire \V2/V3/A1/c1 ;
 wire \V2/V3/A1/A1/c1 ;
 wire \V2/V3/A1/A1/c2 ;
 wire \V2/V3/A1/A1/c3 ;
 wire \V2/V3/A1/A1/M1/c1 ;
 wire \V2/V3/A1/A1/M1/c2 ;
 wire \V2/V3/A1/A1/M1/s1 ;
 wire \V2/V3/A1/A1/M2/c1 ;
 wire \V2/V3/A1/A1/M2/c2 ;
 wire \V2/V3/A1/A1/M2/s1 ;
 wire \V2/V3/A1/A1/M3/c1 ;
 wire \V2/V3/A1/A1/M3/c2 ;
 wire \V2/V3/A1/A1/M3/s1 ;
 wire \V2/V3/A1/A1/M4/c1 ;
 wire \V2/V3/A1/A1/M4/c2 ;
 wire \V2/V3/A1/A1/M4/s1 ;
 wire \V2/V3/A1/A2/c1 ;
 wire \V2/V3/A1/A2/c2 ;
 wire \V2/V3/A1/A2/c3 ;
 wire \V2/V3/A1/A2/M1/c1 ;
 wire \V2/V3/A1/A2/M1/c2 ;
 wire \V2/V3/A1/A2/M1/s1 ;
 wire \V2/V3/A1/A2/M2/c1 ;
 wire \V2/V3/A1/A2/M2/c2 ;
 wire \V2/V3/A1/A2/M2/s1 ;
 wire \V2/V3/A1/A2/M3/c1 ;
 wire \V2/V3/A1/A2/M3/c2 ;
 wire \V2/V3/A1/A2/M3/s1 ;
 wire \V2/V3/A1/A2/M4/c1 ;
 wire \V2/V3/A1/A2/M4/c2 ;
 wire \V2/V3/A1/A2/M4/s1 ;
 wire \V2/V3/A2/c1 ;
 wire \V2/V3/A2/A1/c1 ;
 wire \V2/V3/A2/A1/c2 ;
 wire \V2/V3/A2/A1/c3 ;
 wire \V2/V3/A2/A1/M1/c1 ;
 wire \V2/V3/A2/A1/M1/c2 ;
 wire \V2/V3/A2/A1/M1/s1 ;
 wire \V2/V3/A2/A1/M2/c1 ;
 wire \V2/V3/A2/A1/M2/c2 ;
 wire \V2/V3/A2/A1/M2/s1 ;
 wire \V2/V3/A2/A1/M3/c1 ;
 wire \V2/V3/A2/A1/M3/c2 ;
 wire \V2/V3/A2/A1/M3/s1 ;
 wire \V2/V3/A2/A1/M4/c1 ;
 wire \V2/V3/A2/A1/M4/c2 ;
 wire \V2/V3/A2/A1/M4/s1 ;
 wire \V2/V3/A2/A2/c1 ;
 wire \V2/V3/A2/A2/c2 ;
 wire \V2/V3/A2/A2/c3 ;
 wire \V2/V3/A2/A2/M1/c1 ;
 wire \V2/V3/A2/A2/M1/c2 ;
 wire \V2/V3/A2/A2/M1/s1 ;
 wire \V2/V3/A2/A2/M2/c1 ;
 wire \V2/V3/A2/A2/M2/c2 ;
 wire \V2/V3/A2/A2/M2/s1 ;
 wire \V2/V3/A2/A2/M3/c1 ;
 wire \V2/V3/A2/A2/M3/c2 ;
 wire \V2/V3/A2/A2/M3/s1 ;
 wire \V2/V3/A2/A2/M4/c1 ;
 wire \V2/V3/A2/A2/M4/c2 ;
 wire \V2/V3/A2/A2/M4/s1 ;
 wire \V2/V3/A3/c1 ;
 wire \V2/V3/A3/A1/c1 ;
 wire \V2/V3/A3/A1/c2 ;
 wire \V2/V3/A3/A1/c3 ;
 wire \V2/V3/A3/A1/M1/c1 ;
 wire \V2/V3/A3/A1/M1/c2 ;
 wire \V2/V3/A3/A1/M1/s1 ;
 wire \V2/V3/A3/A1/M2/c1 ;
 wire \V2/V3/A3/A1/M2/c2 ;
 wire \V2/V3/A3/A1/M2/s1 ;
 wire \V2/V3/A3/A1/M3/c1 ;
 wire \V2/V3/A3/A1/M3/c2 ;
 wire \V2/V3/A3/A1/M3/s1 ;
 wire \V2/V3/A3/A1/M4/c1 ;
 wire \V2/V3/A3/A1/M4/c2 ;
 wire \V2/V3/A3/A1/M4/s1 ;
 wire \V2/V3/A3/A2/c1 ;
 wire \V2/V3/A3/A2/c2 ;
 wire \V2/V3/A3/A2/c3 ;
 wire \V2/V3/A3/A2/M1/c1 ;
 wire \V2/V3/A3/A2/M1/c2 ;
 wire \V2/V3/A3/A2/M1/s1 ;
 wire \V2/V3/A3/A2/M2/c1 ;
 wire \V2/V3/A3/A2/M2/c2 ;
 wire \V2/V3/A3/A2/M2/s1 ;
 wire \V2/V3/A3/A2/M3/c1 ;
 wire \V2/V3/A3/A2/M3/c2 ;
 wire \V2/V3/A3/A2/M3/s1 ;
 wire \V2/V3/A3/A2/M4/c1 ;
 wire \V2/V3/A3/A2/M4/c2 ;
 wire \V2/V3/A3/A2/M4/s1 ;
 wire \V2/V3/V1/c1 ;
 wire \V2/V3/V1/c2 ;
 wire \V2/V3/V1/c3 ;
 wire \V2/V3/V1/overflow ;
 wire \V2/V3/V1/A1/c1 ;
 wire \V2/V3/V1/A1/c2 ;
 wire \V2/V3/V1/A1/c3 ;
 wire \V2/V3/V1/A1/M1/c1 ;
 wire \V2/V3/V1/A1/M1/c2 ;
 wire \V2/V3/V1/A1/M1/s1 ;
 wire \V2/V3/V1/A1/M2/c1 ;
 wire \V2/V3/V1/A1/M2/c2 ;
 wire \V2/V3/V1/A1/M2/s1 ;
 wire \V2/V3/V1/A1/M3/c1 ;
 wire \V2/V3/V1/A1/M3/c2 ;
 wire \V2/V3/V1/A1/M3/s1 ;
 wire \V2/V3/V1/A1/M4/c1 ;
 wire \V2/V3/V1/A1/M4/c2 ;
 wire \V2/V3/V1/A1/M4/s1 ;
 wire \V2/V3/V1/A2/c1 ;
 wire \V2/V3/V1/A2/c2 ;
 wire \V2/V3/V1/A2/c3 ;
 wire \V2/V3/V1/A2/M1/c1 ;
 wire \V2/V3/V1/A2/M1/c2 ;
 wire \V2/V3/V1/A2/M1/s1 ;
 wire \V2/V3/V1/A2/M2/c1 ;
 wire \V2/V3/V1/A2/M2/c2 ;
 wire \V2/V3/V1/A2/M2/s1 ;
 wire \V2/V3/V1/A2/M3/c1 ;
 wire \V2/V3/V1/A2/M3/c2 ;
 wire \V2/V3/V1/A2/M3/s1 ;
 wire \V2/V3/V1/A2/M4/c1 ;
 wire \V2/V3/V1/A2/M4/c2 ;
 wire \V2/V3/V1/A2/M4/s1 ;
 wire \V2/V3/V1/A3/c1 ;
 wire \V2/V3/V1/A3/c2 ;
 wire \V2/V3/V1/A3/c3 ;
 wire \V2/V3/V1/A3/M1/c1 ;
 wire \V2/V3/V1/A3/M1/c2 ;
 wire \V2/V3/V1/A3/M1/s1 ;
 wire \V2/V3/V1/A3/M2/c1 ;
 wire \V2/V3/V1/A3/M2/c2 ;
 wire \V2/V3/V1/A3/M2/s1 ;
 wire \V2/V3/V1/A3/M3/c1 ;
 wire \V2/V3/V1/A3/M3/c2 ;
 wire \V2/V3/V1/A3/M3/s1 ;
 wire \V2/V3/V1/A3/M4/c1 ;
 wire \V2/V3/V1/A3/M4/c2 ;
 wire \V2/V3/V1/A3/M4/s1 ;
 wire \V2/V3/V1/V1/w1 ;
 wire \V2/V3/V1/V1/w2 ;
 wire \V2/V3/V1/V1/w3 ;
 wire \V2/V3/V1/V1/w4 ;
 wire \V2/V3/V1/V2/w1 ;
 wire \V2/V3/V1/V2/w2 ;
 wire \V2/V3/V1/V2/w3 ;
 wire \V2/V3/V1/V2/w4 ;
 wire \V2/V3/V1/V3/w1 ;
 wire \V2/V3/V1/V3/w2 ;
 wire \V2/V3/V1/V3/w3 ;
 wire \V2/V3/V1/V3/w4 ;
 wire \V2/V3/V1/V4/w1 ;
 wire \V2/V3/V1/V4/w2 ;
 wire \V2/V3/V1/V4/w3 ;
 wire \V2/V3/V1/V4/w4 ;
 wire \V2/V3/V2/c1 ;
 wire \V2/V3/V2/c2 ;
 wire \V2/V3/V2/c3 ;
 wire \V2/V3/V2/overflow ;
 wire \V2/V3/V2/A1/c1 ;
 wire \V2/V3/V2/A1/c2 ;
 wire \V2/V3/V2/A1/c3 ;
 wire \V2/V3/V2/A1/M1/c1 ;
 wire \V2/V3/V2/A1/M1/c2 ;
 wire \V2/V3/V2/A1/M1/s1 ;
 wire \V2/V3/V2/A1/M2/c1 ;
 wire \V2/V3/V2/A1/M2/c2 ;
 wire \V2/V3/V2/A1/M2/s1 ;
 wire \V2/V3/V2/A1/M3/c1 ;
 wire \V2/V3/V2/A1/M3/c2 ;
 wire \V2/V3/V2/A1/M3/s1 ;
 wire \V2/V3/V2/A1/M4/c1 ;
 wire \V2/V3/V2/A1/M4/c2 ;
 wire \V2/V3/V2/A1/M4/s1 ;
 wire \V2/V3/V2/A2/c1 ;
 wire \V2/V3/V2/A2/c2 ;
 wire \V2/V3/V2/A2/c3 ;
 wire \V2/V3/V2/A2/M1/c1 ;
 wire \V2/V3/V2/A2/M1/c2 ;
 wire \V2/V3/V2/A2/M1/s1 ;
 wire \V2/V3/V2/A2/M2/c1 ;
 wire \V2/V3/V2/A2/M2/c2 ;
 wire \V2/V3/V2/A2/M2/s1 ;
 wire \V2/V3/V2/A2/M3/c1 ;
 wire \V2/V3/V2/A2/M3/c2 ;
 wire \V2/V3/V2/A2/M3/s1 ;
 wire \V2/V3/V2/A2/M4/c1 ;
 wire \V2/V3/V2/A2/M4/c2 ;
 wire \V2/V3/V2/A2/M4/s1 ;
 wire \V2/V3/V2/A3/c1 ;
 wire \V2/V3/V2/A3/c2 ;
 wire \V2/V3/V2/A3/c3 ;
 wire \V2/V3/V2/A3/M1/c1 ;
 wire \V2/V3/V2/A3/M1/c2 ;
 wire \V2/V3/V2/A3/M1/s1 ;
 wire \V2/V3/V2/A3/M2/c1 ;
 wire \V2/V3/V2/A3/M2/c2 ;
 wire \V2/V3/V2/A3/M2/s1 ;
 wire \V2/V3/V2/A3/M3/c1 ;
 wire \V2/V3/V2/A3/M3/c2 ;
 wire \V2/V3/V2/A3/M3/s1 ;
 wire \V2/V3/V2/A3/M4/c1 ;
 wire \V2/V3/V2/A3/M4/c2 ;
 wire \V2/V3/V2/A3/M4/s1 ;
 wire \V2/V3/V2/V1/w1 ;
 wire \V2/V3/V2/V1/w2 ;
 wire \V2/V3/V2/V1/w3 ;
 wire \V2/V3/V2/V1/w4 ;
 wire \V2/V3/V2/V2/w1 ;
 wire \V2/V3/V2/V2/w2 ;
 wire \V2/V3/V2/V2/w3 ;
 wire \V2/V3/V2/V2/w4 ;
 wire \V2/V3/V2/V3/w1 ;
 wire \V2/V3/V2/V3/w2 ;
 wire \V2/V3/V2/V3/w3 ;
 wire \V2/V3/V2/V3/w4 ;
 wire \V2/V3/V2/V4/w1 ;
 wire \V2/V3/V2/V4/w2 ;
 wire \V2/V3/V2/V4/w3 ;
 wire \V2/V3/V2/V4/w4 ;
 wire \V2/V3/V3/c1 ;
 wire \V2/V3/V3/c2 ;
 wire \V2/V3/V3/c3 ;
 wire \V2/V3/V3/overflow ;
 wire \V2/V3/V3/A1/c1 ;
 wire \V2/V3/V3/A1/c2 ;
 wire \V2/V3/V3/A1/c3 ;
 wire \V2/V3/V3/A1/M1/c1 ;
 wire \V2/V3/V3/A1/M1/c2 ;
 wire \V2/V3/V3/A1/M1/s1 ;
 wire \V2/V3/V3/A1/M2/c1 ;
 wire \V2/V3/V3/A1/M2/c2 ;
 wire \V2/V3/V3/A1/M2/s1 ;
 wire \V2/V3/V3/A1/M3/c1 ;
 wire \V2/V3/V3/A1/M3/c2 ;
 wire \V2/V3/V3/A1/M3/s1 ;
 wire \V2/V3/V3/A1/M4/c1 ;
 wire \V2/V3/V3/A1/M4/c2 ;
 wire \V2/V3/V3/A1/M4/s1 ;
 wire \V2/V3/V3/A2/c1 ;
 wire \V2/V3/V3/A2/c2 ;
 wire \V2/V3/V3/A2/c3 ;
 wire \V2/V3/V3/A2/M1/c1 ;
 wire \V2/V3/V3/A2/M1/c2 ;
 wire \V2/V3/V3/A2/M1/s1 ;
 wire \V2/V3/V3/A2/M2/c1 ;
 wire \V2/V3/V3/A2/M2/c2 ;
 wire \V2/V3/V3/A2/M2/s1 ;
 wire \V2/V3/V3/A2/M3/c1 ;
 wire \V2/V3/V3/A2/M3/c2 ;
 wire \V2/V3/V3/A2/M3/s1 ;
 wire \V2/V3/V3/A2/M4/c1 ;
 wire \V2/V3/V3/A2/M4/c2 ;
 wire \V2/V3/V3/A2/M4/s1 ;
 wire \V2/V3/V3/A3/c1 ;
 wire \V2/V3/V3/A3/c2 ;
 wire \V2/V3/V3/A3/c3 ;
 wire \V2/V3/V3/A3/M1/c1 ;
 wire \V2/V3/V3/A3/M1/c2 ;
 wire \V2/V3/V3/A3/M1/s1 ;
 wire \V2/V3/V3/A3/M2/c1 ;
 wire \V2/V3/V3/A3/M2/c2 ;
 wire \V2/V3/V3/A3/M2/s1 ;
 wire \V2/V3/V3/A3/M3/c1 ;
 wire \V2/V3/V3/A3/M3/c2 ;
 wire \V2/V3/V3/A3/M3/s1 ;
 wire \V2/V3/V3/A3/M4/c1 ;
 wire \V2/V3/V3/A3/M4/c2 ;
 wire \V2/V3/V3/A3/M4/s1 ;
 wire \V2/V3/V3/V1/w1 ;
 wire \V2/V3/V3/V1/w2 ;
 wire \V2/V3/V3/V1/w3 ;
 wire \V2/V3/V3/V1/w4 ;
 wire \V2/V3/V3/V2/w1 ;
 wire \V2/V3/V3/V2/w2 ;
 wire \V2/V3/V3/V2/w3 ;
 wire \V2/V3/V3/V2/w4 ;
 wire \V2/V3/V3/V3/w1 ;
 wire \V2/V3/V3/V3/w2 ;
 wire \V2/V3/V3/V3/w3 ;
 wire \V2/V3/V3/V3/w4 ;
 wire \V2/V3/V3/V4/w1 ;
 wire \V2/V3/V3/V4/w2 ;
 wire \V2/V3/V3/V4/w3 ;
 wire \V2/V3/V3/V4/w4 ;
 wire \V2/V3/V4/c1 ;
 wire \V2/V3/V4/c2 ;
 wire \V2/V3/V4/c3 ;
 wire \V2/V3/V4/overflow ;
 wire \V2/V3/V4/A1/c1 ;
 wire \V2/V3/V4/A1/c2 ;
 wire \V2/V3/V4/A1/c3 ;
 wire \V2/V3/V4/A1/M1/c1 ;
 wire \V2/V3/V4/A1/M1/c2 ;
 wire \V2/V3/V4/A1/M1/s1 ;
 wire \V2/V3/V4/A1/M2/c1 ;
 wire \V2/V3/V4/A1/M2/c2 ;
 wire \V2/V3/V4/A1/M2/s1 ;
 wire \V2/V3/V4/A1/M3/c1 ;
 wire \V2/V3/V4/A1/M3/c2 ;
 wire \V2/V3/V4/A1/M3/s1 ;
 wire \V2/V3/V4/A1/M4/c1 ;
 wire \V2/V3/V4/A1/M4/c2 ;
 wire \V2/V3/V4/A1/M4/s1 ;
 wire \V2/V3/V4/A2/c1 ;
 wire \V2/V3/V4/A2/c2 ;
 wire \V2/V3/V4/A2/c3 ;
 wire \V2/V3/V4/A2/M1/c1 ;
 wire \V2/V3/V4/A2/M1/c2 ;
 wire \V2/V3/V4/A2/M1/s1 ;
 wire \V2/V3/V4/A2/M2/c1 ;
 wire \V2/V3/V4/A2/M2/c2 ;
 wire \V2/V3/V4/A2/M2/s1 ;
 wire \V2/V3/V4/A2/M3/c1 ;
 wire \V2/V3/V4/A2/M3/c2 ;
 wire \V2/V3/V4/A2/M3/s1 ;
 wire \V2/V3/V4/A2/M4/c1 ;
 wire \V2/V3/V4/A2/M4/c2 ;
 wire \V2/V3/V4/A2/M4/s1 ;
 wire \V2/V3/V4/A3/c1 ;
 wire \V2/V3/V4/A3/c2 ;
 wire \V2/V3/V4/A3/c3 ;
 wire \V2/V3/V4/A3/M1/c1 ;
 wire \V2/V3/V4/A3/M1/c2 ;
 wire \V2/V3/V4/A3/M1/s1 ;
 wire \V2/V3/V4/A3/M2/c1 ;
 wire \V2/V3/V4/A3/M2/c2 ;
 wire \V2/V3/V4/A3/M2/s1 ;
 wire \V2/V3/V4/A3/M3/c1 ;
 wire \V2/V3/V4/A3/M3/c2 ;
 wire \V2/V3/V4/A3/M3/s1 ;
 wire \V2/V3/V4/A3/M4/c1 ;
 wire \V2/V3/V4/A3/M4/c2 ;
 wire \V2/V3/V4/A3/M4/s1 ;
 wire \V2/V3/V4/V1/w1 ;
 wire \V2/V3/V4/V1/w2 ;
 wire \V2/V3/V4/V1/w3 ;
 wire \V2/V3/V4/V1/w4 ;
 wire \V2/V3/V4/V2/w1 ;
 wire \V2/V3/V4/V2/w2 ;
 wire \V2/V3/V4/V2/w3 ;
 wire \V2/V3/V4/V2/w4 ;
 wire \V2/V3/V4/V3/w1 ;
 wire \V2/V3/V4/V3/w2 ;
 wire \V2/V3/V4/V3/w3 ;
 wire \V2/V3/V4/V3/w4 ;
 wire \V2/V3/V4/V4/w1 ;
 wire \V2/V3/V4/V4/w2 ;
 wire \V2/V3/V4/V4/w3 ;
 wire \V2/V3/V4/V4/w4 ;
 wire \V2/V4/c1 ;
 wire \V2/V4/c2 ;
 wire \V2/V4/c3 ;
 wire \V2/V4/overflow ;
 wire \V2/V4/A1/c1 ;
 wire \V2/V4/A1/A1/c1 ;
 wire \V2/V4/A1/A1/c2 ;
 wire \V2/V4/A1/A1/c3 ;
 wire \V2/V4/A1/A1/M1/c1 ;
 wire \V2/V4/A1/A1/M1/c2 ;
 wire \V2/V4/A1/A1/M1/s1 ;
 wire \V2/V4/A1/A1/M2/c1 ;
 wire \V2/V4/A1/A1/M2/c2 ;
 wire \V2/V4/A1/A1/M2/s1 ;
 wire \V2/V4/A1/A1/M3/c1 ;
 wire \V2/V4/A1/A1/M3/c2 ;
 wire \V2/V4/A1/A1/M3/s1 ;
 wire \V2/V4/A1/A1/M4/c1 ;
 wire \V2/V4/A1/A1/M4/c2 ;
 wire \V2/V4/A1/A1/M4/s1 ;
 wire \V2/V4/A1/A2/c1 ;
 wire \V2/V4/A1/A2/c2 ;
 wire \V2/V4/A1/A2/c3 ;
 wire \V2/V4/A1/A2/M1/c1 ;
 wire \V2/V4/A1/A2/M1/c2 ;
 wire \V2/V4/A1/A2/M1/s1 ;
 wire \V2/V4/A1/A2/M2/c1 ;
 wire \V2/V4/A1/A2/M2/c2 ;
 wire \V2/V4/A1/A2/M2/s1 ;
 wire \V2/V4/A1/A2/M3/c1 ;
 wire \V2/V4/A1/A2/M3/c2 ;
 wire \V2/V4/A1/A2/M3/s1 ;
 wire \V2/V4/A1/A2/M4/c1 ;
 wire \V2/V4/A1/A2/M4/c2 ;
 wire \V2/V4/A1/A2/M4/s1 ;
 wire \V2/V4/A2/c1 ;
 wire \V2/V4/A2/A1/c1 ;
 wire \V2/V4/A2/A1/c2 ;
 wire \V2/V4/A2/A1/c3 ;
 wire \V2/V4/A2/A1/M1/c1 ;
 wire \V2/V4/A2/A1/M1/c2 ;
 wire \V2/V4/A2/A1/M1/s1 ;
 wire \V2/V4/A2/A1/M2/c1 ;
 wire \V2/V4/A2/A1/M2/c2 ;
 wire \V2/V4/A2/A1/M2/s1 ;
 wire \V2/V4/A2/A1/M3/c1 ;
 wire \V2/V4/A2/A1/M3/c2 ;
 wire \V2/V4/A2/A1/M3/s1 ;
 wire \V2/V4/A2/A1/M4/c1 ;
 wire \V2/V4/A2/A1/M4/c2 ;
 wire \V2/V4/A2/A1/M4/s1 ;
 wire \V2/V4/A2/A2/c1 ;
 wire \V2/V4/A2/A2/c2 ;
 wire \V2/V4/A2/A2/c3 ;
 wire \V2/V4/A2/A2/M1/c1 ;
 wire \V2/V4/A2/A2/M1/c2 ;
 wire \V2/V4/A2/A2/M1/s1 ;
 wire \V2/V4/A2/A2/M2/c1 ;
 wire \V2/V4/A2/A2/M2/c2 ;
 wire \V2/V4/A2/A2/M2/s1 ;
 wire \V2/V4/A2/A2/M3/c1 ;
 wire \V2/V4/A2/A2/M3/c2 ;
 wire \V2/V4/A2/A2/M3/s1 ;
 wire \V2/V4/A2/A2/M4/c1 ;
 wire \V2/V4/A2/A2/M4/c2 ;
 wire \V2/V4/A2/A2/M4/s1 ;
 wire \V2/V4/A3/c1 ;
 wire \V2/V4/A3/A1/c1 ;
 wire \V2/V4/A3/A1/c2 ;
 wire \V2/V4/A3/A1/c3 ;
 wire \V2/V4/A3/A1/M1/c1 ;
 wire \V2/V4/A3/A1/M1/c2 ;
 wire \V2/V4/A3/A1/M1/s1 ;
 wire \V2/V4/A3/A1/M2/c1 ;
 wire \V2/V4/A3/A1/M2/c2 ;
 wire \V2/V4/A3/A1/M2/s1 ;
 wire \V2/V4/A3/A1/M3/c1 ;
 wire \V2/V4/A3/A1/M3/c2 ;
 wire \V2/V4/A3/A1/M3/s1 ;
 wire \V2/V4/A3/A1/M4/c1 ;
 wire \V2/V4/A3/A1/M4/c2 ;
 wire \V2/V4/A3/A1/M4/s1 ;
 wire \V2/V4/A3/A2/c1 ;
 wire \V2/V4/A3/A2/c2 ;
 wire \V2/V4/A3/A2/c3 ;
 wire \V2/V4/A3/A2/M1/c1 ;
 wire \V2/V4/A3/A2/M1/c2 ;
 wire \V2/V4/A3/A2/M1/s1 ;
 wire \V2/V4/A3/A2/M2/c1 ;
 wire \V2/V4/A3/A2/M2/c2 ;
 wire \V2/V4/A3/A2/M2/s1 ;
 wire \V2/V4/A3/A2/M3/c1 ;
 wire \V2/V4/A3/A2/M3/c2 ;
 wire \V2/V4/A3/A2/M3/s1 ;
 wire \V2/V4/A3/A2/M4/c1 ;
 wire \V2/V4/A3/A2/M4/c2 ;
 wire \V2/V4/A3/A2/M4/s1 ;
 wire \V2/V4/V1/c1 ;
 wire \V2/V4/V1/c2 ;
 wire \V2/V4/V1/c3 ;
 wire \V2/V4/V1/overflow ;
 wire \V2/V4/V1/A1/c1 ;
 wire \V2/V4/V1/A1/c2 ;
 wire \V2/V4/V1/A1/c3 ;
 wire \V2/V4/V1/A1/M1/c1 ;
 wire \V2/V4/V1/A1/M1/c2 ;
 wire \V2/V4/V1/A1/M1/s1 ;
 wire \V2/V4/V1/A1/M2/c1 ;
 wire \V2/V4/V1/A1/M2/c2 ;
 wire \V2/V4/V1/A1/M2/s1 ;
 wire \V2/V4/V1/A1/M3/c1 ;
 wire \V2/V4/V1/A1/M3/c2 ;
 wire \V2/V4/V1/A1/M3/s1 ;
 wire \V2/V4/V1/A1/M4/c1 ;
 wire \V2/V4/V1/A1/M4/c2 ;
 wire \V2/V4/V1/A1/M4/s1 ;
 wire \V2/V4/V1/A2/c1 ;
 wire \V2/V4/V1/A2/c2 ;
 wire \V2/V4/V1/A2/c3 ;
 wire \V2/V4/V1/A2/M1/c1 ;
 wire \V2/V4/V1/A2/M1/c2 ;
 wire \V2/V4/V1/A2/M1/s1 ;
 wire \V2/V4/V1/A2/M2/c1 ;
 wire \V2/V4/V1/A2/M2/c2 ;
 wire \V2/V4/V1/A2/M2/s1 ;
 wire \V2/V4/V1/A2/M3/c1 ;
 wire \V2/V4/V1/A2/M3/c2 ;
 wire \V2/V4/V1/A2/M3/s1 ;
 wire \V2/V4/V1/A2/M4/c1 ;
 wire \V2/V4/V1/A2/M4/c2 ;
 wire \V2/V4/V1/A2/M4/s1 ;
 wire \V2/V4/V1/A3/c1 ;
 wire \V2/V4/V1/A3/c2 ;
 wire \V2/V4/V1/A3/c3 ;
 wire \V2/V4/V1/A3/M1/c1 ;
 wire \V2/V4/V1/A3/M1/c2 ;
 wire \V2/V4/V1/A3/M1/s1 ;
 wire \V2/V4/V1/A3/M2/c1 ;
 wire \V2/V4/V1/A3/M2/c2 ;
 wire \V2/V4/V1/A3/M2/s1 ;
 wire \V2/V4/V1/A3/M3/c1 ;
 wire \V2/V4/V1/A3/M3/c2 ;
 wire \V2/V4/V1/A3/M3/s1 ;
 wire \V2/V4/V1/A3/M4/c1 ;
 wire \V2/V4/V1/A3/M4/c2 ;
 wire \V2/V4/V1/A3/M4/s1 ;
 wire \V2/V4/V1/V1/w1 ;
 wire \V2/V4/V1/V1/w2 ;
 wire \V2/V4/V1/V1/w3 ;
 wire \V2/V4/V1/V1/w4 ;
 wire \V2/V4/V1/V2/w1 ;
 wire \V2/V4/V1/V2/w2 ;
 wire \V2/V4/V1/V2/w3 ;
 wire \V2/V4/V1/V2/w4 ;
 wire \V2/V4/V1/V3/w1 ;
 wire \V2/V4/V1/V3/w2 ;
 wire \V2/V4/V1/V3/w3 ;
 wire \V2/V4/V1/V3/w4 ;
 wire \V2/V4/V1/V4/w1 ;
 wire \V2/V4/V1/V4/w2 ;
 wire \V2/V4/V1/V4/w3 ;
 wire \V2/V4/V1/V4/w4 ;
 wire \V2/V4/V2/c1 ;
 wire \V2/V4/V2/c2 ;
 wire \V2/V4/V2/c3 ;
 wire \V2/V4/V2/overflow ;
 wire \V2/V4/V2/A1/c1 ;
 wire \V2/V4/V2/A1/c2 ;
 wire \V2/V4/V2/A1/c3 ;
 wire \V2/V4/V2/A1/M1/c1 ;
 wire \V2/V4/V2/A1/M1/c2 ;
 wire \V2/V4/V2/A1/M1/s1 ;
 wire \V2/V4/V2/A1/M2/c1 ;
 wire \V2/V4/V2/A1/M2/c2 ;
 wire \V2/V4/V2/A1/M2/s1 ;
 wire \V2/V4/V2/A1/M3/c1 ;
 wire \V2/V4/V2/A1/M3/c2 ;
 wire \V2/V4/V2/A1/M3/s1 ;
 wire \V2/V4/V2/A1/M4/c1 ;
 wire \V2/V4/V2/A1/M4/c2 ;
 wire \V2/V4/V2/A1/M4/s1 ;
 wire \V2/V4/V2/A2/c1 ;
 wire \V2/V4/V2/A2/c2 ;
 wire \V2/V4/V2/A2/c3 ;
 wire \V2/V4/V2/A2/M1/c1 ;
 wire \V2/V4/V2/A2/M1/c2 ;
 wire \V2/V4/V2/A2/M1/s1 ;
 wire \V2/V4/V2/A2/M2/c1 ;
 wire \V2/V4/V2/A2/M2/c2 ;
 wire \V2/V4/V2/A2/M2/s1 ;
 wire \V2/V4/V2/A2/M3/c1 ;
 wire \V2/V4/V2/A2/M3/c2 ;
 wire \V2/V4/V2/A2/M3/s1 ;
 wire \V2/V4/V2/A2/M4/c1 ;
 wire \V2/V4/V2/A2/M4/c2 ;
 wire \V2/V4/V2/A2/M4/s1 ;
 wire \V2/V4/V2/A3/c1 ;
 wire \V2/V4/V2/A3/c2 ;
 wire \V2/V4/V2/A3/c3 ;
 wire \V2/V4/V2/A3/M1/c1 ;
 wire \V2/V4/V2/A3/M1/c2 ;
 wire \V2/V4/V2/A3/M1/s1 ;
 wire \V2/V4/V2/A3/M2/c1 ;
 wire \V2/V4/V2/A3/M2/c2 ;
 wire \V2/V4/V2/A3/M2/s1 ;
 wire \V2/V4/V2/A3/M3/c1 ;
 wire \V2/V4/V2/A3/M3/c2 ;
 wire \V2/V4/V2/A3/M3/s1 ;
 wire \V2/V4/V2/A3/M4/c1 ;
 wire \V2/V4/V2/A3/M4/c2 ;
 wire \V2/V4/V2/A3/M4/s1 ;
 wire \V2/V4/V2/V1/w1 ;
 wire \V2/V4/V2/V1/w2 ;
 wire \V2/V4/V2/V1/w3 ;
 wire \V2/V4/V2/V1/w4 ;
 wire \V2/V4/V2/V2/w1 ;
 wire \V2/V4/V2/V2/w2 ;
 wire \V2/V4/V2/V2/w3 ;
 wire \V2/V4/V2/V2/w4 ;
 wire \V2/V4/V2/V3/w1 ;
 wire \V2/V4/V2/V3/w2 ;
 wire \V2/V4/V2/V3/w3 ;
 wire \V2/V4/V2/V3/w4 ;
 wire \V2/V4/V2/V4/w1 ;
 wire \V2/V4/V2/V4/w2 ;
 wire \V2/V4/V2/V4/w3 ;
 wire \V2/V4/V2/V4/w4 ;
 wire \V2/V4/V3/c1 ;
 wire \V2/V4/V3/c2 ;
 wire \V2/V4/V3/c3 ;
 wire \V2/V4/V3/overflow ;
 wire \V2/V4/V3/A1/c1 ;
 wire \V2/V4/V3/A1/c2 ;
 wire \V2/V4/V3/A1/c3 ;
 wire \V2/V4/V3/A1/M1/c1 ;
 wire \V2/V4/V3/A1/M1/c2 ;
 wire \V2/V4/V3/A1/M1/s1 ;
 wire \V2/V4/V3/A1/M2/c1 ;
 wire \V2/V4/V3/A1/M2/c2 ;
 wire \V2/V4/V3/A1/M2/s1 ;
 wire \V2/V4/V3/A1/M3/c1 ;
 wire \V2/V4/V3/A1/M3/c2 ;
 wire \V2/V4/V3/A1/M3/s1 ;
 wire \V2/V4/V3/A1/M4/c1 ;
 wire \V2/V4/V3/A1/M4/c2 ;
 wire \V2/V4/V3/A1/M4/s1 ;
 wire \V2/V4/V3/A2/c1 ;
 wire \V2/V4/V3/A2/c2 ;
 wire \V2/V4/V3/A2/c3 ;
 wire \V2/V4/V3/A2/M1/c1 ;
 wire \V2/V4/V3/A2/M1/c2 ;
 wire \V2/V4/V3/A2/M1/s1 ;
 wire \V2/V4/V3/A2/M2/c1 ;
 wire \V2/V4/V3/A2/M2/c2 ;
 wire \V2/V4/V3/A2/M2/s1 ;
 wire \V2/V4/V3/A2/M3/c1 ;
 wire \V2/V4/V3/A2/M3/c2 ;
 wire \V2/V4/V3/A2/M3/s1 ;
 wire \V2/V4/V3/A2/M4/c1 ;
 wire \V2/V4/V3/A2/M4/c2 ;
 wire \V2/V4/V3/A2/M4/s1 ;
 wire \V2/V4/V3/A3/c1 ;
 wire \V2/V4/V3/A3/c2 ;
 wire \V2/V4/V3/A3/c3 ;
 wire \V2/V4/V3/A3/M1/c1 ;
 wire \V2/V4/V3/A3/M1/c2 ;
 wire \V2/V4/V3/A3/M1/s1 ;
 wire \V2/V4/V3/A3/M2/c1 ;
 wire \V2/V4/V3/A3/M2/c2 ;
 wire \V2/V4/V3/A3/M2/s1 ;
 wire \V2/V4/V3/A3/M3/c1 ;
 wire \V2/V4/V3/A3/M3/c2 ;
 wire \V2/V4/V3/A3/M3/s1 ;
 wire \V2/V4/V3/A3/M4/c1 ;
 wire \V2/V4/V3/A3/M4/c2 ;
 wire \V2/V4/V3/A3/M4/s1 ;
 wire \V2/V4/V3/V1/w1 ;
 wire \V2/V4/V3/V1/w2 ;
 wire \V2/V4/V3/V1/w3 ;
 wire \V2/V4/V3/V1/w4 ;
 wire \V2/V4/V3/V2/w1 ;
 wire \V2/V4/V3/V2/w2 ;
 wire \V2/V4/V3/V2/w3 ;
 wire \V2/V4/V3/V2/w4 ;
 wire \V2/V4/V3/V3/w1 ;
 wire \V2/V4/V3/V3/w2 ;
 wire \V2/V4/V3/V3/w3 ;
 wire \V2/V4/V3/V3/w4 ;
 wire \V2/V4/V3/V4/w1 ;
 wire \V2/V4/V3/V4/w2 ;
 wire \V2/V4/V3/V4/w3 ;
 wire \V2/V4/V3/V4/w4 ;
 wire \V2/V4/V4/c1 ;
 wire \V2/V4/V4/c2 ;
 wire \V2/V4/V4/c3 ;
 wire \V2/V4/V4/overflow ;
 wire \V2/V4/V4/A1/c1 ;
 wire \V2/V4/V4/A1/c2 ;
 wire \V2/V4/V4/A1/c3 ;
 wire \V2/V4/V4/A1/M1/c1 ;
 wire \V2/V4/V4/A1/M1/c2 ;
 wire \V2/V4/V4/A1/M1/s1 ;
 wire \V2/V4/V4/A1/M2/c1 ;
 wire \V2/V4/V4/A1/M2/c2 ;
 wire \V2/V4/V4/A1/M2/s1 ;
 wire \V2/V4/V4/A1/M3/c1 ;
 wire \V2/V4/V4/A1/M3/c2 ;
 wire \V2/V4/V4/A1/M3/s1 ;
 wire \V2/V4/V4/A1/M4/c1 ;
 wire \V2/V4/V4/A1/M4/c2 ;
 wire \V2/V4/V4/A1/M4/s1 ;
 wire \V2/V4/V4/A2/c1 ;
 wire \V2/V4/V4/A2/c2 ;
 wire \V2/V4/V4/A2/c3 ;
 wire \V2/V4/V4/A2/M1/c1 ;
 wire \V2/V4/V4/A2/M1/c2 ;
 wire \V2/V4/V4/A2/M1/s1 ;
 wire \V2/V4/V4/A2/M2/c1 ;
 wire \V2/V4/V4/A2/M2/c2 ;
 wire \V2/V4/V4/A2/M2/s1 ;
 wire \V2/V4/V4/A2/M3/c1 ;
 wire \V2/V4/V4/A2/M3/c2 ;
 wire \V2/V4/V4/A2/M3/s1 ;
 wire \V2/V4/V4/A2/M4/c1 ;
 wire \V2/V4/V4/A2/M4/c2 ;
 wire \V2/V4/V4/A2/M4/s1 ;
 wire \V2/V4/V4/A3/c1 ;
 wire \V2/V4/V4/A3/c2 ;
 wire \V2/V4/V4/A3/c3 ;
 wire \V2/V4/V4/A3/M1/c1 ;
 wire \V2/V4/V4/A3/M1/c2 ;
 wire \V2/V4/V4/A3/M1/s1 ;
 wire \V2/V4/V4/A3/M2/c1 ;
 wire \V2/V4/V4/A3/M2/c2 ;
 wire \V2/V4/V4/A3/M2/s1 ;
 wire \V2/V4/V4/A3/M3/c1 ;
 wire \V2/V4/V4/A3/M3/c2 ;
 wire \V2/V4/V4/A3/M3/s1 ;
 wire \V2/V4/V4/A3/M4/c1 ;
 wire \V2/V4/V4/A3/M4/c2 ;
 wire \V2/V4/V4/A3/M4/s1 ;
 wire \V2/V4/V4/V1/w1 ;
 wire \V2/V4/V4/V1/w2 ;
 wire \V2/V4/V4/V1/w3 ;
 wire \V2/V4/V4/V1/w4 ;
 wire \V2/V4/V4/V2/w1 ;
 wire \V2/V4/V4/V2/w2 ;
 wire \V2/V4/V4/V2/w3 ;
 wire \V2/V4/V4/V2/w4 ;
 wire \V2/V4/V4/V3/w1 ;
 wire \V2/V4/V4/V3/w2 ;
 wire \V2/V4/V4/V3/w3 ;
 wire \V2/V4/V4/V3/w4 ;
 wire \V2/V4/V4/V4/w1 ;
 wire \V2/V4/V4/V4/w2 ;
 wire \V2/V4/V4/V4/w3 ;
 wire \V2/V4/V4/V4/w4 ;
 wire \V3/c1 ;
 wire \V3/c2 ;
 wire \V3/c3 ;
 wire \V3/overflow ;
 wire \V3/A1/c1 ;
 wire \V3/A1/A1/c1 ;
 wire \V3/A1/A1/A1/c1 ;
 wire \V3/A1/A1/A1/c2 ;
 wire \V3/A1/A1/A1/c3 ;
 wire \V3/A1/A1/A1/M1/c1 ;
 wire \V3/A1/A1/A1/M1/c2 ;
 wire \V3/A1/A1/A1/M1/s1 ;
 wire \V3/A1/A1/A1/M2/c1 ;
 wire \V3/A1/A1/A1/M2/c2 ;
 wire \V3/A1/A1/A1/M2/s1 ;
 wire \V3/A1/A1/A1/M3/c1 ;
 wire \V3/A1/A1/A1/M3/c2 ;
 wire \V3/A1/A1/A1/M3/s1 ;
 wire \V3/A1/A1/A1/M4/c1 ;
 wire \V3/A1/A1/A1/M4/c2 ;
 wire \V3/A1/A1/A1/M4/s1 ;
 wire \V3/A1/A1/A2/c1 ;
 wire \V3/A1/A1/A2/c2 ;
 wire \V3/A1/A1/A2/c3 ;
 wire \V3/A1/A1/A2/M1/c1 ;
 wire \V3/A1/A1/A2/M1/c2 ;
 wire \V3/A1/A1/A2/M1/s1 ;
 wire \V3/A1/A1/A2/M2/c1 ;
 wire \V3/A1/A1/A2/M2/c2 ;
 wire \V3/A1/A1/A2/M2/s1 ;
 wire \V3/A1/A1/A2/M3/c1 ;
 wire \V3/A1/A1/A2/M3/c2 ;
 wire \V3/A1/A1/A2/M3/s1 ;
 wire \V3/A1/A1/A2/M4/c1 ;
 wire \V3/A1/A1/A2/M4/c2 ;
 wire \V3/A1/A1/A2/M4/s1 ;
 wire \V3/A1/A2/c1 ;
 wire \V3/A1/A2/A1/c1 ;
 wire \V3/A1/A2/A1/c2 ;
 wire \V3/A1/A2/A1/c3 ;
 wire \V3/A1/A2/A1/M1/c1 ;
 wire \V3/A1/A2/A1/M1/c2 ;
 wire \V3/A1/A2/A1/M1/s1 ;
 wire \V3/A1/A2/A1/M2/c1 ;
 wire \V3/A1/A2/A1/M2/c2 ;
 wire \V3/A1/A2/A1/M2/s1 ;
 wire \V3/A1/A2/A1/M3/c1 ;
 wire \V3/A1/A2/A1/M3/c2 ;
 wire \V3/A1/A2/A1/M3/s1 ;
 wire \V3/A1/A2/A1/M4/c1 ;
 wire \V3/A1/A2/A1/M4/c2 ;
 wire \V3/A1/A2/A1/M4/s1 ;
 wire \V3/A1/A2/A2/c1 ;
 wire \V3/A1/A2/A2/c2 ;
 wire \V3/A1/A2/A2/c3 ;
 wire \V3/A1/A2/A2/M1/c1 ;
 wire \V3/A1/A2/A2/M1/c2 ;
 wire \V3/A1/A2/A2/M1/s1 ;
 wire \V3/A1/A2/A2/M2/c1 ;
 wire \V3/A1/A2/A2/M2/c2 ;
 wire \V3/A1/A2/A2/M2/s1 ;
 wire \V3/A1/A2/A2/M3/c1 ;
 wire \V3/A1/A2/A2/M3/c2 ;
 wire \V3/A1/A2/A2/M3/s1 ;
 wire \V3/A1/A2/A2/M4/c1 ;
 wire \V3/A1/A2/A2/M4/c2 ;
 wire \V3/A1/A2/A2/M4/s1 ;
 wire \V3/A2/c1 ;
 wire \V3/A2/A1/c1 ;
 wire \V3/A2/A1/A1/c1 ;
 wire \V3/A2/A1/A1/c2 ;
 wire \V3/A2/A1/A1/c3 ;
 wire \V3/A2/A1/A1/M1/c1 ;
 wire \V3/A2/A1/A1/M1/c2 ;
 wire \V3/A2/A1/A1/M1/s1 ;
 wire \V3/A2/A1/A1/M2/c1 ;
 wire \V3/A2/A1/A1/M2/c2 ;
 wire \V3/A2/A1/A1/M2/s1 ;
 wire \V3/A2/A1/A1/M3/c1 ;
 wire \V3/A2/A1/A1/M3/c2 ;
 wire \V3/A2/A1/A1/M3/s1 ;
 wire \V3/A2/A1/A1/M4/c1 ;
 wire \V3/A2/A1/A1/M4/c2 ;
 wire \V3/A2/A1/A1/M4/s1 ;
 wire \V3/A2/A1/A2/c1 ;
 wire \V3/A2/A1/A2/c2 ;
 wire \V3/A2/A1/A2/c3 ;
 wire \V3/A2/A1/A2/M1/c1 ;
 wire \V3/A2/A1/A2/M1/c2 ;
 wire \V3/A2/A1/A2/M1/s1 ;
 wire \V3/A2/A1/A2/M2/c1 ;
 wire \V3/A2/A1/A2/M2/c2 ;
 wire \V3/A2/A1/A2/M2/s1 ;
 wire \V3/A2/A1/A2/M3/c1 ;
 wire \V3/A2/A1/A2/M3/c2 ;
 wire \V3/A2/A1/A2/M3/s1 ;
 wire \V3/A2/A1/A2/M4/c1 ;
 wire \V3/A2/A1/A2/M4/c2 ;
 wire \V3/A2/A1/A2/M4/s1 ;
 wire \V3/A2/A2/c1 ;
 wire \V3/A2/A2/A1/c1 ;
 wire \V3/A2/A2/A1/c2 ;
 wire \V3/A2/A2/A1/c3 ;
 wire \V3/A2/A2/A1/M1/c1 ;
 wire \V3/A2/A2/A1/M1/c2 ;
 wire \V3/A2/A2/A1/M1/s1 ;
 wire \V3/A2/A2/A1/M2/c1 ;
 wire \V3/A2/A2/A1/M2/c2 ;
 wire \V3/A2/A2/A1/M2/s1 ;
 wire \V3/A2/A2/A1/M3/c1 ;
 wire \V3/A2/A2/A1/M3/c2 ;
 wire \V3/A2/A2/A1/M3/s1 ;
 wire \V3/A2/A2/A1/M4/c1 ;
 wire \V3/A2/A2/A1/M4/c2 ;
 wire \V3/A2/A2/A1/M4/s1 ;
 wire \V3/A2/A2/A2/c1 ;
 wire \V3/A2/A2/A2/c2 ;
 wire \V3/A2/A2/A2/c3 ;
 wire \V3/A2/A2/A2/M1/c1 ;
 wire \V3/A2/A2/A2/M1/c2 ;
 wire \V3/A2/A2/A2/M1/s1 ;
 wire \V3/A2/A2/A2/M2/c1 ;
 wire \V3/A2/A2/A2/M2/c2 ;
 wire \V3/A2/A2/A2/M2/s1 ;
 wire \V3/A2/A2/A2/M3/c1 ;
 wire \V3/A2/A2/A2/M3/c2 ;
 wire \V3/A2/A2/A2/M3/s1 ;
 wire \V3/A2/A2/A2/M4/c1 ;
 wire \V3/A2/A2/A2/M4/c2 ;
 wire \V3/A2/A2/A2/M4/s1 ;
 wire \V3/A3/c1 ;
 wire \V3/A3/A1/c1 ;
 wire \V3/A3/A1/A1/c1 ;
 wire \V3/A3/A1/A1/c2 ;
 wire \V3/A3/A1/A1/c3 ;
 wire \V3/A3/A1/A1/M1/c1 ;
 wire \V3/A3/A1/A1/M1/c2 ;
 wire \V3/A3/A1/A1/M1/s1 ;
 wire \V3/A3/A1/A1/M2/c1 ;
 wire \V3/A3/A1/A1/M2/c2 ;
 wire \V3/A3/A1/A1/M2/s1 ;
 wire \V3/A3/A1/A1/M3/c1 ;
 wire \V3/A3/A1/A1/M3/c2 ;
 wire \V3/A3/A1/A1/M3/s1 ;
 wire \V3/A3/A1/A1/M4/c1 ;
 wire \V3/A3/A1/A1/M4/c2 ;
 wire \V3/A3/A1/A1/M4/s1 ;
 wire \V3/A3/A1/A2/c1 ;
 wire \V3/A3/A1/A2/c2 ;
 wire \V3/A3/A1/A2/c3 ;
 wire \V3/A3/A1/A2/M1/c1 ;
 wire \V3/A3/A1/A2/M1/c2 ;
 wire \V3/A3/A1/A2/M1/s1 ;
 wire \V3/A3/A1/A2/M2/c1 ;
 wire \V3/A3/A1/A2/M2/c2 ;
 wire \V3/A3/A1/A2/M2/s1 ;
 wire \V3/A3/A1/A2/M3/c1 ;
 wire \V3/A3/A1/A2/M3/c2 ;
 wire \V3/A3/A1/A2/M3/s1 ;
 wire \V3/A3/A1/A2/M4/c1 ;
 wire \V3/A3/A1/A2/M4/c2 ;
 wire \V3/A3/A1/A2/M4/s1 ;
 wire \V3/A3/A2/c1 ;
 wire \V3/A3/A2/A1/c1 ;
 wire \V3/A3/A2/A1/c2 ;
 wire \V3/A3/A2/A1/c3 ;
 wire \V3/A3/A2/A1/M1/c1 ;
 wire \V3/A3/A2/A1/M1/c2 ;
 wire \V3/A3/A2/A1/M1/s1 ;
 wire \V3/A3/A2/A1/M2/c1 ;
 wire \V3/A3/A2/A1/M2/c2 ;
 wire \V3/A3/A2/A1/M2/s1 ;
 wire \V3/A3/A2/A1/M3/c1 ;
 wire \V3/A3/A2/A1/M3/c2 ;
 wire \V3/A3/A2/A1/M3/s1 ;
 wire \V3/A3/A2/A1/M4/c1 ;
 wire \V3/A3/A2/A1/M4/c2 ;
 wire \V3/A3/A2/A1/M4/s1 ;
 wire \V3/A3/A2/A2/c1 ;
 wire \V3/A3/A2/A2/c2 ;
 wire \V3/A3/A2/A2/c3 ;
 wire \V3/A3/A2/A2/M1/c1 ;
 wire \V3/A3/A2/A2/M1/c2 ;
 wire \V3/A3/A2/A2/M1/s1 ;
 wire \V3/A3/A2/A2/M2/c1 ;
 wire \V3/A3/A2/A2/M2/c2 ;
 wire \V3/A3/A2/A2/M2/s1 ;
 wire \V3/A3/A2/A2/M3/c1 ;
 wire \V3/A3/A2/A2/M3/c2 ;
 wire \V3/A3/A2/A2/M3/s1 ;
 wire \V3/A3/A2/A2/M4/c1 ;
 wire \V3/A3/A2/A2/M4/c2 ;
 wire \V3/A3/A2/A2/M4/s1 ;
 wire \V3/V1/c1 ;
 wire \V3/V1/c2 ;
 wire \V3/V1/c3 ;
 wire \V3/V1/overflow ;
 wire \V3/V1/A1/c1 ;
 wire \V3/V1/A1/A1/c1 ;
 wire \V3/V1/A1/A1/c2 ;
 wire \V3/V1/A1/A1/c3 ;
 wire \V3/V1/A1/A1/M1/c1 ;
 wire \V3/V1/A1/A1/M1/c2 ;
 wire \V3/V1/A1/A1/M1/s1 ;
 wire \V3/V1/A1/A1/M2/c1 ;
 wire \V3/V1/A1/A1/M2/c2 ;
 wire \V3/V1/A1/A1/M2/s1 ;
 wire \V3/V1/A1/A1/M3/c1 ;
 wire \V3/V1/A1/A1/M3/c2 ;
 wire \V3/V1/A1/A1/M3/s1 ;
 wire \V3/V1/A1/A1/M4/c1 ;
 wire \V3/V1/A1/A1/M4/c2 ;
 wire \V3/V1/A1/A1/M4/s1 ;
 wire \V3/V1/A1/A2/c1 ;
 wire \V3/V1/A1/A2/c2 ;
 wire \V3/V1/A1/A2/c3 ;
 wire \V3/V1/A1/A2/M1/c1 ;
 wire \V3/V1/A1/A2/M1/c2 ;
 wire \V3/V1/A1/A2/M1/s1 ;
 wire \V3/V1/A1/A2/M2/c1 ;
 wire \V3/V1/A1/A2/M2/c2 ;
 wire \V3/V1/A1/A2/M2/s1 ;
 wire \V3/V1/A1/A2/M3/c1 ;
 wire \V3/V1/A1/A2/M3/c2 ;
 wire \V3/V1/A1/A2/M3/s1 ;
 wire \V3/V1/A1/A2/M4/c1 ;
 wire \V3/V1/A1/A2/M4/c2 ;
 wire \V3/V1/A1/A2/M4/s1 ;
 wire \V3/V1/A2/c1 ;
 wire \V3/V1/A2/A1/c1 ;
 wire \V3/V1/A2/A1/c2 ;
 wire \V3/V1/A2/A1/c3 ;
 wire \V3/V1/A2/A1/M1/c1 ;
 wire \V3/V1/A2/A1/M1/c2 ;
 wire \V3/V1/A2/A1/M1/s1 ;
 wire \V3/V1/A2/A1/M2/c1 ;
 wire \V3/V1/A2/A1/M2/c2 ;
 wire \V3/V1/A2/A1/M2/s1 ;
 wire \V3/V1/A2/A1/M3/c1 ;
 wire \V3/V1/A2/A1/M3/c2 ;
 wire \V3/V1/A2/A1/M3/s1 ;
 wire \V3/V1/A2/A1/M4/c1 ;
 wire \V3/V1/A2/A1/M4/c2 ;
 wire \V3/V1/A2/A1/M4/s1 ;
 wire \V3/V1/A2/A2/c1 ;
 wire \V3/V1/A2/A2/c2 ;
 wire \V3/V1/A2/A2/c3 ;
 wire \V3/V1/A2/A2/M1/c1 ;
 wire \V3/V1/A2/A2/M1/c2 ;
 wire \V3/V1/A2/A2/M1/s1 ;
 wire \V3/V1/A2/A2/M2/c1 ;
 wire \V3/V1/A2/A2/M2/c2 ;
 wire \V3/V1/A2/A2/M2/s1 ;
 wire \V3/V1/A2/A2/M3/c1 ;
 wire \V3/V1/A2/A2/M3/c2 ;
 wire \V3/V1/A2/A2/M3/s1 ;
 wire \V3/V1/A2/A2/M4/c1 ;
 wire \V3/V1/A2/A2/M4/c2 ;
 wire \V3/V1/A2/A2/M4/s1 ;
 wire \V3/V1/A3/c1 ;
 wire \V3/V1/A3/A1/c1 ;
 wire \V3/V1/A3/A1/c2 ;
 wire \V3/V1/A3/A1/c3 ;
 wire \V3/V1/A3/A1/M1/c1 ;
 wire \V3/V1/A3/A1/M1/c2 ;
 wire \V3/V1/A3/A1/M1/s1 ;
 wire \V3/V1/A3/A1/M2/c1 ;
 wire \V3/V1/A3/A1/M2/c2 ;
 wire \V3/V1/A3/A1/M2/s1 ;
 wire \V3/V1/A3/A1/M3/c1 ;
 wire \V3/V1/A3/A1/M3/c2 ;
 wire \V3/V1/A3/A1/M3/s1 ;
 wire \V3/V1/A3/A1/M4/c1 ;
 wire \V3/V1/A3/A1/M4/c2 ;
 wire \V3/V1/A3/A1/M4/s1 ;
 wire \V3/V1/A3/A2/c1 ;
 wire \V3/V1/A3/A2/c2 ;
 wire \V3/V1/A3/A2/c3 ;
 wire \V3/V1/A3/A2/M1/c1 ;
 wire \V3/V1/A3/A2/M1/c2 ;
 wire \V3/V1/A3/A2/M1/s1 ;
 wire \V3/V1/A3/A2/M2/c1 ;
 wire \V3/V1/A3/A2/M2/c2 ;
 wire \V3/V1/A3/A2/M2/s1 ;
 wire \V3/V1/A3/A2/M3/c1 ;
 wire \V3/V1/A3/A2/M3/c2 ;
 wire \V3/V1/A3/A2/M3/s1 ;
 wire \V3/V1/A3/A2/M4/c1 ;
 wire \V3/V1/A3/A2/M4/c2 ;
 wire \V3/V1/A3/A2/M4/s1 ;
 wire \V3/V1/V1/c1 ;
 wire \V3/V1/V1/c2 ;
 wire \V3/V1/V1/c3 ;
 wire \V3/V1/V1/overflow ;
 wire \V3/V1/V1/A1/c1 ;
 wire \V3/V1/V1/A1/c2 ;
 wire \V3/V1/V1/A1/c3 ;
 wire \V3/V1/V1/A1/M1/c1 ;
 wire \V3/V1/V1/A1/M1/c2 ;
 wire \V3/V1/V1/A1/M1/s1 ;
 wire \V3/V1/V1/A1/M2/c1 ;
 wire \V3/V1/V1/A1/M2/c2 ;
 wire \V3/V1/V1/A1/M2/s1 ;
 wire \V3/V1/V1/A1/M3/c1 ;
 wire \V3/V1/V1/A1/M3/c2 ;
 wire \V3/V1/V1/A1/M3/s1 ;
 wire \V3/V1/V1/A1/M4/c1 ;
 wire \V3/V1/V1/A1/M4/c2 ;
 wire \V3/V1/V1/A1/M4/s1 ;
 wire \V3/V1/V1/A2/c1 ;
 wire \V3/V1/V1/A2/c2 ;
 wire \V3/V1/V1/A2/c3 ;
 wire \V3/V1/V1/A2/M1/c1 ;
 wire \V3/V1/V1/A2/M1/c2 ;
 wire \V3/V1/V1/A2/M1/s1 ;
 wire \V3/V1/V1/A2/M2/c1 ;
 wire \V3/V1/V1/A2/M2/c2 ;
 wire \V3/V1/V1/A2/M2/s1 ;
 wire \V3/V1/V1/A2/M3/c1 ;
 wire \V3/V1/V1/A2/M3/c2 ;
 wire \V3/V1/V1/A2/M3/s1 ;
 wire \V3/V1/V1/A2/M4/c1 ;
 wire \V3/V1/V1/A2/M4/c2 ;
 wire \V3/V1/V1/A2/M4/s1 ;
 wire \V3/V1/V1/A3/c1 ;
 wire \V3/V1/V1/A3/c2 ;
 wire \V3/V1/V1/A3/c3 ;
 wire \V3/V1/V1/A3/M1/c1 ;
 wire \V3/V1/V1/A3/M1/c2 ;
 wire \V3/V1/V1/A3/M1/s1 ;
 wire \V3/V1/V1/A3/M2/c1 ;
 wire \V3/V1/V1/A3/M2/c2 ;
 wire \V3/V1/V1/A3/M2/s1 ;
 wire \V3/V1/V1/A3/M3/c1 ;
 wire \V3/V1/V1/A3/M3/c2 ;
 wire \V3/V1/V1/A3/M3/s1 ;
 wire \V3/V1/V1/A3/M4/c1 ;
 wire \V3/V1/V1/A3/M4/c2 ;
 wire \V3/V1/V1/A3/M4/s1 ;
 wire \V3/V1/V1/V1/w1 ;
 wire \V3/V1/V1/V1/w2 ;
 wire \V3/V1/V1/V1/w3 ;
 wire \V3/V1/V1/V1/w4 ;
 wire \V3/V1/V1/V2/w1 ;
 wire \V3/V1/V1/V2/w2 ;
 wire \V3/V1/V1/V2/w3 ;
 wire \V3/V1/V1/V2/w4 ;
 wire \V3/V1/V1/V3/w1 ;
 wire \V3/V1/V1/V3/w2 ;
 wire \V3/V1/V1/V3/w3 ;
 wire \V3/V1/V1/V3/w4 ;
 wire \V3/V1/V1/V4/w1 ;
 wire \V3/V1/V1/V4/w2 ;
 wire \V3/V1/V1/V4/w3 ;
 wire \V3/V1/V1/V4/w4 ;
 wire \V3/V1/V2/c1 ;
 wire \V3/V1/V2/c2 ;
 wire \V3/V1/V2/c3 ;
 wire \V3/V1/V2/overflow ;
 wire \V3/V1/V2/A1/c1 ;
 wire \V3/V1/V2/A1/c2 ;
 wire \V3/V1/V2/A1/c3 ;
 wire \V3/V1/V2/A1/M1/c1 ;
 wire \V3/V1/V2/A1/M1/c2 ;
 wire \V3/V1/V2/A1/M1/s1 ;
 wire \V3/V1/V2/A1/M2/c1 ;
 wire \V3/V1/V2/A1/M2/c2 ;
 wire \V3/V1/V2/A1/M2/s1 ;
 wire \V3/V1/V2/A1/M3/c1 ;
 wire \V3/V1/V2/A1/M3/c2 ;
 wire \V3/V1/V2/A1/M3/s1 ;
 wire \V3/V1/V2/A1/M4/c1 ;
 wire \V3/V1/V2/A1/M4/c2 ;
 wire \V3/V1/V2/A1/M4/s1 ;
 wire \V3/V1/V2/A2/c1 ;
 wire \V3/V1/V2/A2/c2 ;
 wire \V3/V1/V2/A2/c3 ;
 wire \V3/V1/V2/A2/M1/c1 ;
 wire \V3/V1/V2/A2/M1/c2 ;
 wire \V3/V1/V2/A2/M1/s1 ;
 wire \V3/V1/V2/A2/M2/c1 ;
 wire \V3/V1/V2/A2/M2/c2 ;
 wire \V3/V1/V2/A2/M2/s1 ;
 wire \V3/V1/V2/A2/M3/c1 ;
 wire \V3/V1/V2/A2/M3/c2 ;
 wire \V3/V1/V2/A2/M3/s1 ;
 wire \V3/V1/V2/A2/M4/c1 ;
 wire \V3/V1/V2/A2/M4/c2 ;
 wire \V3/V1/V2/A2/M4/s1 ;
 wire \V3/V1/V2/A3/c1 ;
 wire \V3/V1/V2/A3/c2 ;
 wire \V3/V1/V2/A3/c3 ;
 wire \V3/V1/V2/A3/M1/c1 ;
 wire \V3/V1/V2/A3/M1/c2 ;
 wire \V3/V1/V2/A3/M1/s1 ;
 wire \V3/V1/V2/A3/M2/c1 ;
 wire \V3/V1/V2/A3/M2/c2 ;
 wire \V3/V1/V2/A3/M2/s1 ;
 wire \V3/V1/V2/A3/M3/c1 ;
 wire \V3/V1/V2/A3/M3/c2 ;
 wire \V3/V1/V2/A3/M3/s1 ;
 wire \V3/V1/V2/A3/M4/c1 ;
 wire \V3/V1/V2/A3/M4/c2 ;
 wire \V3/V1/V2/A3/M4/s1 ;
 wire \V3/V1/V2/V1/w1 ;
 wire \V3/V1/V2/V1/w2 ;
 wire \V3/V1/V2/V1/w3 ;
 wire \V3/V1/V2/V1/w4 ;
 wire \V3/V1/V2/V2/w1 ;
 wire \V3/V1/V2/V2/w2 ;
 wire \V3/V1/V2/V2/w3 ;
 wire \V3/V1/V2/V2/w4 ;
 wire \V3/V1/V2/V3/w1 ;
 wire \V3/V1/V2/V3/w2 ;
 wire \V3/V1/V2/V3/w3 ;
 wire \V3/V1/V2/V3/w4 ;
 wire \V3/V1/V2/V4/w1 ;
 wire \V3/V1/V2/V4/w2 ;
 wire \V3/V1/V2/V4/w3 ;
 wire \V3/V1/V2/V4/w4 ;
 wire \V3/V1/V3/c1 ;
 wire \V3/V1/V3/c2 ;
 wire \V3/V1/V3/c3 ;
 wire \V3/V1/V3/overflow ;
 wire \V3/V1/V3/A1/c1 ;
 wire \V3/V1/V3/A1/c2 ;
 wire \V3/V1/V3/A1/c3 ;
 wire \V3/V1/V3/A1/M1/c1 ;
 wire \V3/V1/V3/A1/M1/c2 ;
 wire \V3/V1/V3/A1/M1/s1 ;
 wire \V3/V1/V3/A1/M2/c1 ;
 wire \V3/V1/V3/A1/M2/c2 ;
 wire \V3/V1/V3/A1/M2/s1 ;
 wire \V3/V1/V3/A1/M3/c1 ;
 wire \V3/V1/V3/A1/M3/c2 ;
 wire \V3/V1/V3/A1/M3/s1 ;
 wire \V3/V1/V3/A1/M4/c1 ;
 wire \V3/V1/V3/A1/M4/c2 ;
 wire \V3/V1/V3/A1/M4/s1 ;
 wire \V3/V1/V3/A2/c1 ;
 wire \V3/V1/V3/A2/c2 ;
 wire \V3/V1/V3/A2/c3 ;
 wire \V3/V1/V3/A2/M1/c1 ;
 wire \V3/V1/V3/A2/M1/c2 ;
 wire \V3/V1/V3/A2/M1/s1 ;
 wire \V3/V1/V3/A2/M2/c1 ;
 wire \V3/V1/V3/A2/M2/c2 ;
 wire \V3/V1/V3/A2/M2/s1 ;
 wire \V3/V1/V3/A2/M3/c1 ;
 wire \V3/V1/V3/A2/M3/c2 ;
 wire \V3/V1/V3/A2/M3/s1 ;
 wire \V3/V1/V3/A2/M4/c1 ;
 wire \V3/V1/V3/A2/M4/c2 ;
 wire \V3/V1/V3/A2/M4/s1 ;
 wire \V3/V1/V3/A3/c1 ;
 wire \V3/V1/V3/A3/c2 ;
 wire \V3/V1/V3/A3/c3 ;
 wire \V3/V1/V3/A3/M1/c1 ;
 wire \V3/V1/V3/A3/M1/c2 ;
 wire \V3/V1/V3/A3/M1/s1 ;
 wire \V3/V1/V3/A3/M2/c1 ;
 wire \V3/V1/V3/A3/M2/c2 ;
 wire \V3/V1/V3/A3/M2/s1 ;
 wire \V3/V1/V3/A3/M3/c1 ;
 wire \V3/V1/V3/A3/M3/c2 ;
 wire \V3/V1/V3/A3/M3/s1 ;
 wire \V3/V1/V3/A3/M4/c1 ;
 wire \V3/V1/V3/A3/M4/c2 ;
 wire \V3/V1/V3/A3/M4/s1 ;
 wire \V3/V1/V3/V1/w1 ;
 wire \V3/V1/V3/V1/w2 ;
 wire \V3/V1/V3/V1/w3 ;
 wire \V3/V1/V3/V1/w4 ;
 wire \V3/V1/V3/V2/w1 ;
 wire \V3/V1/V3/V2/w2 ;
 wire \V3/V1/V3/V2/w3 ;
 wire \V3/V1/V3/V2/w4 ;
 wire \V3/V1/V3/V3/w1 ;
 wire \V3/V1/V3/V3/w2 ;
 wire \V3/V1/V3/V3/w3 ;
 wire \V3/V1/V3/V3/w4 ;
 wire \V3/V1/V3/V4/w1 ;
 wire \V3/V1/V3/V4/w2 ;
 wire \V3/V1/V3/V4/w3 ;
 wire \V3/V1/V3/V4/w4 ;
 wire \V3/V1/V4/c1 ;
 wire \V3/V1/V4/c2 ;
 wire \V3/V1/V4/c3 ;
 wire \V3/V1/V4/overflow ;
 wire \V3/V1/V4/A1/c1 ;
 wire \V3/V1/V4/A1/c2 ;
 wire \V3/V1/V4/A1/c3 ;
 wire \V3/V1/V4/A1/M1/c1 ;
 wire \V3/V1/V4/A1/M1/c2 ;
 wire \V3/V1/V4/A1/M1/s1 ;
 wire \V3/V1/V4/A1/M2/c1 ;
 wire \V3/V1/V4/A1/M2/c2 ;
 wire \V3/V1/V4/A1/M2/s1 ;
 wire \V3/V1/V4/A1/M3/c1 ;
 wire \V3/V1/V4/A1/M3/c2 ;
 wire \V3/V1/V4/A1/M3/s1 ;
 wire \V3/V1/V4/A1/M4/c1 ;
 wire \V3/V1/V4/A1/M4/c2 ;
 wire \V3/V1/V4/A1/M4/s1 ;
 wire \V3/V1/V4/A2/c1 ;
 wire \V3/V1/V4/A2/c2 ;
 wire \V3/V1/V4/A2/c3 ;
 wire \V3/V1/V4/A2/M1/c1 ;
 wire \V3/V1/V4/A2/M1/c2 ;
 wire \V3/V1/V4/A2/M1/s1 ;
 wire \V3/V1/V4/A2/M2/c1 ;
 wire \V3/V1/V4/A2/M2/c2 ;
 wire \V3/V1/V4/A2/M2/s1 ;
 wire \V3/V1/V4/A2/M3/c1 ;
 wire \V3/V1/V4/A2/M3/c2 ;
 wire \V3/V1/V4/A2/M3/s1 ;
 wire \V3/V1/V4/A2/M4/c1 ;
 wire \V3/V1/V4/A2/M4/c2 ;
 wire \V3/V1/V4/A2/M4/s1 ;
 wire \V3/V1/V4/A3/c1 ;
 wire \V3/V1/V4/A3/c2 ;
 wire \V3/V1/V4/A3/c3 ;
 wire \V3/V1/V4/A3/M1/c1 ;
 wire \V3/V1/V4/A3/M1/c2 ;
 wire \V3/V1/V4/A3/M1/s1 ;
 wire \V3/V1/V4/A3/M2/c1 ;
 wire \V3/V1/V4/A3/M2/c2 ;
 wire \V3/V1/V4/A3/M2/s1 ;
 wire \V3/V1/V4/A3/M3/c1 ;
 wire \V3/V1/V4/A3/M3/c2 ;
 wire \V3/V1/V4/A3/M3/s1 ;
 wire \V3/V1/V4/A3/M4/c1 ;
 wire \V3/V1/V4/A3/M4/c2 ;
 wire \V3/V1/V4/A3/M4/s1 ;
 wire \V3/V1/V4/V1/w1 ;
 wire \V3/V1/V4/V1/w2 ;
 wire \V3/V1/V4/V1/w3 ;
 wire \V3/V1/V4/V1/w4 ;
 wire \V3/V1/V4/V2/w1 ;
 wire \V3/V1/V4/V2/w2 ;
 wire \V3/V1/V4/V2/w3 ;
 wire \V3/V1/V4/V2/w4 ;
 wire \V3/V1/V4/V3/w1 ;
 wire \V3/V1/V4/V3/w2 ;
 wire \V3/V1/V4/V3/w3 ;
 wire \V3/V1/V4/V3/w4 ;
 wire \V3/V1/V4/V4/w1 ;
 wire \V3/V1/V4/V4/w2 ;
 wire \V3/V1/V4/V4/w3 ;
 wire \V3/V1/V4/V4/w4 ;
 wire \V3/V2/c1 ;
 wire \V3/V2/c2 ;
 wire \V3/V2/c3 ;
 wire \V3/V2/overflow ;
 wire \V3/V2/A1/c1 ;
 wire \V3/V2/A1/A1/c1 ;
 wire \V3/V2/A1/A1/c2 ;
 wire \V3/V2/A1/A1/c3 ;
 wire \V3/V2/A1/A1/M1/c1 ;
 wire \V3/V2/A1/A1/M1/c2 ;
 wire \V3/V2/A1/A1/M1/s1 ;
 wire \V3/V2/A1/A1/M2/c1 ;
 wire \V3/V2/A1/A1/M2/c2 ;
 wire \V3/V2/A1/A1/M2/s1 ;
 wire \V3/V2/A1/A1/M3/c1 ;
 wire \V3/V2/A1/A1/M3/c2 ;
 wire \V3/V2/A1/A1/M3/s1 ;
 wire \V3/V2/A1/A1/M4/c1 ;
 wire \V3/V2/A1/A1/M4/c2 ;
 wire \V3/V2/A1/A1/M4/s1 ;
 wire \V3/V2/A1/A2/c1 ;
 wire \V3/V2/A1/A2/c2 ;
 wire \V3/V2/A1/A2/c3 ;
 wire \V3/V2/A1/A2/M1/c1 ;
 wire \V3/V2/A1/A2/M1/c2 ;
 wire \V3/V2/A1/A2/M1/s1 ;
 wire \V3/V2/A1/A2/M2/c1 ;
 wire \V3/V2/A1/A2/M2/c2 ;
 wire \V3/V2/A1/A2/M2/s1 ;
 wire \V3/V2/A1/A2/M3/c1 ;
 wire \V3/V2/A1/A2/M3/c2 ;
 wire \V3/V2/A1/A2/M3/s1 ;
 wire \V3/V2/A1/A2/M4/c1 ;
 wire \V3/V2/A1/A2/M4/c2 ;
 wire \V3/V2/A1/A2/M4/s1 ;
 wire \V3/V2/A2/c1 ;
 wire \V3/V2/A2/A1/c1 ;
 wire \V3/V2/A2/A1/c2 ;
 wire \V3/V2/A2/A1/c3 ;
 wire \V3/V2/A2/A1/M1/c1 ;
 wire \V3/V2/A2/A1/M1/c2 ;
 wire \V3/V2/A2/A1/M1/s1 ;
 wire \V3/V2/A2/A1/M2/c1 ;
 wire \V3/V2/A2/A1/M2/c2 ;
 wire \V3/V2/A2/A1/M2/s1 ;
 wire \V3/V2/A2/A1/M3/c1 ;
 wire \V3/V2/A2/A1/M3/c2 ;
 wire \V3/V2/A2/A1/M3/s1 ;
 wire \V3/V2/A2/A1/M4/c1 ;
 wire \V3/V2/A2/A1/M4/c2 ;
 wire \V3/V2/A2/A1/M4/s1 ;
 wire \V3/V2/A2/A2/c1 ;
 wire \V3/V2/A2/A2/c2 ;
 wire \V3/V2/A2/A2/c3 ;
 wire \V3/V2/A2/A2/M1/c1 ;
 wire \V3/V2/A2/A2/M1/c2 ;
 wire \V3/V2/A2/A2/M1/s1 ;
 wire \V3/V2/A2/A2/M2/c1 ;
 wire \V3/V2/A2/A2/M2/c2 ;
 wire \V3/V2/A2/A2/M2/s1 ;
 wire \V3/V2/A2/A2/M3/c1 ;
 wire \V3/V2/A2/A2/M3/c2 ;
 wire \V3/V2/A2/A2/M3/s1 ;
 wire \V3/V2/A2/A2/M4/c1 ;
 wire \V3/V2/A2/A2/M4/c2 ;
 wire \V3/V2/A2/A2/M4/s1 ;
 wire \V3/V2/A3/c1 ;
 wire \V3/V2/A3/A1/c1 ;
 wire \V3/V2/A3/A1/c2 ;
 wire \V3/V2/A3/A1/c3 ;
 wire \V3/V2/A3/A1/M1/c1 ;
 wire \V3/V2/A3/A1/M1/c2 ;
 wire \V3/V2/A3/A1/M1/s1 ;
 wire \V3/V2/A3/A1/M2/c1 ;
 wire \V3/V2/A3/A1/M2/c2 ;
 wire \V3/V2/A3/A1/M2/s1 ;
 wire \V3/V2/A3/A1/M3/c1 ;
 wire \V3/V2/A3/A1/M3/c2 ;
 wire \V3/V2/A3/A1/M3/s1 ;
 wire \V3/V2/A3/A1/M4/c1 ;
 wire \V3/V2/A3/A1/M4/c2 ;
 wire \V3/V2/A3/A1/M4/s1 ;
 wire \V3/V2/A3/A2/c1 ;
 wire \V3/V2/A3/A2/c2 ;
 wire \V3/V2/A3/A2/c3 ;
 wire \V3/V2/A3/A2/M1/c1 ;
 wire \V3/V2/A3/A2/M1/c2 ;
 wire \V3/V2/A3/A2/M1/s1 ;
 wire \V3/V2/A3/A2/M2/c1 ;
 wire \V3/V2/A3/A2/M2/c2 ;
 wire \V3/V2/A3/A2/M2/s1 ;
 wire \V3/V2/A3/A2/M3/c1 ;
 wire \V3/V2/A3/A2/M3/c2 ;
 wire \V3/V2/A3/A2/M3/s1 ;
 wire \V3/V2/A3/A2/M4/c1 ;
 wire \V3/V2/A3/A2/M4/c2 ;
 wire \V3/V2/A3/A2/M4/s1 ;
 wire \V3/V2/V1/c1 ;
 wire \V3/V2/V1/c2 ;
 wire \V3/V2/V1/c3 ;
 wire \V3/V2/V1/overflow ;
 wire \V3/V2/V1/A1/c1 ;
 wire \V3/V2/V1/A1/c2 ;
 wire \V3/V2/V1/A1/c3 ;
 wire \V3/V2/V1/A1/M1/c1 ;
 wire \V3/V2/V1/A1/M1/c2 ;
 wire \V3/V2/V1/A1/M1/s1 ;
 wire \V3/V2/V1/A1/M2/c1 ;
 wire \V3/V2/V1/A1/M2/c2 ;
 wire \V3/V2/V1/A1/M2/s1 ;
 wire \V3/V2/V1/A1/M3/c1 ;
 wire \V3/V2/V1/A1/M3/c2 ;
 wire \V3/V2/V1/A1/M3/s1 ;
 wire \V3/V2/V1/A1/M4/c1 ;
 wire \V3/V2/V1/A1/M4/c2 ;
 wire \V3/V2/V1/A1/M4/s1 ;
 wire \V3/V2/V1/A2/c1 ;
 wire \V3/V2/V1/A2/c2 ;
 wire \V3/V2/V1/A2/c3 ;
 wire \V3/V2/V1/A2/M1/c1 ;
 wire \V3/V2/V1/A2/M1/c2 ;
 wire \V3/V2/V1/A2/M1/s1 ;
 wire \V3/V2/V1/A2/M2/c1 ;
 wire \V3/V2/V1/A2/M2/c2 ;
 wire \V3/V2/V1/A2/M2/s1 ;
 wire \V3/V2/V1/A2/M3/c1 ;
 wire \V3/V2/V1/A2/M3/c2 ;
 wire \V3/V2/V1/A2/M3/s1 ;
 wire \V3/V2/V1/A2/M4/c1 ;
 wire \V3/V2/V1/A2/M4/c2 ;
 wire \V3/V2/V1/A2/M4/s1 ;
 wire \V3/V2/V1/A3/c1 ;
 wire \V3/V2/V1/A3/c2 ;
 wire \V3/V2/V1/A3/c3 ;
 wire \V3/V2/V1/A3/M1/c1 ;
 wire \V3/V2/V1/A3/M1/c2 ;
 wire \V3/V2/V1/A3/M1/s1 ;
 wire \V3/V2/V1/A3/M2/c1 ;
 wire \V3/V2/V1/A3/M2/c2 ;
 wire \V3/V2/V1/A3/M2/s1 ;
 wire \V3/V2/V1/A3/M3/c1 ;
 wire \V3/V2/V1/A3/M3/c2 ;
 wire \V3/V2/V1/A3/M3/s1 ;
 wire \V3/V2/V1/A3/M4/c1 ;
 wire \V3/V2/V1/A3/M4/c2 ;
 wire \V3/V2/V1/A3/M4/s1 ;
 wire \V3/V2/V1/V1/w1 ;
 wire \V3/V2/V1/V1/w2 ;
 wire \V3/V2/V1/V1/w3 ;
 wire \V3/V2/V1/V1/w4 ;
 wire \V3/V2/V1/V2/w1 ;
 wire \V3/V2/V1/V2/w2 ;
 wire \V3/V2/V1/V2/w3 ;
 wire \V3/V2/V1/V2/w4 ;
 wire \V3/V2/V1/V3/w1 ;
 wire \V3/V2/V1/V3/w2 ;
 wire \V3/V2/V1/V3/w3 ;
 wire \V3/V2/V1/V3/w4 ;
 wire \V3/V2/V1/V4/w1 ;
 wire \V3/V2/V1/V4/w2 ;
 wire \V3/V2/V1/V4/w3 ;
 wire \V3/V2/V1/V4/w4 ;
 wire \V3/V2/V2/c1 ;
 wire \V3/V2/V2/c2 ;
 wire \V3/V2/V2/c3 ;
 wire \V3/V2/V2/overflow ;
 wire \V3/V2/V2/A1/c1 ;
 wire \V3/V2/V2/A1/c2 ;
 wire \V3/V2/V2/A1/c3 ;
 wire \V3/V2/V2/A1/M1/c1 ;
 wire \V3/V2/V2/A1/M1/c2 ;
 wire \V3/V2/V2/A1/M1/s1 ;
 wire \V3/V2/V2/A1/M2/c1 ;
 wire \V3/V2/V2/A1/M2/c2 ;
 wire \V3/V2/V2/A1/M2/s1 ;
 wire \V3/V2/V2/A1/M3/c1 ;
 wire \V3/V2/V2/A1/M3/c2 ;
 wire \V3/V2/V2/A1/M3/s1 ;
 wire \V3/V2/V2/A1/M4/c1 ;
 wire \V3/V2/V2/A1/M4/c2 ;
 wire \V3/V2/V2/A1/M4/s1 ;
 wire \V3/V2/V2/A2/c1 ;
 wire \V3/V2/V2/A2/c2 ;
 wire \V3/V2/V2/A2/c3 ;
 wire \V3/V2/V2/A2/M1/c1 ;
 wire \V3/V2/V2/A2/M1/c2 ;
 wire \V3/V2/V2/A2/M1/s1 ;
 wire \V3/V2/V2/A2/M2/c1 ;
 wire \V3/V2/V2/A2/M2/c2 ;
 wire \V3/V2/V2/A2/M2/s1 ;
 wire \V3/V2/V2/A2/M3/c1 ;
 wire \V3/V2/V2/A2/M3/c2 ;
 wire \V3/V2/V2/A2/M3/s1 ;
 wire \V3/V2/V2/A2/M4/c1 ;
 wire \V3/V2/V2/A2/M4/c2 ;
 wire \V3/V2/V2/A2/M4/s1 ;
 wire \V3/V2/V2/A3/c1 ;
 wire \V3/V2/V2/A3/c2 ;
 wire \V3/V2/V2/A3/c3 ;
 wire \V3/V2/V2/A3/M1/c1 ;
 wire \V3/V2/V2/A3/M1/c2 ;
 wire \V3/V2/V2/A3/M1/s1 ;
 wire \V3/V2/V2/A3/M2/c1 ;
 wire \V3/V2/V2/A3/M2/c2 ;
 wire \V3/V2/V2/A3/M2/s1 ;
 wire \V3/V2/V2/A3/M3/c1 ;
 wire \V3/V2/V2/A3/M3/c2 ;
 wire \V3/V2/V2/A3/M3/s1 ;
 wire \V3/V2/V2/A3/M4/c1 ;
 wire \V3/V2/V2/A3/M4/c2 ;
 wire \V3/V2/V2/A3/M4/s1 ;
 wire \V3/V2/V2/V1/w1 ;
 wire \V3/V2/V2/V1/w2 ;
 wire \V3/V2/V2/V1/w3 ;
 wire \V3/V2/V2/V1/w4 ;
 wire \V3/V2/V2/V2/w1 ;
 wire \V3/V2/V2/V2/w2 ;
 wire \V3/V2/V2/V2/w3 ;
 wire \V3/V2/V2/V2/w4 ;
 wire \V3/V2/V2/V3/w1 ;
 wire \V3/V2/V2/V3/w2 ;
 wire \V3/V2/V2/V3/w3 ;
 wire \V3/V2/V2/V3/w4 ;
 wire \V3/V2/V2/V4/w1 ;
 wire \V3/V2/V2/V4/w2 ;
 wire \V3/V2/V2/V4/w3 ;
 wire \V3/V2/V2/V4/w4 ;
 wire \V3/V2/V3/c1 ;
 wire \V3/V2/V3/c2 ;
 wire \V3/V2/V3/c3 ;
 wire \V3/V2/V3/overflow ;
 wire \V3/V2/V3/A1/c1 ;
 wire \V3/V2/V3/A1/c2 ;
 wire \V3/V2/V3/A1/c3 ;
 wire \V3/V2/V3/A1/M1/c1 ;
 wire \V3/V2/V3/A1/M1/c2 ;
 wire \V3/V2/V3/A1/M1/s1 ;
 wire \V3/V2/V3/A1/M2/c1 ;
 wire \V3/V2/V3/A1/M2/c2 ;
 wire \V3/V2/V3/A1/M2/s1 ;
 wire \V3/V2/V3/A1/M3/c1 ;
 wire \V3/V2/V3/A1/M3/c2 ;
 wire \V3/V2/V3/A1/M3/s1 ;
 wire \V3/V2/V3/A1/M4/c1 ;
 wire \V3/V2/V3/A1/M4/c2 ;
 wire \V3/V2/V3/A1/M4/s1 ;
 wire \V3/V2/V3/A2/c1 ;
 wire \V3/V2/V3/A2/c2 ;
 wire \V3/V2/V3/A2/c3 ;
 wire \V3/V2/V3/A2/M1/c1 ;
 wire \V3/V2/V3/A2/M1/c2 ;
 wire \V3/V2/V3/A2/M1/s1 ;
 wire \V3/V2/V3/A2/M2/c1 ;
 wire \V3/V2/V3/A2/M2/c2 ;
 wire \V3/V2/V3/A2/M2/s1 ;
 wire \V3/V2/V3/A2/M3/c1 ;
 wire \V3/V2/V3/A2/M3/c2 ;
 wire \V3/V2/V3/A2/M3/s1 ;
 wire \V3/V2/V3/A2/M4/c1 ;
 wire \V3/V2/V3/A2/M4/c2 ;
 wire \V3/V2/V3/A2/M4/s1 ;
 wire \V3/V2/V3/A3/c1 ;
 wire \V3/V2/V3/A3/c2 ;
 wire \V3/V2/V3/A3/c3 ;
 wire \V3/V2/V3/A3/M1/c1 ;
 wire \V3/V2/V3/A3/M1/c2 ;
 wire \V3/V2/V3/A3/M1/s1 ;
 wire \V3/V2/V3/A3/M2/c1 ;
 wire \V3/V2/V3/A3/M2/c2 ;
 wire \V3/V2/V3/A3/M2/s1 ;
 wire \V3/V2/V3/A3/M3/c1 ;
 wire \V3/V2/V3/A3/M3/c2 ;
 wire \V3/V2/V3/A3/M3/s1 ;
 wire \V3/V2/V3/A3/M4/c1 ;
 wire \V3/V2/V3/A3/M4/c2 ;
 wire \V3/V2/V3/A3/M4/s1 ;
 wire \V3/V2/V3/V1/w1 ;
 wire \V3/V2/V3/V1/w2 ;
 wire \V3/V2/V3/V1/w3 ;
 wire \V3/V2/V3/V1/w4 ;
 wire \V3/V2/V3/V2/w1 ;
 wire \V3/V2/V3/V2/w2 ;
 wire \V3/V2/V3/V2/w3 ;
 wire \V3/V2/V3/V2/w4 ;
 wire \V3/V2/V3/V3/w1 ;
 wire \V3/V2/V3/V3/w2 ;
 wire \V3/V2/V3/V3/w3 ;
 wire \V3/V2/V3/V3/w4 ;
 wire \V3/V2/V3/V4/w1 ;
 wire \V3/V2/V3/V4/w2 ;
 wire \V3/V2/V3/V4/w3 ;
 wire \V3/V2/V3/V4/w4 ;
 wire \V3/V2/V4/c1 ;
 wire \V3/V2/V4/c2 ;
 wire \V3/V2/V4/c3 ;
 wire \V3/V2/V4/overflow ;
 wire \V3/V2/V4/A1/c1 ;
 wire \V3/V2/V4/A1/c2 ;
 wire \V3/V2/V4/A1/c3 ;
 wire \V3/V2/V4/A1/M1/c1 ;
 wire \V3/V2/V4/A1/M1/c2 ;
 wire \V3/V2/V4/A1/M1/s1 ;
 wire \V3/V2/V4/A1/M2/c1 ;
 wire \V3/V2/V4/A1/M2/c2 ;
 wire \V3/V2/V4/A1/M2/s1 ;
 wire \V3/V2/V4/A1/M3/c1 ;
 wire \V3/V2/V4/A1/M3/c2 ;
 wire \V3/V2/V4/A1/M3/s1 ;
 wire \V3/V2/V4/A1/M4/c1 ;
 wire \V3/V2/V4/A1/M4/c2 ;
 wire \V3/V2/V4/A1/M4/s1 ;
 wire \V3/V2/V4/A2/c1 ;
 wire \V3/V2/V4/A2/c2 ;
 wire \V3/V2/V4/A2/c3 ;
 wire \V3/V2/V4/A2/M1/c1 ;
 wire \V3/V2/V4/A2/M1/c2 ;
 wire \V3/V2/V4/A2/M1/s1 ;
 wire \V3/V2/V4/A2/M2/c1 ;
 wire \V3/V2/V4/A2/M2/c2 ;
 wire \V3/V2/V4/A2/M2/s1 ;
 wire \V3/V2/V4/A2/M3/c1 ;
 wire \V3/V2/V4/A2/M3/c2 ;
 wire \V3/V2/V4/A2/M3/s1 ;
 wire \V3/V2/V4/A2/M4/c1 ;
 wire \V3/V2/V4/A2/M4/c2 ;
 wire \V3/V2/V4/A2/M4/s1 ;
 wire \V3/V2/V4/A3/c1 ;
 wire \V3/V2/V4/A3/c2 ;
 wire \V3/V2/V4/A3/c3 ;
 wire \V3/V2/V4/A3/M1/c1 ;
 wire \V3/V2/V4/A3/M1/c2 ;
 wire \V3/V2/V4/A3/M1/s1 ;
 wire \V3/V2/V4/A3/M2/c1 ;
 wire \V3/V2/V4/A3/M2/c2 ;
 wire \V3/V2/V4/A3/M2/s1 ;
 wire \V3/V2/V4/A3/M3/c1 ;
 wire \V3/V2/V4/A3/M3/c2 ;
 wire \V3/V2/V4/A3/M3/s1 ;
 wire \V3/V2/V4/A3/M4/c1 ;
 wire \V3/V2/V4/A3/M4/c2 ;
 wire \V3/V2/V4/A3/M4/s1 ;
 wire \V3/V2/V4/V1/w1 ;
 wire \V3/V2/V4/V1/w2 ;
 wire \V3/V2/V4/V1/w3 ;
 wire \V3/V2/V4/V1/w4 ;
 wire \V3/V2/V4/V2/w1 ;
 wire \V3/V2/V4/V2/w2 ;
 wire \V3/V2/V4/V2/w3 ;
 wire \V3/V2/V4/V2/w4 ;
 wire \V3/V2/V4/V3/w1 ;
 wire \V3/V2/V4/V3/w2 ;
 wire \V3/V2/V4/V3/w3 ;
 wire \V3/V2/V4/V3/w4 ;
 wire \V3/V2/V4/V4/w1 ;
 wire \V3/V2/V4/V4/w2 ;
 wire \V3/V2/V4/V4/w3 ;
 wire \V3/V2/V4/V4/w4 ;
 wire \V3/V3/c1 ;
 wire \V3/V3/c2 ;
 wire \V3/V3/c3 ;
 wire \V3/V3/overflow ;
 wire \V3/V3/A1/c1 ;
 wire \V3/V3/A1/A1/c1 ;
 wire \V3/V3/A1/A1/c2 ;
 wire \V3/V3/A1/A1/c3 ;
 wire \V3/V3/A1/A1/M1/c1 ;
 wire \V3/V3/A1/A1/M1/c2 ;
 wire \V3/V3/A1/A1/M1/s1 ;
 wire \V3/V3/A1/A1/M2/c1 ;
 wire \V3/V3/A1/A1/M2/c2 ;
 wire \V3/V3/A1/A1/M2/s1 ;
 wire \V3/V3/A1/A1/M3/c1 ;
 wire \V3/V3/A1/A1/M3/c2 ;
 wire \V3/V3/A1/A1/M3/s1 ;
 wire \V3/V3/A1/A1/M4/c1 ;
 wire \V3/V3/A1/A1/M4/c2 ;
 wire \V3/V3/A1/A1/M4/s1 ;
 wire \V3/V3/A1/A2/c1 ;
 wire \V3/V3/A1/A2/c2 ;
 wire \V3/V3/A1/A2/c3 ;
 wire \V3/V3/A1/A2/M1/c1 ;
 wire \V3/V3/A1/A2/M1/c2 ;
 wire \V3/V3/A1/A2/M1/s1 ;
 wire \V3/V3/A1/A2/M2/c1 ;
 wire \V3/V3/A1/A2/M2/c2 ;
 wire \V3/V3/A1/A2/M2/s1 ;
 wire \V3/V3/A1/A2/M3/c1 ;
 wire \V3/V3/A1/A2/M3/c2 ;
 wire \V3/V3/A1/A2/M3/s1 ;
 wire \V3/V3/A1/A2/M4/c1 ;
 wire \V3/V3/A1/A2/M4/c2 ;
 wire \V3/V3/A1/A2/M4/s1 ;
 wire \V3/V3/A2/c1 ;
 wire \V3/V3/A2/A1/c1 ;
 wire \V3/V3/A2/A1/c2 ;
 wire \V3/V3/A2/A1/c3 ;
 wire \V3/V3/A2/A1/M1/c1 ;
 wire \V3/V3/A2/A1/M1/c2 ;
 wire \V3/V3/A2/A1/M1/s1 ;
 wire \V3/V3/A2/A1/M2/c1 ;
 wire \V3/V3/A2/A1/M2/c2 ;
 wire \V3/V3/A2/A1/M2/s1 ;
 wire \V3/V3/A2/A1/M3/c1 ;
 wire \V3/V3/A2/A1/M3/c2 ;
 wire \V3/V3/A2/A1/M3/s1 ;
 wire \V3/V3/A2/A1/M4/c1 ;
 wire \V3/V3/A2/A1/M4/c2 ;
 wire \V3/V3/A2/A1/M4/s1 ;
 wire \V3/V3/A2/A2/c1 ;
 wire \V3/V3/A2/A2/c2 ;
 wire \V3/V3/A2/A2/c3 ;
 wire \V3/V3/A2/A2/M1/c1 ;
 wire \V3/V3/A2/A2/M1/c2 ;
 wire \V3/V3/A2/A2/M1/s1 ;
 wire \V3/V3/A2/A2/M2/c1 ;
 wire \V3/V3/A2/A2/M2/c2 ;
 wire \V3/V3/A2/A2/M2/s1 ;
 wire \V3/V3/A2/A2/M3/c1 ;
 wire \V3/V3/A2/A2/M3/c2 ;
 wire \V3/V3/A2/A2/M3/s1 ;
 wire \V3/V3/A2/A2/M4/c1 ;
 wire \V3/V3/A2/A2/M4/c2 ;
 wire \V3/V3/A2/A2/M4/s1 ;
 wire \V3/V3/A3/c1 ;
 wire \V3/V3/A3/A1/c1 ;
 wire \V3/V3/A3/A1/c2 ;
 wire \V3/V3/A3/A1/c3 ;
 wire \V3/V3/A3/A1/M1/c1 ;
 wire \V3/V3/A3/A1/M1/c2 ;
 wire \V3/V3/A3/A1/M1/s1 ;
 wire \V3/V3/A3/A1/M2/c1 ;
 wire \V3/V3/A3/A1/M2/c2 ;
 wire \V3/V3/A3/A1/M2/s1 ;
 wire \V3/V3/A3/A1/M3/c1 ;
 wire \V3/V3/A3/A1/M3/c2 ;
 wire \V3/V3/A3/A1/M3/s1 ;
 wire \V3/V3/A3/A1/M4/c1 ;
 wire \V3/V3/A3/A1/M4/c2 ;
 wire \V3/V3/A3/A1/M4/s1 ;
 wire \V3/V3/A3/A2/c1 ;
 wire \V3/V3/A3/A2/c2 ;
 wire \V3/V3/A3/A2/c3 ;
 wire \V3/V3/A3/A2/M1/c1 ;
 wire \V3/V3/A3/A2/M1/c2 ;
 wire \V3/V3/A3/A2/M1/s1 ;
 wire \V3/V3/A3/A2/M2/c1 ;
 wire \V3/V3/A3/A2/M2/c2 ;
 wire \V3/V3/A3/A2/M2/s1 ;
 wire \V3/V3/A3/A2/M3/c1 ;
 wire \V3/V3/A3/A2/M3/c2 ;
 wire \V3/V3/A3/A2/M3/s1 ;
 wire \V3/V3/A3/A2/M4/c1 ;
 wire \V3/V3/A3/A2/M4/c2 ;
 wire \V3/V3/A3/A2/M4/s1 ;
 wire \V3/V3/V1/c1 ;
 wire \V3/V3/V1/c2 ;
 wire \V3/V3/V1/c3 ;
 wire \V3/V3/V1/overflow ;
 wire \V3/V3/V1/A1/c1 ;
 wire \V3/V3/V1/A1/c2 ;
 wire \V3/V3/V1/A1/c3 ;
 wire \V3/V3/V1/A1/M1/c1 ;
 wire \V3/V3/V1/A1/M1/c2 ;
 wire \V3/V3/V1/A1/M1/s1 ;
 wire \V3/V3/V1/A1/M2/c1 ;
 wire \V3/V3/V1/A1/M2/c2 ;
 wire \V3/V3/V1/A1/M2/s1 ;
 wire \V3/V3/V1/A1/M3/c1 ;
 wire \V3/V3/V1/A1/M3/c2 ;
 wire \V3/V3/V1/A1/M3/s1 ;
 wire \V3/V3/V1/A1/M4/c1 ;
 wire \V3/V3/V1/A1/M4/c2 ;
 wire \V3/V3/V1/A1/M4/s1 ;
 wire \V3/V3/V1/A2/c1 ;
 wire \V3/V3/V1/A2/c2 ;
 wire \V3/V3/V1/A2/c3 ;
 wire \V3/V3/V1/A2/M1/c1 ;
 wire \V3/V3/V1/A2/M1/c2 ;
 wire \V3/V3/V1/A2/M1/s1 ;
 wire \V3/V3/V1/A2/M2/c1 ;
 wire \V3/V3/V1/A2/M2/c2 ;
 wire \V3/V3/V1/A2/M2/s1 ;
 wire \V3/V3/V1/A2/M3/c1 ;
 wire \V3/V3/V1/A2/M3/c2 ;
 wire \V3/V3/V1/A2/M3/s1 ;
 wire \V3/V3/V1/A2/M4/c1 ;
 wire \V3/V3/V1/A2/M4/c2 ;
 wire \V3/V3/V1/A2/M4/s1 ;
 wire \V3/V3/V1/A3/c1 ;
 wire \V3/V3/V1/A3/c2 ;
 wire \V3/V3/V1/A3/c3 ;
 wire \V3/V3/V1/A3/M1/c1 ;
 wire \V3/V3/V1/A3/M1/c2 ;
 wire \V3/V3/V1/A3/M1/s1 ;
 wire \V3/V3/V1/A3/M2/c1 ;
 wire \V3/V3/V1/A3/M2/c2 ;
 wire \V3/V3/V1/A3/M2/s1 ;
 wire \V3/V3/V1/A3/M3/c1 ;
 wire \V3/V3/V1/A3/M3/c2 ;
 wire \V3/V3/V1/A3/M3/s1 ;
 wire \V3/V3/V1/A3/M4/c1 ;
 wire \V3/V3/V1/A3/M4/c2 ;
 wire \V3/V3/V1/A3/M4/s1 ;
 wire \V3/V3/V1/V1/w1 ;
 wire \V3/V3/V1/V1/w2 ;
 wire \V3/V3/V1/V1/w3 ;
 wire \V3/V3/V1/V1/w4 ;
 wire \V3/V3/V1/V2/w1 ;
 wire \V3/V3/V1/V2/w2 ;
 wire \V3/V3/V1/V2/w3 ;
 wire \V3/V3/V1/V2/w4 ;
 wire \V3/V3/V1/V3/w1 ;
 wire \V3/V3/V1/V3/w2 ;
 wire \V3/V3/V1/V3/w3 ;
 wire \V3/V3/V1/V3/w4 ;
 wire \V3/V3/V1/V4/w1 ;
 wire \V3/V3/V1/V4/w2 ;
 wire \V3/V3/V1/V4/w3 ;
 wire \V3/V3/V1/V4/w4 ;
 wire \V3/V3/V2/c1 ;
 wire \V3/V3/V2/c2 ;
 wire \V3/V3/V2/c3 ;
 wire \V3/V3/V2/overflow ;
 wire \V3/V3/V2/A1/c1 ;
 wire \V3/V3/V2/A1/c2 ;
 wire \V3/V3/V2/A1/c3 ;
 wire \V3/V3/V2/A1/M1/c1 ;
 wire \V3/V3/V2/A1/M1/c2 ;
 wire \V3/V3/V2/A1/M1/s1 ;
 wire \V3/V3/V2/A1/M2/c1 ;
 wire \V3/V3/V2/A1/M2/c2 ;
 wire \V3/V3/V2/A1/M2/s1 ;
 wire \V3/V3/V2/A1/M3/c1 ;
 wire \V3/V3/V2/A1/M3/c2 ;
 wire \V3/V3/V2/A1/M3/s1 ;
 wire \V3/V3/V2/A1/M4/c1 ;
 wire \V3/V3/V2/A1/M4/c2 ;
 wire \V3/V3/V2/A1/M4/s1 ;
 wire \V3/V3/V2/A2/c1 ;
 wire \V3/V3/V2/A2/c2 ;
 wire \V3/V3/V2/A2/c3 ;
 wire \V3/V3/V2/A2/M1/c1 ;
 wire \V3/V3/V2/A2/M1/c2 ;
 wire \V3/V3/V2/A2/M1/s1 ;
 wire \V3/V3/V2/A2/M2/c1 ;
 wire \V3/V3/V2/A2/M2/c2 ;
 wire \V3/V3/V2/A2/M2/s1 ;
 wire \V3/V3/V2/A2/M3/c1 ;
 wire \V3/V3/V2/A2/M3/c2 ;
 wire \V3/V3/V2/A2/M3/s1 ;
 wire \V3/V3/V2/A2/M4/c1 ;
 wire \V3/V3/V2/A2/M4/c2 ;
 wire \V3/V3/V2/A2/M4/s1 ;
 wire \V3/V3/V2/A3/c1 ;
 wire \V3/V3/V2/A3/c2 ;
 wire \V3/V3/V2/A3/c3 ;
 wire \V3/V3/V2/A3/M1/c1 ;
 wire \V3/V3/V2/A3/M1/c2 ;
 wire \V3/V3/V2/A3/M1/s1 ;
 wire \V3/V3/V2/A3/M2/c1 ;
 wire \V3/V3/V2/A3/M2/c2 ;
 wire \V3/V3/V2/A3/M2/s1 ;
 wire \V3/V3/V2/A3/M3/c1 ;
 wire \V3/V3/V2/A3/M3/c2 ;
 wire \V3/V3/V2/A3/M3/s1 ;
 wire \V3/V3/V2/A3/M4/c1 ;
 wire \V3/V3/V2/A3/M4/c2 ;
 wire \V3/V3/V2/A3/M4/s1 ;
 wire \V3/V3/V2/V1/w1 ;
 wire \V3/V3/V2/V1/w2 ;
 wire \V3/V3/V2/V1/w3 ;
 wire \V3/V3/V2/V1/w4 ;
 wire \V3/V3/V2/V2/w1 ;
 wire \V3/V3/V2/V2/w2 ;
 wire \V3/V3/V2/V2/w3 ;
 wire \V3/V3/V2/V2/w4 ;
 wire \V3/V3/V2/V3/w1 ;
 wire \V3/V3/V2/V3/w2 ;
 wire \V3/V3/V2/V3/w3 ;
 wire \V3/V3/V2/V3/w4 ;
 wire \V3/V3/V2/V4/w1 ;
 wire \V3/V3/V2/V4/w2 ;
 wire \V3/V3/V2/V4/w3 ;
 wire \V3/V3/V2/V4/w4 ;
 wire \V3/V3/V3/c1 ;
 wire \V3/V3/V3/c2 ;
 wire \V3/V3/V3/c3 ;
 wire \V3/V3/V3/overflow ;
 wire \V3/V3/V3/A1/c1 ;
 wire \V3/V3/V3/A1/c2 ;
 wire \V3/V3/V3/A1/c3 ;
 wire \V3/V3/V3/A1/M1/c1 ;
 wire \V3/V3/V3/A1/M1/c2 ;
 wire \V3/V3/V3/A1/M1/s1 ;
 wire \V3/V3/V3/A1/M2/c1 ;
 wire \V3/V3/V3/A1/M2/c2 ;
 wire \V3/V3/V3/A1/M2/s1 ;
 wire \V3/V3/V3/A1/M3/c1 ;
 wire \V3/V3/V3/A1/M3/c2 ;
 wire \V3/V3/V3/A1/M3/s1 ;
 wire \V3/V3/V3/A1/M4/c1 ;
 wire \V3/V3/V3/A1/M4/c2 ;
 wire \V3/V3/V3/A1/M4/s1 ;
 wire \V3/V3/V3/A2/c1 ;
 wire \V3/V3/V3/A2/c2 ;
 wire \V3/V3/V3/A2/c3 ;
 wire \V3/V3/V3/A2/M1/c1 ;
 wire \V3/V3/V3/A2/M1/c2 ;
 wire \V3/V3/V3/A2/M1/s1 ;
 wire \V3/V3/V3/A2/M2/c1 ;
 wire \V3/V3/V3/A2/M2/c2 ;
 wire \V3/V3/V3/A2/M2/s1 ;
 wire \V3/V3/V3/A2/M3/c1 ;
 wire \V3/V3/V3/A2/M3/c2 ;
 wire \V3/V3/V3/A2/M3/s1 ;
 wire \V3/V3/V3/A2/M4/c1 ;
 wire \V3/V3/V3/A2/M4/c2 ;
 wire \V3/V3/V3/A2/M4/s1 ;
 wire \V3/V3/V3/A3/c1 ;
 wire \V3/V3/V3/A3/c2 ;
 wire \V3/V3/V3/A3/c3 ;
 wire \V3/V3/V3/A3/M1/c1 ;
 wire \V3/V3/V3/A3/M1/c2 ;
 wire \V3/V3/V3/A3/M1/s1 ;
 wire \V3/V3/V3/A3/M2/c1 ;
 wire \V3/V3/V3/A3/M2/c2 ;
 wire \V3/V3/V3/A3/M2/s1 ;
 wire \V3/V3/V3/A3/M3/c1 ;
 wire \V3/V3/V3/A3/M3/c2 ;
 wire \V3/V3/V3/A3/M3/s1 ;
 wire \V3/V3/V3/A3/M4/c1 ;
 wire \V3/V3/V3/A3/M4/c2 ;
 wire \V3/V3/V3/A3/M4/s1 ;
 wire \V3/V3/V3/V1/w1 ;
 wire \V3/V3/V3/V1/w2 ;
 wire \V3/V3/V3/V1/w3 ;
 wire \V3/V3/V3/V1/w4 ;
 wire \V3/V3/V3/V2/w1 ;
 wire \V3/V3/V3/V2/w2 ;
 wire \V3/V3/V3/V2/w3 ;
 wire \V3/V3/V3/V2/w4 ;
 wire \V3/V3/V3/V3/w1 ;
 wire \V3/V3/V3/V3/w2 ;
 wire \V3/V3/V3/V3/w3 ;
 wire \V3/V3/V3/V3/w4 ;
 wire \V3/V3/V3/V4/w1 ;
 wire \V3/V3/V3/V4/w2 ;
 wire \V3/V3/V3/V4/w3 ;
 wire \V3/V3/V3/V4/w4 ;
 wire \V3/V3/V4/c1 ;
 wire \V3/V3/V4/c2 ;
 wire \V3/V3/V4/c3 ;
 wire \V3/V3/V4/overflow ;
 wire \V3/V3/V4/A1/c1 ;
 wire \V3/V3/V4/A1/c2 ;
 wire \V3/V3/V4/A1/c3 ;
 wire \V3/V3/V4/A1/M1/c1 ;
 wire \V3/V3/V4/A1/M1/c2 ;
 wire \V3/V3/V4/A1/M1/s1 ;
 wire \V3/V3/V4/A1/M2/c1 ;
 wire \V3/V3/V4/A1/M2/c2 ;
 wire \V3/V3/V4/A1/M2/s1 ;
 wire \V3/V3/V4/A1/M3/c1 ;
 wire \V3/V3/V4/A1/M3/c2 ;
 wire \V3/V3/V4/A1/M3/s1 ;
 wire \V3/V3/V4/A1/M4/c1 ;
 wire \V3/V3/V4/A1/M4/c2 ;
 wire \V3/V3/V4/A1/M4/s1 ;
 wire \V3/V3/V4/A2/c1 ;
 wire \V3/V3/V4/A2/c2 ;
 wire \V3/V3/V4/A2/c3 ;
 wire \V3/V3/V4/A2/M1/c1 ;
 wire \V3/V3/V4/A2/M1/c2 ;
 wire \V3/V3/V4/A2/M1/s1 ;
 wire \V3/V3/V4/A2/M2/c1 ;
 wire \V3/V3/V4/A2/M2/c2 ;
 wire \V3/V3/V4/A2/M2/s1 ;
 wire \V3/V3/V4/A2/M3/c1 ;
 wire \V3/V3/V4/A2/M3/c2 ;
 wire \V3/V3/V4/A2/M3/s1 ;
 wire \V3/V3/V4/A2/M4/c1 ;
 wire \V3/V3/V4/A2/M4/c2 ;
 wire \V3/V3/V4/A2/M4/s1 ;
 wire \V3/V3/V4/A3/c1 ;
 wire \V3/V3/V4/A3/c2 ;
 wire \V3/V3/V4/A3/c3 ;
 wire \V3/V3/V4/A3/M1/c1 ;
 wire \V3/V3/V4/A3/M1/c2 ;
 wire \V3/V3/V4/A3/M1/s1 ;
 wire \V3/V3/V4/A3/M2/c1 ;
 wire \V3/V3/V4/A3/M2/c2 ;
 wire \V3/V3/V4/A3/M2/s1 ;
 wire \V3/V3/V4/A3/M3/c1 ;
 wire \V3/V3/V4/A3/M3/c2 ;
 wire \V3/V3/V4/A3/M3/s1 ;
 wire \V3/V3/V4/A3/M4/c1 ;
 wire \V3/V3/V4/A3/M4/c2 ;
 wire \V3/V3/V4/A3/M4/s1 ;
 wire \V3/V3/V4/V1/w1 ;
 wire \V3/V3/V4/V1/w2 ;
 wire \V3/V3/V4/V1/w3 ;
 wire \V3/V3/V4/V1/w4 ;
 wire \V3/V3/V4/V2/w1 ;
 wire \V3/V3/V4/V2/w2 ;
 wire \V3/V3/V4/V2/w3 ;
 wire \V3/V3/V4/V2/w4 ;
 wire \V3/V3/V4/V3/w1 ;
 wire \V3/V3/V4/V3/w2 ;
 wire \V3/V3/V4/V3/w3 ;
 wire \V3/V3/V4/V3/w4 ;
 wire \V3/V3/V4/V4/w1 ;
 wire \V3/V3/V4/V4/w2 ;
 wire \V3/V3/V4/V4/w3 ;
 wire \V3/V3/V4/V4/w4 ;
 wire \V3/V4/c1 ;
 wire \V3/V4/c2 ;
 wire \V3/V4/c3 ;
 wire \V3/V4/overflow ;
 wire \V3/V4/A1/c1 ;
 wire \V3/V4/A1/A1/c1 ;
 wire \V3/V4/A1/A1/c2 ;
 wire \V3/V4/A1/A1/c3 ;
 wire \V3/V4/A1/A1/M1/c1 ;
 wire \V3/V4/A1/A1/M1/c2 ;
 wire \V3/V4/A1/A1/M1/s1 ;
 wire \V3/V4/A1/A1/M2/c1 ;
 wire \V3/V4/A1/A1/M2/c2 ;
 wire \V3/V4/A1/A1/M2/s1 ;
 wire \V3/V4/A1/A1/M3/c1 ;
 wire \V3/V4/A1/A1/M3/c2 ;
 wire \V3/V4/A1/A1/M3/s1 ;
 wire \V3/V4/A1/A1/M4/c1 ;
 wire \V3/V4/A1/A1/M4/c2 ;
 wire \V3/V4/A1/A1/M4/s1 ;
 wire \V3/V4/A1/A2/c1 ;
 wire \V3/V4/A1/A2/c2 ;
 wire \V3/V4/A1/A2/c3 ;
 wire \V3/V4/A1/A2/M1/c1 ;
 wire \V3/V4/A1/A2/M1/c2 ;
 wire \V3/V4/A1/A2/M1/s1 ;
 wire \V3/V4/A1/A2/M2/c1 ;
 wire \V3/V4/A1/A2/M2/c2 ;
 wire \V3/V4/A1/A2/M2/s1 ;
 wire \V3/V4/A1/A2/M3/c1 ;
 wire \V3/V4/A1/A2/M3/c2 ;
 wire \V3/V4/A1/A2/M3/s1 ;
 wire \V3/V4/A1/A2/M4/c1 ;
 wire \V3/V4/A1/A2/M4/c2 ;
 wire \V3/V4/A1/A2/M4/s1 ;
 wire \V3/V4/A2/c1 ;
 wire \V3/V4/A2/A1/c1 ;
 wire \V3/V4/A2/A1/c2 ;
 wire \V3/V4/A2/A1/c3 ;
 wire \V3/V4/A2/A1/M1/c1 ;
 wire \V3/V4/A2/A1/M1/c2 ;
 wire \V3/V4/A2/A1/M1/s1 ;
 wire \V3/V4/A2/A1/M2/c1 ;
 wire \V3/V4/A2/A1/M2/c2 ;
 wire \V3/V4/A2/A1/M2/s1 ;
 wire \V3/V4/A2/A1/M3/c1 ;
 wire \V3/V4/A2/A1/M3/c2 ;
 wire \V3/V4/A2/A1/M3/s1 ;
 wire \V3/V4/A2/A1/M4/c1 ;
 wire \V3/V4/A2/A1/M4/c2 ;
 wire \V3/V4/A2/A1/M4/s1 ;
 wire \V3/V4/A2/A2/c1 ;
 wire \V3/V4/A2/A2/c2 ;
 wire \V3/V4/A2/A2/c3 ;
 wire \V3/V4/A2/A2/M1/c1 ;
 wire \V3/V4/A2/A2/M1/c2 ;
 wire \V3/V4/A2/A2/M1/s1 ;
 wire \V3/V4/A2/A2/M2/c1 ;
 wire \V3/V4/A2/A2/M2/c2 ;
 wire \V3/V4/A2/A2/M2/s1 ;
 wire \V3/V4/A2/A2/M3/c1 ;
 wire \V3/V4/A2/A2/M3/c2 ;
 wire \V3/V4/A2/A2/M3/s1 ;
 wire \V3/V4/A2/A2/M4/c1 ;
 wire \V3/V4/A2/A2/M4/c2 ;
 wire \V3/V4/A2/A2/M4/s1 ;
 wire \V3/V4/A3/c1 ;
 wire \V3/V4/A3/A1/c1 ;
 wire \V3/V4/A3/A1/c2 ;
 wire \V3/V4/A3/A1/c3 ;
 wire \V3/V4/A3/A1/M1/c1 ;
 wire \V3/V4/A3/A1/M1/c2 ;
 wire \V3/V4/A3/A1/M1/s1 ;
 wire \V3/V4/A3/A1/M2/c1 ;
 wire \V3/V4/A3/A1/M2/c2 ;
 wire \V3/V4/A3/A1/M2/s1 ;
 wire \V3/V4/A3/A1/M3/c1 ;
 wire \V3/V4/A3/A1/M3/c2 ;
 wire \V3/V4/A3/A1/M3/s1 ;
 wire \V3/V4/A3/A1/M4/c1 ;
 wire \V3/V4/A3/A1/M4/c2 ;
 wire \V3/V4/A3/A1/M4/s1 ;
 wire \V3/V4/A3/A2/c1 ;
 wire \V3/V4/A3/A2/c2 ;
 wire \V3/V4/A3/A2/c3 ;
 wire \V3/V4/A3/A2/M1/c1 ;
 wire \V3/V4/A3/A2/M1/c2 ;
 wire \V3/V4/A3/A2/M1/s1 ;
 wire \V3/V4/A3/A2/M2/c1 ;
 wire \V3/V4/A3/A2/M2/c2 ;
 wire \V3/V4/A3/A2/M2/s1 ;
 wire \V3/V4/A3/A2/M3/c1 ;
 wire \V3/V4/A3/A2/M3/c2 ;
 wire \V3/V4/A3/A2/M3/s1 ;
 wire \V3/V4/A3/A2/M4/c1 ;
 wire \V3/V4/A3/A2/M4/c2 ;
 wire \V3/V4/A3/A2/M4/s1 ;
 wire \V3/V4/V1/c1 ;
 wire \V3/V4/V1/c2 ;
 wire \V3/V4/V1/c3 ;
 wire \V3/V4/V1/overflow ;
 wire \V3/V4/V1/A1/c1 ;
 wire \V3/V4/V1/A1/c2 ;
 wire \V3/V4/V1/A1/c3 ;
 wire \V3/V4/V1/A1/M1/c1 ;
 wire \V3/V4/V1/A1/M1/c2 ;
 wire \V3/V4/V1/A1/M1/s1 ;
 wire \V3/V4/V1/A1/M2/c1 ;
 wire \V3/V4/V1/A1/M2/c2 ;
 wire \V3/V4/V1/A1/M2/s1 ;
 wire \V3/V4/V1/A1/M3/c1 ;
 wire \V3/V4/V1/A1/M3/c2 ;
 wire \V3/V4/V1/A1/M3/s1 ;
 wire \V3/V4/V1/A1/M4/c1 ;
 wire \V3/V4/V1/A1/M4/c2 ;
 wire \V3/V4/V1/A1/M4/s1 ;
 wire \V3/V4/V1/A2/c1 ;
 wire \V3/V4/V1/A2/c2 ;
 wire \V3/V4/V1/A2/c3 ;
 wire \V3/V4/V1/A2/M1/c1 ;
 wire \V3/V4/V1/A2/M1/c2 ;
 wire \V3/V4/V1/A2/M1/s1 ;
 wire \V3/V4/V1/A2/M2/c1 ;
 wire \V3/V4/V1/A2/M2/c2 ;
 wire \V3/V4/V1/A2/M2/s1 ;
 wire \V3/V4/V1/A2/M3/c1 ;
 wire \V3/V4/V1/A2/M3/c2 ;
 wire \V3/V4/V1/A2/M3/s1 ;
 wire \V3/V4/V1/A2/M4/c1 ;
 wire \V3/V4/V1/A2/M4/c2 ;
 wire \V3/V4/V1/A2/M4/s1 ;
 wire \V3/V4/V1/A3/c1 ;
 wire \V3/V4/V1/A3/c2 ;
 wire \V3/V4/V1/A3/c3 ;
 wire \V3/V4/V1/A3/M1/c1 ;
 wire \V3/V4/V1/A3/M1/c2 ;
 wire \V3/V4/V1/A3/M1/s1 ;
 wire \V3/V4/V1/A3/M2/c1 ;
 wire \V3/V4/V1/A3/M2/c2 ;
 wire \V3/V4/V1/A3/M2/s1 ;
 wire \V3/V4/V1/A3/M3/c1 ;
 wire \V3/V4/V1/A3/M3/c2 ;
 wire \V3/V4/V1/A3/M3/s1 ;
 wire \V3/V4/V1/A3/M4/c1 ;
 wire \V3/V4/V1/A3/M4/c2 ;
 wire \V3/V4/V1/A3/M4/s1 ;
 wire \V3/V4/V1/V1/w1 ;
 wire \V3/V4/V1/V1/w2 ;
 wire \V3/V4/V1/V1/w3 ;
 wire \V3/V4/V1/V1/w4 ;
 wire \V3/V4/V1/V2/w1 ;
 wire \V3/V4/V1/V2/w2 ;
 wire \V3/V4/V1/V2/w3 ;
 wire \V3/V4/V1/V2/w4 ;
 wire \V3/V4/V1/V3/w1 ;
 wire \V3/V4/V1/V3/w2 ;
 wire \V3/V4/V1/V3/w3 ;
 wire \V3/V4/V1/V3/w4 ;
 wire \V3/V4/V1/V4/w1 ;
 wire \V3/V4/V1/V4/w2 ;
 wire \V3/V4/V1/V4/w3 ;
 wire \V3/V4/V1/V4/w4 ;
 wire \V3/V4/V2/c1 ;
 wire \V3/V4/V2/c2 ;
 wire \V3/V4/V2/c3 ;
 wire \V3/V4/V2/overflow ;
 wire \V3/V4/V2/A1/c1 ;
 wire \V3/V4/V2/A1/c2 ;
 wire \V3/V4/V2/A1/c3 ;
 wire \V3/V4/V2/A1/M1/c1 ;
 wire \V3/V4/V2/A1/M1/c2 ;
 wire \V3/V4/V2/A1/M1/s1 ;
 wire \V3/V4/V2/A1/M2/c1 ;
 wire \V3/V4/V2/A1/M2/c2 ;
 wire \V3/V4/V2/A1/M2/s1 ;
 wire \V3/V4/V2/A1/M3/c1 ;
 wire \V3/V4/V2/A1/M3/c2 ;
 wire \V3/V4/V2/A1/M3/s1 ;
 wire \V3/V4/V2/A1/M4/c1 ;
 wire \V3/V4/V2/A1/M4/c2 ;
 wire \V3/V4/V2/A1/M4/s1 ;
 wire \V3/V4/V2/A2/c1 ;
 wire \V3/V4/V2/A2/c2 ;
 wire \V3/V4/V2/A2/c3 ;
 wire \V3/V4/V2/A2/M1/c1 ;
 wire \V3/V4/V2/A2/M1/c2 ;
 wire \V3/V4/V2/A2/M1/s1 ;
 wire \V3/V4/V2/A2/M2/c1 ;
 wire \V3/V4/V2/A2/M2/c2 ;
 wire \V3/V4/V2/A2/M2/s1 ;
 wire \V3/V4/V2/A2/M3/c1 ;
 wire \V3/V4/V2/A2/M3/c2 ;
 wire \V3/V4/V2/A2/M3/s1 ;
 wire \V3/V4/V2/A2/M4/c1 ;
 wire \V3/V4/V2/A2/M4/c2 ;
 wire \V3/V4/V2/A2/M4/s1 ;
 wire \V3/V4/V2/A3/c1 ;
 wire \V3/V4/V2/A3/c2 ;
 wire \V3/V4/V2/A3/c3 ;
 wire \V3/V4/V2/A3/M1/c1 ;
 wire \V3/V4/V2/A3/M1/c2 ;
 wire \V3/V4/V2/A3/M1/s1 ;
 wire \V3/V4/V2/A3/M2/c1 ;
 wire \V3/V4/V2/A3/M2/c2 ;
 wire \V3/V4/V2/A3/M2/s1 ;
 wire \V3/V4/V2/A3/M3/c1 ;
 wire \V3/V4/V2/A3/M3/c2 ;
 wire \V3/V4/V2/A3/M3/s1 ;
 wire \V3/V4/V2/A3/M4/c1 ;
 wire \V3/V4/V2/A3/M4/c2 ;
 wire \V3/V4/V2/A3/M4/s1 ;
 wire \V3/V4/V2/V1/w1 ;
 wire \V3/V4/V2/V1/w2 ;
 wire \V3/V4/V2/V1/w3 ;
 wire \V3/V4/V2/V1/w4 ;
 wire \V3/V4/V2/V2/w1 ;
 wire \V3/V4/V2/V2/w2 ;
 wire \V3/V4/V2/V2/w3 ;
 wire \V3/V4/V2/V2/w4 ;
 wire \V3/V4/V2/V3/w1 ;
 wire \V3/V4/V2/V3/w2 ;
 wire \V3/V4/V2/V3/w3 ;
 wire \V3/V4/V2/V3/w4 ;
 wire \V3/V4/V2/V4/w1 ;
 wire \V3/V4/V2/V4/w2 ;
 wire \V3/V4/V2/V4/w3 ;
 wire \V3/V4/V2/V4/w4 ;
 wire \V3/V4/V3/c1 ;
 wire \V3/V4/V3/c2 ;
 wire \V3/V4/V3/c3 ;
 wire \V3/V4/V3/overflow ;
 wire \V3/V4/V3/A1/c1 ;
 wire \V3/V4/V3/A1/c2 ;
 wire \V3/V4/V3/A1/c3 ;
 wire \V3/V4/V3/A1/M1/c1 ;
 wire \V3/V4/V3/A1/M1/c2 ;
 wire \V3/V4/V3/A1/M1/s1 ;
 wire \V3/V4/V3/A1/M2/c1 ;
 wire \V3/V4/V3/A1/M2/c2 ;
 wire \V3/V4/V3/A1/M2/s1 ;
 wire \V3/V4/V3/A1/M3/c1 ;
 wire \V3/V4/V3/A1/M3/c2 ;
 wire \V3/V4/V3/A1/M3/s1 ;
 wire \V3/V4/V3/A1/M4/c1 ;
 wire \V3/V4/V3/A1/M4/c2 ;
 wire \V3/V4/V3/A1/M4/s1 ;
 wire \V3/V4/V3/A2/c1 ;
 wire \V3/V4/V3/A2/c2 ;
 wire \V3/V4/V3/A2/c3 ;
 wire \V3/V4/V3/A2/M1/c1 ;
 wire \V3/V4/V3/A2/M1/c2 ;
 wire \V3/V4/V3/A2/M1/s1 ;
 wire \V3/V4/V3/A2/M2/c1 ;
 wire \V3/V4/V3/A2/M2/c2 ;
 wire \V3/V4/V3/A2/M2/s1 ;
 wire \V3/V4/V3/A2/M3/c1 ;
 wire \V3/V4/V3/A2/M3/c2 ;
 wire \V3/V4/V3/A2/M3/s1 ;
 wire \V3/V4/V3/A2/M4/c1 ;
 wire \V3/V4/V3/A2/M4/c2 ;
 wire \V3/V4/V3/A2/M4/s1 ;
 wire \V3/V4/V3/A3/c1 ;
 wire \V3/V4/V3/A3/c2 ;
 wire \V3/V4/V3/A3/c3 ;
 wire \V3/V4/V3/A3/M1/c1 ;
 wire \V3/V4/V3/A3/M1/c2 ;
 wire \V3/V4/V3/A3/M1/s1 ;
 wire \V3/V4/V3/A3/M2/c1 ;
 wire \V3/V4/V3/A3/M2/c2 ;
 wire \V3/V4/V3/A3/M2/s1 ;
 wire \V3/V4/V3/A3/M3/c1 ;
 wire \V3/V4/V3/A3/M3/c2 ;
 wire \V3/V4/V3/A3/M3/s1 ;
 wire \V3/V4/V3/A3/M4/c1 ;
 wire \V3/V4/V3/A3/M4/c2 ;
 wire \V3/V4/V3/A3/M4/s1 ;
 wire \V3/V4/V3/V1/w1 ;
 wire \V3/V4/V3/V1/w2 ;
 wire \V3/V4/V3/V1/w3 ;
 wire \V3/V4/V3/V1/w4 ;
 wire \V3/V4/V3/V2/w1 ;
 wire \V3/V4/V3/V2/w2 ;
 wire \V3/V4/V3/V2/w3 ;
 wire \V3/V4/V3/V2/w4 ;
 wire \V3/V4/V3/V3/w1 ;
 wire \V3/V4/V3/V3/w2 ;
 wire \V3/V4/V3/V3/w3 ;
 wire \V3/V4/V3/V3/w4 ;
 wire \V3/V4/V3/V4/w1 ;
 wire \V3/V4/V3/V4/w2 ;
 wire \V3/V4/V3/V4/w3 ;
 wire \V3/V4/V3/V4/w4 ;
 wire \V3/V4/V4/c1 ;
 wire \V3/V4/V4/c2 ;
 wire \V3/V4/V4/c3 ;
 wire \V3/V4/V4/overflow ;
 wire \V3/V4/V4/A1/c1 ;
 wire \V3/V4/V4/A1/c2 ;
 wire \V3/V4/V4/A1/c3 ;
 wire \V3/V4/V4/A1/M1/c1 ;
 wire \V3/V4/V4/A1/M1/c2 ;
 wire \V3/V4/V4/A1/M1/s1 ;
 wire \V3/V4/V4/A1/M2/c1 ;
 wire \V3/V4/V4/A1/M2/c2 ;
 wire \V3/V4/V4/A1/M2/s1 ;
 wire \V3/V4/V4/A1/M3/c1 ;
 wire \V3/V4/V4/A1/M3/c2 ;
 wire \V3/V4/V4/A1/M3/s1 ;
 wire \V3/V4/V4/A1/M4/c1 ;
 wire \V3/V4/V4/A1/M4/c2 ;
 wire \V3/V4/V4/A1/M4/s1 ;
 wire \V3/V4/V4/A2/c1 ;
 wire \V3/V4/V4/A2/c2 ;
 wire \V3/V4/V4/A2/c3 ;
 wire \V3/V4/V4/A2/M1/c1 ;
 wire \V3/V4/V4/A2/M1/c2 ;
 wire \V3/V4/V4/A2/M1/s1 ;
 wire \V3/V4/V4/A2/M2/c1 ;
 wire \V3/V4/V4/A2/M2/c2 ;
 wire \V3/V4/V4/A2/M2/s1 ;
 wire \V3/V4/V4/A2/M3/c1 ;
 wire \V3/V4/V4/A2/M3/c2 ;
 wire \V3/V4/V4/A2/M3/s1 ;
 wire \V3/V4/V4/A2/M4/c1 ;
 wire \V3/V4/V4/A2/M4/c2 ;
 wire \V3/V4/V4/A2/M4/s1 ;
 wire \V3/V4/V4/A3/c1 ;
 wire \V3/V4/V4/A3/c2 ;
 wire \V3/V4/V4/A3/c3 ;
 wire \V3/V4/V4/A3/M1/c1 ;
 wire \V3/V4/V4/A3/M1/c2 ;
 wire \V3/V4/V4/A3/M1/s1 ;
 wire \V3/V4/V4/A3/M2/c1 ;
 wire \V3/V4/V4/A3/M2/c2 ;
 wire \V3/V4/V4/A3/M2/s1 ;
 wire \V3/V4/V4/A3/M3/c1 ;
 wire \V3/V4/V4/A3/M3/c2 ;
 wire \V3/V4/V4/A3/M3/s1 ;
 wire \V3/V4/V4/A3/M4/c1 ;
 wire \V3/V4/V4/A3/M4/c2 ;
 wire \V3/V4/V4/A3/M4/s1 ;
 wire \V3/V4/V4/V1/w1 ;
 wire \V3/V4/V4/V1/w2 ;
 wire \V3/V4/V4/V1/w3 ;
 wire \V3/V4/V4/V1/w4 ;
 wire \V3/V4/V4/V2/w1 ;
 wire \V3/V4/V4/V2/w2 ;
 wire \V3/V4/V4/V2/w3 ;
 wire \V3/V4/V4/V2/w4 ;
 wire \V3/V4/V4/V3/w1 ;
 wire \V3/V4/V4/V3/w2 ;
 wire \V3/V4/V4/V3/w3 ;
 wire \V3/V4/V4/V3/w4 ;
 wire \V3/V4/V4/V4/w1 ;
 wire \V3/V4/V4/V4/w2 ;
 wire \V3/V4/V4/V4/w3 ;
 wire \V3/V4/V4/V4/w4 ;
 wire \V4/c1 ;
 wire \V4/c2 ;
 wire \V4/c3 ;
 wire \V4/overflow ;
 wire \V4/A1/c1 ;
 wire \V4/A1/A1/c1 ;
 wire \V4/A1/A1/A1/c1 ;
 wire \V4/A1/A1/A1/c2 ;
 wire \V4/A1/A1/A1/c3 ;
 wire \V4/A1/A1/A1/M1/c1 ;
 wire \V4/A1/A1/A1/M1/c2 ;
 wire \V4/A1/A1/A1/M1/s1 ;
 wire \V4/A1/A1/A1/M2/c1 ;
 wire \V4/A1/A1/A1/M2/c2 ;
 wire \V4/A1/A1/A1/M2/s1 ;
 wire \V4/A1/A1/A1/M3/c1 ;
 wire \V4/A1/A1/A1/M3/c2 ;
 wire \V4/A1/A1/A1/M3/s1 ;
 wire \V4/A1/A1/A1/M4/c1 ;
 wire \V4/A1/A1/A1/M4/c2 ;
 wire \V4/A1/A1/A1/M4/s1 ;
 wire \V4/A1/A1/A2/c1 ;
 wire \V4/A1/A1/A2/c2 ;
 wire \V4/A1/A1/A2/c3 ;
 wire \V4/A1/A1/A2/M1/c1 ;
 wire \V4/A1/A1/A2/M1/c2 ;
 wire \V4/A1/A1/A2/M1/s1 ;
 wire \V4/A1/A1/A2/M2/c1 ;
 wire \V4/A1/A1/A2/M2/c2 ;
 wire \V4/A1/A1/A2/M2/s1 ;
 wire \V4/A1/A1/A2/M3/c1 ;
 wire \V4/A1/A1/A2/M3/c2 ;
 wire \V4/A1/A1/A2/M3/s1 ;
 wire \V4/A1/A1/A2/M4/c1 ;
 wire \V4/A1/A1/A2/M4/c2 ;
 wire \V4/A1/A1/A2/M4/s1 ;
 wire \V4/A1/A2/c1 ;
 wire \V4/A1/A2/A1/c1 ;
 wire \V4/A1/A2/A1/c2 ;
 wire \V4/A1/A2/A1/c3 ;
 wire \V4/A1/A2/A1/M1/c1 ;
 wire \V4/A1/A2/A1/M1/c2 ;
 wire \V4/A1/A2/A1/M1/s1 ;
 wire \V4/A1/A2/A1/M2/c1 ;
 wire \V4/A1/A2/A1/M2/c2 ;
 wire \V4/A1/A2/A1/M2/s1 ;
 wire \V4/A1/A2/A1/M3/c1 ;
 wire \V4/A1/A2/A1/M3/c2 ;
 wire \V4/A1/A2/A1/M3/s1 ;
 wire \V4/A1/A2/A1/M4/c1 ;
 wire \V4/A1/A2/A1/M4/c2 ;
 wire \V4/A1/A2/A1/M4/s1 ;
 wire \V4/A1/A2/A2/c1 ;
 wire \V4/A1/A2/A2/c2 ;
 wire \V4/A1/A2/A2/c3 ;
 wire \V4/A1/A2/A2/M1/c1 ;
 wire \V4/A1/A2/A2/M1/c2 ;
 wire \V4/A1/A2/A2/M1/s1 ;
 wire \V4/A1/A2/A2/M2/c1 ;
 wire \V4/A1/A2/A2/M2/c2 ;
 wire \V4/A1/A2/A2/M2/s1 ;
 wire \V4/A1/A2/A2/M3/c1 ;
 wire \V4/A1/A2/A2/M3/c2 ;
 wire \V4/A1/A2/A2/M3/s1 ;
 wire \V4/A1/A2/A2/M4/c1 ;
 wire \V4/A1/A2/A2/M4/c2 ;
 wire \V4/A1/A2/A2/M4/s1 ;
 wire \V4/A2/c1 ;
 wire \V4/A2/A1/c1 ;
 wire \V4/A2/A1/A1/c1 ;
 wire \V4/A2/A1/A1/c2 ;
 wire \V4/A2/A1/A1/c3 ;
 wire \V4/A2/A1/A1/M1/c1 ;
 wire \V4/A2/A1/A1/M1/c2 ;
 wire \V4/A2/A1/A1/M1/s1 ;
 wire \V4/A2/A1/A1/M2/c1 ;
 wire \V4/A2/A1/A1/M2/c2 ;
 wire \V4/A2/A1/A1/M2/s1 ;
 wire \V4/A2/A1/A1/M3/c1 ;
 wire \V4/A2/A1/A1/M3/c2 ;
 wire \V4/A2/A1/A1/M3/s1 ;
 wire \V4/A2/A1/A1/M4/c1 ;
 wire \V4/A2/A1/A1/M4/c2 ;
 wire \V4/A2/A1/A1/M4/s1 ;
 wire \V4/A2/A1/A2/c1 ;
 wire \V4/A2/A1/A2/c2 ;
 wire \V4/A2/A1/A2/c3 ;
 wire \V4/A2/A1/A2/M1/c1 ;
 wire \V4/A2/A1/A2/M1/c2 ;
 wire \V4/A2/A1/A2/M1/s1 ;
 wire \V4/A2/A1/A2/M2/c1 ;
 wire \V4/A2/A1/A2/M2/c2 ;
 wire \V4/A2/A1/A2/M2/s1 ;
 wire \V4/A2/A1/A2/M3/c1 ;
 wire \V4/A2/A1/A2/M3/c2 ;
 wire \V4/A2/A1/A2/M3/s1 ;
 wire \V4/A2/A1/A2/M4/c1 ;
 wire \V4/A2/A1/A2/M4/c2 ;
 wire \V4/A2/A1/A2/M4/s1 ;
 wire \V4/A2/A2/c1 ;
 wire \V4/A2/A2/A1/c1 ;
 wire \V4/A2/A2/A1/c2 ;
 wire \V4/A2/A2/A1/c3 ;
 wire \V4/A2/A2/A1/M1/c1 ;
 wire \V4/A2/A2/A1/M1/c2 ;
 wire \V4/A2/A2/A1/M1/s1 ;
 wire \V4/A2/A2/A1/M2/c1 ;
 wire \V4/A2/A2/A1/M2/c2 ;
 wire \V4/A2/A2/A1/M2/s1 ;
 wire \V4/A2/A2/A1/M3/c1 ;
 wire \V4/A2/A2/A1/M3/c2 ;
 wire \V4/A2/A2/A1/M3/s1 ;
 wire \V4/A2/A2/A1/M4/c1 ;
 wire \V4/A2/A2/A1/M4/c2 ;
 wire \V4/A2/A2/A1/M4/s1 ;
 wire \V4/A2/A2/A2/c1 ;
 wire \V4/A2/A2/A2/c2 ;
 wire \V4/A2/A2/A2/c3 ;
 wire \V4/A2/A2/A2/M1/c1 ;
 wire \V4/A2/A2/A2/M1/c2 ;
 wire \V4/A2/A2/A2/M1/s1 ;
 wire \V4/A2/A2/A2/M2/c1 ;
 wire \V4/A2/A2/A2/M2/c2 ;
 wire \V4/A2/A2/A2/M2/s1 ;
 wire \V4/A2/A2/A2/M3/c1 ;
 wire \V4/A2/A2/A2/M3/c2 ;
 wire \V4/A2/A2/A2/M3/s1 ;
 wire \V4/A2/A2/A2/M4/c1 ;
 wire \V4/A2/A2/A2/M4/c2 ;
 wire \V4/A2/A2/A2/M4/s1 ;
 wire \V4/A3/c1 ;
 wire \V4/A3/A1/c1 ;
 wire \V4/A3/A1/A1/c1 ;
 wire \V4/A3/A1/A1/c2 ;
 wire \V4/A3/A1/A1/c3 ;
 wire \V4/A3/A1/A1/M1/c1 ;
 wire \V4/A3/A1/A1/M1/c2 ;
 wire \V4/A3/A1/A1/M1/s1 ;
 wire \V4/A3/A1/A1/M2/c1 ;
 wire \V4/A3/A1/A1/M2/c2 ;
 wire \V4/A3/A1/A1/M2/s1 ;
 wire \V4/A3/A1/A1/M3/c1 ;
 wire \V4/A3/A1/A1/M3/c2 ;
 wire \V4/A3/A1/A1/M3/s1 ;
 wire \V4/A3/A1/A1/M4/c1 ;
 wire \V4/A3/A1/A1/M4/c2 ;
 wire \V4/A3/A1/A1/M4/s1 ;
 wire \V4/A3/A1/A2/c1 ;
 wire \V4/A3/A1/A2/c2 ;
 wire \V4/A3/A1/A2/c3 ;
 wire \V4/A3/A1/A2/M1/c1 ;
 wire \V4/A3/A1/A2/M1/c2 ;
 wire \V4/A3/A1/A2/M1/s1 ;
 wire \V4/A3/A1/A2/M2/c1 ;
 wire \V4/A3/A1/A2/M2/c2 ;
 wire \V4/A3/A1/A2/M2/s1 ;
 wire \V4/A3/A1/A2/M3/c1 ;
 wire \V4/A3/A1/A2/M3/c2 ;
 wire \V4/A3/A1/A2/M3/s1 ;
 wire \V4/A3/A1/A2/M4/c1 ;
 wire \V4/A3/A1/A2/M4/c2 ;
 wire \V4/A3/A1/A2/M4/s1 ;
 wire \V4/A3/A2/c1 ;
 wire \V4/A3/A2/A1/c1 ;
 wire \V4/A3/A2/A1/c2 ;
 wire \V4/A3/A2/A1/c3 ;
 wire \V4/A3/A2/A1/M1/c1 ;
 wire \V4/A3/A2/A1/M1/c2 ;
 wire \V4/A3/A2/A1/M1/s1 ;
 wire \V4/A3/A2/A1/M2/c1 ;
 wire \V4/A3/A2/A1/M2/c2 ;
 wire \V4/A3/A2/A1/M2/s1 ;
 wire \V4/A3/A2/A1/M3/c1 ;
 wire \V4/A3/A2/A1/M3/c2 ;
 wire \V4/A3/A2/A1/M3/s1 ;
 wire \V4/A3/A2/A1/M4/c1 ;
 wire \V4/A3/A2/A1/M4/c2 ;
 wire \V4/A3/A2/A1/M4/s1 ;
 wire \V4/A3/A2/A2/c1 ;
 wire \V4/A3/A2/A2/c2 ;
 wire \V4/A3/A2/A2/c3 ;
 wire \V4/A3/A2/A2/M1/c1 ;
 wire \V4/A3/A2/A2/M1/c2 ;
 wire \V4/A3/A2/A2/M1/s1 ;
 wire \V4/A3/A2/A2/M2/c1 ;
 wire \V4/A3/A2/A2/M2/c2 ;
 wire \V4/A3/A2/A2/M2/s1 ;
 wire \V4/A3/A2/A2/M3/c1 ;
 wire \V4/A3/A2/A2/M3/c2 ;
 wire \V4/A3/A2/A2/M3/s1 ;
 wire \V4/A3/A2/A2/M4/c1 ;
 wire \V4/A3/A2/A2/M4/c2 ;
 wire \V4/A3/A2/A2/M4/s1 ;
 wire \V4/V1/c1 ;
 wire \V4/V1/c2 ;
 wire \V4/V1/c3 ;
 wire \V4/V1/overflow ;
 wire \V4/V1/A1/c1 ;
 wire \V4/V1/A1/A1/c1 ;
 wire \V4/V1/A1/A1/c2 ;
 wire \V4/V1/A1/A1/c3 ;
 wire \V4/V1/A1/A1/M1/c1 ;
 wire \V4/V1/A1/A1/M1/c2 ;
 wire \V4/V1/A1/A1/M1/s1 ;
 wire \V4/V1/A1/A1/M2/c1 ;
 wire \V4/V1/A1/A1/M2/c2 ;
 wire \V4/V1/A1/A1/M2/s1 ;
 wire \V4/V1/A1/A1/M3/c1 ;
 wire \V4/V1/A1/A1/M3/c2 ;
 wire \V4/V1/A1/A1/M3/s1 ;
 wire \V4/V1/A1/A1/M4/c1 ;
 wire \V4/V1/A1/A1/M4/c2 ;
 wire \V4/V1/A1/A1/M4/s1 ;
 wire \V4/V1/A1/A2/c1 ;
 wire \V4/V1/A1/A2/c2 ;
 wire \V4/V1/A1/A2/c3 ;
 wire \V4/V1/A1/A2/M1/c1 ;
 wire \V4/V1/A1/A2/M1/c2 ;
 wire \V4/V1/A1/A2/M1/s1 ;
 wire \V4/V1/A1/A2/M2/c1 ;
 wire \V4/V1/A1/A2/M2/c2 ;
 wire \V4/V1/A1/A2/M2/s1 ;
 wire \V4/V1/A1/A2/M3/c1 ;
 wire \V4/V1/A1/A2/M3/c2 ;
 wire \V4/V1/A1/A2/M3/s1 ;
 wire \V4/V1/A1/A2/M4/c1 ;
 wire \V4/V1/A1/A2/M4/c2 ;
 wire \V4/V1/A1/A2/M4/s1 ;
 wire \V4/V1/A2/c1 ;
 wire \V4/V1/A2/A1/c1 ;
 wire \V4/V1/A2/A1/c2 ;
 wire \V4/V1/A2/A1/c3 ;
 wire \V4/V1/A2/A1/M1/c1 ;
 wire \V4/V1/A2/A1/M1/c2 ;
 wire \V4/V1/A2/A1/M1/s1 ;
 wire \V4/V1/A2/A1/M2/c1 ;
 wire \V4/V1/A2/A1/M2/c2 ;
 wire \V4/V1/A2/A1/M2/s1 ;
 wire \V4/V1/A2/A1/M3/c1 ;
 wire \V4/V1/A2/A1/M3/c2 ;
 wire \V4/V1/A2/A1/M3/s1 ;
 wire \V4/V1/A2/A1/M4/c1 ;
 wire \V4/V1/A2/A1/M4/c2 ;
 wire \V4/V1/A2/A1/M4/s1 ;
 wire \V4/V1/A2/A2/c1 ;
 wire \V4/V1/A2/A2/c2 ;
 wire \V4/V1/A2/A2/c3 ;
 wire \V4/V1/A2/A2/M1/c1 ;
 wire \V4/V1/A2/A2/M1/c2 ;
 wire \V4/V1/A2/A2/M1/s1 ;
 wire \V4/V1/A2/A2/M2/c1 ;
 wire \V4/V1/A2/A2/M2/c2 ;
 wire \V4/V1/A2/A2/M2/s1 ;
 wire \V4/V1/A2/A2/M3/c1 ;
 wire \V4/V1/A2/A2/M3/c2 ;
 wire \V4/V1/A2/A2/M3/s1 ;
 wire \V4/V1/A2/A2/M4/c1 ;
 wire \V4/V1/A2/A2/M4/c2 ;
 wire \V4/V1/A2/A2/M4/s1 ;
 wire \V4/V1/A3/c1 ;
 wire \V4/V1/A3/A1/c1 ;
 wire \V4/V1/A3/A1/c2 ;
 wire \V4/V1/A3/A1/c3 ;
 wire \V4/V1/A3/A1/M1/c1 ;
 wire \V4/V1/A3/A1/M1/c2 ;
 wire \V4/V1/A3/A1/M1/s1 ;
 wire \V4/V1/A3/A1/M2/c1 ;
 wire \V4/V1/A3/A1/M2/c2 ;
 wire \V4/V1/A3/A1/M2/s1 ;
 wire \V4/V1/A3/A1/M3/c1 ;
 wire \V4/V1/A3/A1/M3/c2 ;
 wire \V4/V1/A3/A1/M3/s1 ;
 wire \V4/V1/A3/A1/M4/c1 ;
 wire \V4/V1/A3/A1/M4/c2 ;
 wire \V4/V1/A3/A1/M4/s1 ;
 wire \V4/V1/A3/A2/c1 ;
 wire \V4/V1/A3/A2/c2 ;
 wire \V4/V1/A3/A2/c3 ;
 wire \V4/V1/A3/A2/M1/c1 ;
 wire \V4/V1/A3/A2/M1/c2 ;
 wire \V4/V1/A3/A2/M1/s1 ;
 wire \V4/V1/A3/A2/M2/c1 ;
 wire \V4/V1/A3/A2/M2/c2 ;
 wire \V4/V1/A3/A2/M2/s1 ;
 wire \V4/V1/A3/A2/M3/c1 ;
 wire \V4/V1/A3/A2/M3/c2 ;
 wire \V4/V1/A3/A2/M3/s1 ;
 wire \V4/V1/A3/A2/M4/c1 ;
 wire \V4/V1/A3/A2/M4/c2 ;
 wire \V4/V1/A3/A2/M4/s1 ;
 wire \V4/V1/V1/c1 ;
 wire \V4/V1/V1/c2 ;
 wire \V4/V1/V1/c3 ;
 wire \V4/V1/V1/overflow ;
 wire \V4/V1/V1/A1/c1 ;
 wire \V4/V1/V1/A1/c2 ;
 wire \V4/V1/V1/A1/c3 ;
 wire \V4/V1/V1/A1/M1/c1 ;
 wire \V4/V1/V1/A1/M1/c2 ;
 wire \V4/V1/V1/A1/M1/s1 ;
 wire \V4/V1/V1/A1/M2/c1 ;
 wire \V4/V1/V1/A1/M2/c2 ;
 wire \V4/V1/V1/A1/M2/s1 ;
 wire \V4/V1/V1/A1/M3/c1 ;
 wire \V4/V1/V1/A1/M3/c2 ;
 wire \V4/V1/V1/A1/M3/s1 ;
 wire \V4/V1/V1/A1/M4/c1 ;
 wire \V4/V1/V1/A1/M4/c2 ;
 wire \V4/V1/V1/A1/M4/s1 ;
 wire \V4/V1/V1/A2/c1 ;
 wire \V4/V1/V1/A2/c2 ;
 wire \V4/V1/V1/A2/c3 ;
 wire \V4/V1/V1/A2/M1/c1 ;
 wire \V4/V1/V1/A2/M1/c2 ;
 wire \V4/V1/V1/A2/M1/s1 ;
 wire \V4/V1/V1/A2/M2/c1 ;
 wire \V4/V1/V1/A2/M2/c2 ;
 wire \V4/V1/V1/A2/M2/s1 ;
 wire \V4/V1/V1/A2/M3/c1 ;
 wire \V4/V1/V1/A2/M3/c2 ;
 wire \V4/V1/V1/A2/M3/s1 ;
 wire \V4/V1/V1/A2/M4/c1 ;
 wire \V4/V1/V1/A2/M4/c2 ;
 wire \V4/V1/V1/A2/M4/s1 ;
 wire \V4/V1/V1/A3/c1 ;
 wire \V4/V1/V1/A3/c2 ;
 wire \V4/V1/V1/A3/c3 ;
 wire \V4/V1/V1/A3/M1/c1 ;
 wire \V4/V1/V1/A3/M1/c2 ;
 wire \V4/V1/V1/A3/M1/s1 ;
 wire \V4/V1/V1/A3/M2/c1 ;
 wire \V4/V1/V1/A3/M2/c2 ;
 wire \V4/V1/V1/A3/M2/s1 ;
 wire \V4/V1/V1/A3/M3/c1 ;
 wire \V4/V1/V1/A3/M3/c2 ;
 wire \V4/V1/V1/A3/M3/s1 ;
 wire \V4/V1/V1/A3/M4/c1 ;
 wire \V4/V1/V1/A3/M4/c2 ;
 wire \V4/V1/V1/A3/M4/s1 ;
 wire \V4/V1/V1/V1/w1 ;
 wire \V4/V1/V1/V1/w2 ;
 wire \V4/V1/V1/V1/w3 ;
 wire \V4/V1/V1/V1/w4 ;
 wire \V4/V1/V1/V2/w1 ;
 wire \V4/V1/V1/V2/w2 ;
 wire \V4/V1/V1/V2/w3 ;
 wire \V4/V1/V1/V2/w4 ;
 wire \V4/V1/V1/V3/w1 ;
 wire \V4/V1/V1/V3/w2 ;
 wire \V4/V1/V1/V3/w3 ;
 wire \V4/V1/V1/V3/w4 ;
 wire \V4/V1/V1/V4/w1 ;
 wire \V4/V1/V1/V4/w2 ;
 wire \V4/V1/V1/V4/w3 ;
 wire \V4/V1/V1/V4/w4 ;
 wire \V4/V1/V2/c1 ;
 wire \V4/V1/V2/c2 ;
 wire \V4/V1/V2/c3 ;
 wire \V4/V1/V2/overflow ;
 wire \V4/V1/V2/A1/c1 ;
 wire \V4/V1/V2/A1/c2 ;
 wire \V4/V1/V2/A1/c3 ;
 wire \V4/V1/V2/A1/M1/c1 ;
 wire \V4/V1/V2/A1/M1/c2 ;
 wire \V4/V1/V2/A1/M1/s1 ;
 wire \V4/V1/V2/A1/M2/c1 ;
 wire \V4/V1/V2/A1/M2/c2 ;
 wire \V4/V1/V2/A1/M2/s1 ;
 wire \V4/V1/V2/A1/M3/c1 ;
 wire \V4/V1/V2/A1/M3/c2 ;
 wire \V4/V1/V2/A1/M3/s1 ;
 wire \V4/V1/V2/A1/M4/c1 ;
 wire \V4/V1/V2/A1/M4/c2 ;
 wire \V4/V1/V2/A1/M4/s1 ;
 wire \V4/V1/V2/A2/c1 ;
 wire \V4/V1/V2/A2/c2 ;
 wire \V4/V1/V2/A2/c3 ;
 wire \V4/V1/V2/A2/M1/c1 ;
 wire \V4/V1/V2/A2/M1/c2 ;
 wire \V4/V1/V2/A2/M1/s1 ;
 wire \V4/V1/V2/A2/M2/c1 ;
 wire \V4/V1/V2/A2/M2/c2 ;
 wire \V4/V1/V2/A2/M2/s1 ;
 wire \V4/V1/V2/A2/M3/c1 ;
 wire \V4/V1/V2/A2/M3/c2 ;
 wire \V4/V1/V2/A2/M3/s1 ;
 wire \V4/V1/V2/A2/M4/c1 ;
 wire \V4/V1/V2/A2/M4/c2 ;
 wire \V4/V1/V2/A2/M4/s1 ;
 wire \V4/V1/V2/A3/c1 ;
 wire \V4/V1/V2/A3/c2 ;
 wire \V4/V1/V2/A3/c3 ;
 wire \V4/V1/V2/A3/M1/c1 ;
 wire \V4/V1/V2/A3/M1/c2 ;
 wire \V4/V1/V2/A3/M1/s1 ;
 wire \V4/V1/V2/A3/M2/c1 ;
 wire \V4/V1/V2/A3/M2/c2 ;
 wire \V4/V1/V2/A3/M2/s1 ;
 wire \V4/V1/V2/A3/M3/c1 ;
 wire \V4/V1/V2/A3/M3/c2 ;
 wire \V4/V1/V2/A3/M3/s1 ;
 wire \V4/V1/V2/A3/M4/c1 ;
 wire \V4/V1/V2/A3/M4/c2 ;
 wire \V4/V1/V2/A3/M4/s1 ;
 wire \V4/V1/V2/V1/w1 ;
 wire \V4/V1/V2/V1/w2 ;
 wire \V4/V1/V2/V1/w3 ;
 wire \V4/V1/V2/V1/w4 ;
 wire \V4/V1/V2/V2/w1 ;
 wire \V4/V1/V2/V2/w2 ;
 wire \V4/V1/V2/V2/w3 ;
 wire \V4/V1/V2/V2/w4 ;
 wire \V4/V1/V2/V3/w1 ;
 wire \V4/V1/V2/V3/w2 ;
 wire \V4/V1/V2/V3/w3 ;
 wire \V4/V1/V2/V3/w4 ;
 wire \V4/V1/V2/V4/w1 ;
 wire \V4/V1/V2/V4/w2 ;
 wire \V4/V1/V2/V4/w3 ;
 wire \V4/V1/V2/V4/w4 ;
 wire \V4/V1/V3/c1 ;
 wire \V4/V1/V3/c2 ;
 wire \V4/V1/V3/c3 ;
 wire \V4/V1/V3/overflow ;
 wire \V4/V1/V3/A1/c1 ;
 wire \V4/V1/V3/A1/c2 ;
 wire \V4/V1/V3/A1/c3 ;
 wire \V4/V1/V3/A1/M1/c1 ;
 wire \V4/V1/V3/A1/M1/c2 ;
 wire \V4/V1/V3/A1/M1/s1 ;
 wire \V4/V1/V3/A1/M2/c1 ;
 wire \V4/V1/V3/A1/M2/c2 ;
 wire \V4/V1/V3/A1/M2/s1 ;
 wire \V4/V1/V3/A1/M3/c1 ;
 wire \V4/V1/V3/A1/M3/c2 ;
 wire \V4/V1/V3/A1/M3/s1 ;
 wire \V4/V1/V3/A1/M4/c1 ;
 wire \V4/V1/V3/A1/M4/c2 ;
 wire \V4/V1/V3/A1/M4/s1 ;
 wire \V4/V1/V3/A2/c1 ;
 wire \V4/V1/V3/A2/c2 ;
 wire \V4/V1/V3/A2/c3 ;
 wire \V4/V1/V3/A2/M1/c1 ;
 wire \V4/V1/V3/A2/M1/c2 ;
 wire \V4/V1/V3/A2/M1/s1 ;
 wire \V4/V1/V3/A2/M2/c1 ;
 wire \V4/V1/V3/A2/M2/c2 ;
 wire \V4/V1/V3/A2/M2/s1 ;
 wire \V4/V1/V3/A2/M3/c1 ;
 wire \V4/V1/V3/A2/M3/c2 ;
 wire \V4/V1/V3/A2/M3/s1 ;
 wire \V4/V1/V3/A2/M4/c1 ;
 wire \V4/V1/V3/A2/M4/c2 ;
 wire \V4/V1/V3/A2/M4/s1 ;
 wire \V4/V1/V3/A3/c1 ;
 wire \V4/V1/V3/A3/c2 ;
 wire \V4/V1/V3/A3/c3 ;
 wire \V4/V1/V3/A3/M1/c1 ;
 wire \V4/V1/V3/A3/M1/c2 ;
 wire \V4/V1/V3/A3/M1/s1 ;
 wire \V4/V1/V3/A3/M2/c1 ;
 wire \V4/V1/V3/A3/M2/c2 ;
 wire \V4/V1/V3/A3/M2/s1 ;
 wire \V4/V1/V3/A3/M3/c1 ;
 wire \V4/V1/V3/A3/M3/c2 ;
 wire \V4/V1/V3/A3/M3/s1 ;
 wire \V4/V1/V3/A3/M4/c1 ;
 wire \V4/V1/V3/A3/M4/c2 ;
 wire \V4/V1/V3/A3/M4/s1 ;
 wire \V4/V1/V3/V1/w1 ;
 wire \V4/V1/V3/V1/w2 ;
 wire \V4/V1/V3/V1/w3 ;
 wire \V4/V1/V3/V1/w4 ;
 wire \V4/V1/V3/V2/w1 ;
 wire \V4/V1/V3/V2/w2 ;
 wire \V4/V1/V3/V2/w3 ;
 wire \V4/V1/V3/V2/w4 ;
 wire \V4/V1/V3/V3/w1 ;
 wire \V4/V1/V3/V3/w2 ;
 wire \V4/V1/V3/V3/w3 ;
 wire \V4/V1/V3/V3/w4 ;
 wire \V4/V1/V3/V4/w1 ;
 wire \V4/V1/V3/V4/w2 ;
 wire \V4/V1/V3/V4/w3 ;
 wire \V4/V1/V3/V4/w4 ;
 wire \V4/V1/V4/c1 ;
 wire \V4/V1/V4/c2 ;
 wire \V4/V1/V4/c3 ;
 wire \V4/V1/V4/overflow ;
 wire \V4/V1/V4/A1/c1 ;
 wire \V4/V1/V4/A1/c2 ;
 wire \V4/V1/V4/A1/c3 ;
 wire \V4/V1/V4/A1/M1/c1 ;
 wire \V4/V1/V4/A1/M1/c2 ;
 wire \V4/V1/V4/A1/M1/s1 ;
 wire \V4/V1/V4/A1/M2/c1 ;
 wire \V4/V1/V4/A1/M2/c2 ;
 wire \V4/V1/V4/A1/M2/s1 ;
 wire \V4/V1/V4/A1/M3/c1 ;
 wire \V4/V1/V4/A1/M3/c2 ;
 wire \V4/V1/V4/A1/M3/s1 ;
 wire \V4/V1/V4/A1/M4/c1 ;
 wire \V4/V1/V4/A1/M4/c2 ;
 wire \V4/V1/V4/A1/M4/s1 ;
 wire \V4/V1/V4/A2/c1 ;
 wire \V4/V1/V4/A2/c2 ;
 wire \V4/V1/V4/A2/c3 ;
 wire \V4/V1/V4/A2/M1/c1 ;
 wire \V4/V1/V4/A2/M1/c2 ;
 wire \V4/V1/V4/A2/M1/s1 ;
 wire \V4/V1/V4/A2/M2/c1 ;
 wire \V4/V1/V4/A2/M2/c2 ;
 wire \V4/V1/V4/A2/M2/s1 ;
 wire \V4/V1/V4/A2/M3/c1 ;
 wire \V4/V1/V4/A2/M3/c2 ;
 wire \V4/V1/V4/A2/M3/s1 ;
 wire \V4/V1/V4/A2/M4/c1 ;
 wire \V4/V1/V4/A2/M4/c2 ;
 wire \V4/V1/V4/A2/M4/s1 ;
 wire \V4/V1/V4/A3/c1 ;
 wire \V4/V1/V4/A3/c2 ;
 wire \V4/V1/V4/A3/c3 ;
 wire \V4/V1/V4/A3/M1/c1 ;
 wire \V4/V1/V4/A3/M1/c2 ;
 wire \V4/V1/V4/A3/M1/s1 ;
 wire \V4/V1/V4/A3/M2/c1 ;
 wire \V4/V1/V4/A3/M2/c2 ;
 wire \V4/V1/V4/A3/M2/s1 ;
 wire \V4/V1/V4/A3/M3/c1 ;
 wire \V4/V1/V4/A3/M3/c2 ;
 wire \V4/V1/V4/A3/M3/s1 ;
 wire \V4/V1/V4/A3/M4/c1 ;
 wire \V4/V1/V4/A3/M4/c2 ;
 wire \V4/V1/V4/A3/M4/s1 ;
 wire \V4/V1/V4/V1/w1 ;
 wire \V4/V1/V4/V1/w2 ;
 wire \V4/V1/V4/V1/w3 ;
 wire \V4/V1/V4/V1/w4 ;
 wire \V4/V1/V4/V2/w1 ;
 wire \V4/V1/V4/V2/w2 ;
 wire \V4/V1/V4/V2/w3 ;
 wire \V4/V1/V4/V2/w4 ;
 wire \V4/V1/V4/V3/w1 ;
 wire \V4/V1/V4/V3/w2 ;
 wire \V4/V1/V4/V3/w3 ;
 wire \V4/V1/V4/V3/w4 ;
 wire \V4/V1/V4/V4/w1 ;
 wire \V4/V1/V4/V4/w2 ;
 wire \V4/V1/V4/V4/w3 ;
 wire \V4/V1/V4/V4/w4 ;
 wire \V4/V2/c1 ;
 wire \V4/V2/c2 ;
 wire \V4/V2/c3 ;
 wire \V4/V2/overflow ;
 wire \V4/V2/A1/c1 ;
 wire \V4/V2/A1/A1/c1 ;
 wire \V4/V2/A1/A1/c2 ;
 wire \V4/V2/A1/A1/c3 ;
 wire \V4/V2/A1/A1/M1/c1 ;
 wire \V4/V2/A1/A1/M1/c2 ;
 wire \V4/V2/A1/A1/M1/s1 ;
 wire \V4/V2/A1/A1/M2/c1 ;
 wire \V4/V2/A1/A1/M2/c2 ;
 wire \V4/V2/A1/A1/M2/s1 ;
 wire \V4/V2/A1/A1/M3/c1 ;
 wire \V4/V2/A1/A1/M3/c2 ;
 wire \V4/V2/A1/A1/M3/s1 ;
 wire \V4/V2/A1/A1/M4/c1 ;
 wire \V4/V2/A1/A1/M4/c2 ;
 wire \V4/V2/A1/A1/M4/s1 ;
 wire \V4/V2/A1/A2/c1 ;
 wire \V4/V2/A1/A2/c2 ;
 wire \V4/V2/A1/A2/c3 ;
 wire \V4/V2/A1/A2/M1/c1 ;
 wire \V4/V2/A1/A2/M1/c2 ;
 wire \V4/V2/A1/A2/M1/s1 ;
 wire \V4/V2/A1/A2/M2/c1 ;
 wire \V4/V2/A1/A2/M2/c2 ;
 wire \V4/V2/A1/A2/M2/s1 ;
 wire \V4/V2/A1/A2/M3/c1 ;
 wire \V4/V2/A1/A2/M3/c2 ;
 wire \V4/V2/A1/A2/M3/s1 ;
 wire \V4/V2/A1/A2/M4/c1 ;
 wire \V4/V2/A1/A2/M4/c2 ;
 wire \V4/V2/A1/A2/M4/s1 ;
 wire \V4/V2/A2/c1 ;
 wire \V4/V2/A2/A1/c1 ;
 wire \V4/V2/A2/A1/c2 ;
 wire \V4/V2/A2/A1/c3 ;
 wire \V4/V2/A2/A1/M1/c1 ;
 wire \V4/V2/A2/A1/M1/c2 ;
 wire \V4/V2/A2/A1/M1/s1 ;
 wire \V4/V2/A2/A1/M2/c1 ;
 wire \V4/V2/A2/A1/M2/c2 ;
 wire \V4/V2/A2/A1/M2/s1 ;
 wire \V4/V2/A2/A1/M3/c1 ;
 wire \V4/V2/A2/A1/M3/c2 ;
 wire \V4/V2/A2/A1/M3/s1 ;
 wire \V4/V2/A2/A1/M4/c1 ;
 wire \V4/V2/A2/A1/M4/c2 ;
 wire \V4/V2/A2/A1/M4/s1 ;
 wire \V4/V2/A2/A2/c1 ;
 wire \V4/V2/A2/A2/c2 ;
 wire \V4/V2/A2/A2/c3 ;
 wire \V4/V2/A2/A2/M1/c1 ;
 wire \V4/V2/A2/A2/M1/c2 ;
 wire \V4/V2/A2/A2/M1/s1 ;
 wire \V4/V2/A2/A2/M2/c1 ;
 wire \V4/V2/A2/A2/M2/c2 ;
 wire \V4/V2/A2/A2/M2/s1 ;
 wire \V4/V2/A2/A2/M3/c1 ;
 wire \V4/V2/A2/A2/M3/c2 ;
 wire \V4/V2/A2/A2/M3/s1 ;
 wire \V4/V2/A2/A2/M4/c1 ;
 wire \V4/V2/A2/A2/M4/c2 ;
 wire \V4/V2/A2/A2/M4/s1 ;
 wire \V4/V2/A3/c1 ;
 wire \V4/V2/A3/A1/c1 ;
 wire \V4/V2/A3/A1/c2 ;
 wire \V4/V2/A3/A1/c3 ;
 wire \V4/V2/A3/A1/M1/c1 ;
 wire \V4/V2/A3/A1/M1/c2 ;
 wire \V4/V2/A3/A1/M1/s1 ;
 wire \V4/V2/A3/A1/M2/c1 ;
 wire \V4/V2/A3/A1/M2/c2 ;
 wire \V4/V2/A3/A1/M2/s1 ;
 wire \V4/V2/A3/A1/M3/c1 ;
 wire \V4/V2/A3/A1/M3/c2 ;
 wire \V4/V2/A3/A1/M3/s1 ;
 wire \V4/V2/A3/A1/M4/c1 ;
 wire \V4/V2/A3/A1/M4/c2 ;
 wire \V4/V2/A3/A1/M4/s1 ;
 wire \V4/V2/A3/A2/c1 ;
 wire \V4/V2/A3/A2/c2 ;
 wire \V4/V2/A3/A2/c3 ;
 wire \V4/V2/A3/A2/M1/c1 ;
 wire \V4/V2/A3/A2/M1/c2 ;
 wire \V4/V2/A3/A2/M1/s1 ;
 wire \V4/V2/A3/A2/M2/c1 ;
 wire \V4/V2/A3/A2/M2/c2 ;
 wire \V4/V2/A3/A2/M2/s1 ;
 wire \V4/V2/A3/A2/M3/c1 ;
 wire \V4/V2/A3/A2/M3/c2 ;
 wire \V4/V2/A3/A2/M3/s1 ;
 wire \V4/V2/A3/A2/M4/c1 ;
 wire \V4/V2/A3/A2/M4/c2 ;
 wire \V4/V2/A3/A2/M4/s1 ;
 wire \V4/V2/V1/c1 ;
 wire \V4/V2/V1/c2 ;
 wire \V4/V2/V1/c3 ;
 wire \V4/V2/V1/overflow ;
 wire \V4/V2/V1/A1/c1 ;
 wire \V4/V2/V1/A1/c2 ;
 wire \V4/V2/V1/A1/c3 ;
 wire \V4/V2/V1/A1/M1/c1 ;
 wire \V4/V2/V1/A1/M1/c2 ;
 wire \V4/V2/V1/A1/M1/s1 ;
 wire \V4/V2/V1/A1/M2/c1 ;
 wire \V4/V2/V1/A1/M2/c2 ;
 wire \V4/V2/V1/A1/M2/s1 ;
 wire \V4/V2/V1/A1/M3/c1 ;
 wire \V4/V2/V1/A1/M3/c2 ;
 wire \V4/V2/V1/A1/M3/s1 ;
 wire \V4/V2/V1/A1/M4/c1 ;
 wire \V4/V2/V1/A1/M4/c2 ;
 wire \V4/V2/V1/A1/M4/s1 ;
 wire \V4/V2/V1/A2/c1 ;
 wire \V4/V2/V1/A2/c2 ;
 wire \V4/V2/V1/A2/c3 ;
 wire \V4/V2/V1/A2/M1/c1 ;
 wire \V4/V2/V1/A2/M1/c2 ;
 wire \V4/V2/V1/A2/M1/s1 ;
 wire \V4/V2/V1/A2/M2/c1 ;
 wire \V4/V2/V1/A2/M2/c2 ;
 wire \V4/V2/V1/A2/M2/s1 ;
 wire \V4/V2/V1/A2/M3/c1 ;
 wire \V4/V2/V1/A2/M3/c2 ;
 wire \V4/V2/V1/A2/M3/s1 ;
 wire \V4/V2/V1/A2/M4/c1 ;
 wire \V4/V2/V1/A2/M4/c2 ;
 wire \V4/V2/V1/A2/M4/s1 ;
 wire \V4/V2/V1/A3/c1 ;
 wire \V4/V2/V1/A3/c2 ;
 wire \V4/V2/V1/A3/c3 ;
 wire \V4/V2/V1/A3/M1/c1 ;
 wire \V4/V2/V1/A3/M1/c2 ;
 wire \V4/V2/V1/A3/M1/s1 ;
 wire \V4/V2/V1/A3/M2/c1 ;
 wire \V4/V2/V1/A3/M2/c2 ;
 wire \V4/V2/V1/A3/M2/s1 ;
 wire \V4/V2/V1/A3/M3/c1 ;
 wire \V4/V2/V1/A3/M3/c2 ;
 wire \V4/V2/V1/A3/M3/s1 ;
 wire \V4/V2/V1/A3/M4/c1 ;
 wire \V4/V2/V1/A3/M4/c2 ;
 wire \V4/V2/V1/A3/M4/s1 ;
 wire \V4/V2/V1/V1/w1 ;
 wire \V4/V2/V1/V1/w2 ;
 wire \V4/V2/V1/V1/w3 ;
 wire \V4/V2/V1/V1/w4 ;
 wire \V4/V2/V1/V2/w1 ;
 wire \V4/V2/V1/V2/w2 ;
 wire \V4/V2/V1/V2/w3 ;
 wire \V4/V2/V1/V2/w4 ;
 wire \V4/V2/V1/V3/w1 ;
 wire \V4/V2/V1/V3/w2 ;
 wire \V4/V2/V1/V3/w3 ;
 wire \V4/V2/V1/V3/w4 ;
 wire \V4/V2/V1/V4/w1 ;
 wire \V4/V2/V1/V4/w2 ;
 wire \V4/V2/V1/V4/w3 ;
 wire \V4/V2/V1/V4/w4 ;
 wire \V4/V2/V2/c1 ;
 wire \V4/V2/V2/c2 ;
 wire \V4/V2/V2/c3 ;
 wire \V4/V2/V2/overflow ;
 wire \V4/V2/V2/A1/c1 ;
 wire \V4/V2/V2/A1/c2 ;
 wire \V4/V2/V2/A1/c3 ;
 wire \V4/V2/V2/A1/M1/c1 ;
 wire \V4/V2/V2/A1/M1/c2 ;
 wire \V4/V2/V2/A1/M1/s1 ;
 wire \V4/V2/V2/A1/M2/c1 ;
 wire \V4/V2/V2/A1/M2/c2 ;
 wire \V4/V2/V2/A1/M2/s1 ;
 wire \V4/V2/V2/A1/M3/c1 ;
 wire \V4/V2/V2/A1/M3/c2 ;
 wire \V4/V2/V2/A1/M3/s1 ;
 wire \V4/V2/V2/A1/M4/c1 ;
 wire \V4/V2/V2/A1/M4/c2 ;
 wire \V4/V2/V2/A1/M4/s1 ;
 wire \V4/V2/V2/A2/c1 ;
 wire \V4/V2/V2/A2/c2 ;
 wire \V4/V2/V2/A2/c3 ;
 wire \V4/V2/V2/A2/M1/c1 ;
 wire \V4/V2/V2/A2/M1/c2 ;
 wire \V4/V2/V2/A2/M1/s1 ;
 wire \V4/V2/V2/A2/M2/c1 ;
 wire \V4/V2/V2/A2/M2/c2 ;
 wire \V4/V2/V2/A2/M2/s1 ;
 wire \V4/V2/V2/A2/M3/c1 ;
 wire \V4/V2/V2/A2/M3/c2 ;
 wire \V4/V2/V2/A2/M3/s1 ;
 wire \V4/V2/V2/A2/M4/c1 ;
 wire \V4/V2/V2/A2/M4/c2 ;
 wire \V4/V2/V2/A2/M4/s1 ;
 wire \V4/V2/V2/A3/c1 ;
 wire \V4/V2/V2/A3/c2 ;
 wire \V4/V2/V2/A3/c3 ;
 wire \V4/V2/V2/A3/M1/c1 ;
 wire \V4/V2/V2/A3/M1/c2 ;
 wire \V4/V2/V2/A3/M1/s1 ;
 wire \V4/V2/V2/A3/M2/c1 ;
 wire \V4/V2/V2/A3/M2/c2 ;
 wire \V4/V2/V2/A3/M2/s1 ;
 wire \V4/V2/V2/A3/M3/c1 ;
 wire \V4/V2/V2/A3/M3/c2 ;
 wire \V4/V2/V2/A3/M3/s1 ;
 wire \V4/V2/V2/A3/M4/c1 ;
 wire \V4/V2/V2/A3/M4/c2 ;
 wire \V4/V2/V2/A3/M4/s1 ;
 wire \V4/V2/V2/V1/w1 ;
 wire \V4/V2/V2/V1/w2 ;
 wire \V4/V2/V2/V1/w3 ;
 wire \V4/V2/V2/V1/w4 ;
 wire \V4/V2/V2/V2/w1 ;
 wire \V4/V2/V2/V2/w2 ;
 wire \V4/V2/V2/V2/w3 ;
 wire \V4/V2/V2/V2/w4 ;
 wire \V4/V2/V2/V3/w1 ;
 wire \V4/V2/V2/V3/w2 ;
 wire \V4/V2/V2/V3/w3 ;
 wire \V4/V2/V2/V3/w4 ;
 wire \V4/V2/V2/V4/w1 ;
 wire \V4/V2/V2/V4/w2 ;
 wire \V4/V2/V2/V4/w3 ;
 wire \V4/V2/V2/V4/w4 ;
 wire \V4/V2/V3/c1 ;
 wire \V4/V2/V3/c2 ;
 wire \V4/V2/V3/c3 ;
 wire \V4/V2/V3/overflow ;
 wire \V4/V2/V3/A1/c1 ;
 wire \V4/V2/V3/A1/c2 ;
 wire \V4/V2/V3/A1/c3 ;
 wire \V4/V2/V3/A1/M1/c1 ;
 wire \V4/V2/V3/A1/M1/c2 ;
 wire \V4/V2/V3/A1/M1/s1 ;
 wire \V4/V2/V3/A1/M2/c1 ;
 wire \V4/V2/V3/A1/M2/c2 ;
 wire \V4/V2/V3/A1/M2/s1 ;
 wire \V4/V2/V3/A1/M3/c1 ;
 wire \V4/V2/V3/A1/M3/c2 ;
 wire \V4/V2/V3/A1/M3/s1 ;
 wire \V4/V2/V3/A1/M4/c1 ;
 wire \V4/V2/V3/A1/M4/c2 ;
 wire \V4/V2/V3/A1/M4/s1 ;
 wire \V4/V2/V3/A2/c1 ;
 wire \V4/V2/V3/A2/c2 ;
 wire \V4/V2/V3/A2/c3 ;
 wire \V4/V2/V3/A2/M1/c1 ;
 wire \V4/V2/V3/A2/M1/c2 ;
 wire \V4/V2/V3/A2/M1/s1 ;
 wire \V4/V2/V3/A2/M2/c1 ;
 wire \V4/V2/V3/A2/M2/c2 ;
 wire \V4/V2/V3/A2/M2/s1 ;
 wire \V4/V2/V3/A2/M3/c1 ;
 wire \V4/V2/V3/A2/M3/c2 ;
 wire \V4/V2/V3/A2/M3/s1 ;
 wire \V4/V2/V3/A2/M4/c1 ;
 wire \V4/V2/V3/A2/M4/c2 ;
 wire \V4/V2/V3/A2/M4/s1 ;
 wire \V4/V2/V3/A3/c1 ;
 wire \V4/V2/V3/A3/c2 ;
 wire \V4/V2/V3/A3/c3 ;
 wire \V4/V2/V3/A3/M1/c1 ;
 wire \V4/V2/V3/A3/M1/c2 ;
 wire \V4/V2/V3/A3/M1/s1 ;
 wire \V4/V2/V3/A3/M2/c1 ;
 wire \V4/V2/V3/A3/M2/c2 ;
 wire \V4/V2/V3/A3/M2/s1 ;
 wire \V4/V2/V3/A3/M3/c1 ;
 wire \V4/V2/V3/A3/M3/c2 ;
 wire \V4/V2/V3/A3/M3/s1 ;
 wire \V4/V2/V3/A3/M4/c1 ;
 wire \V4/V2/V3/A3/M4/c2 ;
 wire \V4/V2/V3/A3/M4/s1 ;
 wire \V4/V2/V3/V1/w1 ;
 wire \V4/V2/V3/V1/w2 ;
 wire \V4/V2/V3/V1/w3 ;
 wire \V4/V2/V3/V1/w4 ;
 wire \V4/V2/V3/V2/w1 ;
 wire \V4/V2/V3/V2/w2 ;
 wire \V4/V2/V3/V2/w3 ;
 wire \V4/V2/V3/V2/w4 ;
 wire \V4/V2/V3/V3/w1 ;
 wire \V4/V2/V3/V3/w2 ;
 wire \V4/V2/V3/V3/w3 ;
 wire \V4/V2/V3/V3/w4 ;
 wire \V4/V2/V3/V4/w1 ;
 wire \V4/V2/V3/V4/w2 ;
 wire \V4/V2/V3/V4/w3 ;
 wire \V4/V2/V3/V4/w4 ;
 wire \V4/V2/V4/c1 ;
 wire \V4/V2/V4/c2 ;
 wire \V4/V2/V4/c3 ;
 wire \V4/V2/V4/overflow ;
 wire \V4/V2/V4/A1/c1 ;
 wire \V4/V2/V4/A1/c2 ;
 wire \V4/V2/V4/A1/c3 ;
 wire \V4/V2/V4/A1/M1/c1 ;
 wire \V4/V2/V4/A1/M1/c2 ;
 wire \V4/V2/V4/A1/M1/s1 ;
 wire \V4/V2/V4/A1/M2/c1 ;
 wire \V4/V2/V4/A1/M2/c2 ;
 wire \V4/V2/V4/A1/M2/s1 ;
 wire \V4/V2/V4/A1/M3/c1 ;
 wire \V4/V2/V4/A1/M3/c2 ;
 wire \V4/V2/V4/A1/M3/s1 ;
 wire \V4/V2/V4/A1/M4/c1 ;
 wire \V4/V2/V4/A1/M4/c2 ;
 wire \V4/V2/V4/A1/M4/s1 ;
 wire \V4/V2/V4/A2/c1 ;
 wire \V4/V2/V4/A2/c2 ;
 wire \V4/V2/V4/A2/c3 ;
 wire \V4/V2/V4/A2/M1/c1 ;
 wire \V4/V2/V4/A2/M1/c2 ;
 wire \V4/V2/V4/A2/M1/s1 ;
 wire \V4/V2/V4/A2/M2/c1 ;
 wire \V4/V2/V4/A2/M2/c2 ;
 wire \V4/V2/V4/A2/M2/s1 ;
 wire \V4/V2/V4/A2/M3/c1 ;
 wire \V4/V2/V4/A2/M3/c2 ;
 wire \V4/V2/V4/A2/M3/s1 ;
 wire \V4/V2/V4/A2/M4/c1 ;
 wire \V4/V2/V4/A2/M4/c2 ;
 wire \V4/V2/V4/A2/M4/s1 ;
 wire \V4/V2/V4/A3/c1 ;
 wire \V4/V2/V4/A3/c2 ;
 wire \V4/V2/V4/A3/c3 ;
 wire \V4/V2/V4/A3/M1/c1 ;
 wire \V4/V2/V4/A3/M1/c2 ;
 wire \V4/V2/V4/A3/M1/s1 ;
 wire \V4/V2/V4/A3/M2/c1 ;
 wire \V4/V2/V4/A3/M2/c2 ;
 wire \V4/V2/V4/A3/M2/s1 ;
 wire \V4/V2/V4/A3/M3/c1 ;
 wire \V4/V2/V4/A3/M3/c2 ;
 wire \V4/V2/V4/A3/M3/s1 ;
 wire \V4/V2/V4/A3/M4/c1 ;
 wire \V4/V2/V4/A3/M4/c2 ;
 wire \V4/V2/V4/A3/M4/s1 ;
 wire \V4/V2/V4/V1/w1 ;
 wire \V4/V2/V4/V1/w2 ;
 wire \V4/V2/V4/V1/w3 ;
 wire \V4/V2/V4/V1/w4 ;
 wire \V4/V2/V4/V2/w1 ;
 wire \V4/V2/V4/V2/w2 ;
 wire \V4/V2/V4/V2/w3 ;
 wire \V4/V2/V4/V2/w4 ;
 wire \V4/V2/V4/V3/w1 ;
 wire \V4/V2/V4/V3/w2 ;
 wire \V4/V2/V4/V3/w3 ;
 wire \V4/V2/V4/V3/w4 ;
 wire \V4/V2/V4/V4/w1 ;
 wire \V4/V2/V4/V4/w2 ;
 wire \V4/V2/V4/V4/w3 ;
 wire \V4/V2/V4/V4/w4 ;
 wire \V4/V3/c1 ;
 wire \V4/V3/c2 ;
 wire \V4/V3/c3 ;
 wire \V4/V3/overflow ;
 wire \V4/V3/A1/c1 ;
 wire \V4/V3/A1/A1/c1 ;
 wire \V4/V3/A1/A1/c2 ;
 wire \V4/V3/A1/A1/c3 ;
 wire \V4/V3/A1/A1/M1/c1 ;
 wire \V4/V3/A1/A1/M1/c2 ;
 wire \V4/V3/A1/A1/M1/s1 ;
 wire \V4/V3/A1/A1/M2/c1 ;
 wire \V4/V3/A1/A1/M2/c2 ;
 wire \V4/V3/A1/A1/M2/s1 ;
 wire \V4/V3/A1/A1/M3/c1 ;
 wire \V4/V3/A1/A1/M3/c2 ;
 wire \V4/V3/A1/A1/M3/s1 ;
 wire \V4/V3/A1/A1/M4/c1 ;
 wire \V4/V3/A1/A1/M4/c2 ;
 wire \V4/V3/A1/A1/M4/s1 ;
 wire \V4/V3/A1/A2/c1 ;
 wire \V4/V3/A1/A2/c2 ;
 wire \V4/V3/A1/A2/c3 ;
 wire \V4/V3/A1/A2/M1/c1 ;
 wire \V4/V3/A1/A2/M1/c2 ;
 wire \V4/V3/A1/A2/M1/s1 ;
 wire \V4/V3/A1/A2/M2/c1 ;
 wire \V4/V3/A1/A2/M2/c2 ;
 wire \V4/V3/A1/A2/M2/s1 ;
 wire \V4/V3/A1/A2/M3/c1 ;
 wire \V4/V3/A1/A2/M3/c2 ;
 wire \V4/V3/A1/A2/M3/s1 ;
 wire \V4/V3/A1/A2/M4/c1 ;
 wire \V4/V3/A1/A2/M4/c2 ;
 wire \V4/V3/A1/A2/M4/s1 ;
 wire \V4/V3/A2/c1 ;
 wire \V4/V3/A2/A1/c1 ;
 wire \V4/V3/A2/A1/c2 ;
 wire \V4/V3/A2/A1/c3 ;
 wire \V4/V3/A2/A1/M1/c1 ;
 wire \V4/V3/A2/A1/M1/c2 ;
 wire \V4/V3/A2/A1/M1/s1 ;
 wire \V4/V3/A2/A1/M2/c1 ;
 wire \V4/V3/A2/A1/M2/c2 ;
 wire \V4/V3/A2/A1/M2/s1 ;
 wire \V4/V3/A2/A1/M3/c1 ;
 wire \V4/V3/A2/A1/M3/c2 ;
 wire \V4/V3/A2/A1/M3/s1 ;
 wire \V4/V3/A2/A1/M4/c1 ;
 wire \V4/V3/A2/A1/M4/c2 ;
 wire \V4/V3/A2/A1/M4/s1 ;
 wire \V4/V3/A2/A2/c1 ;
 wire \V4/V3/A2/A2/c2 ;
 wire \V4/V3/A2/A2/c3 ;
 wire \V4/V3/A2/A2/M1/c1 ;
 wire \V4/V3/A2/A2/M1/c2 ;
 wire \V4/V3/A2/A2/M1/s1 ;
 wire \V4/V3/A2/A2/M2/c1 ;
 wire \V4/V3/A2/A2/M2/c2 ;
 wire \V4/V3/A2/A2/M2/s1 ;
 wire \V4/V3/A2/A2/M3/c1 ;
 wire \V4/V3/A2/A2/M3/c2 ;
 wire \V4/V3/A2/A2/M3/s1 ;
 wire \V4/V3/A2/A2/M4/c1 ;
 wire \V4/V3/A2/A2/M4/c2 ;
 wire \V4/V3/A2/A2/M4/s1 ;
 wire \V4/V3/A3/c1 ;
 wire \V4/V3/A3/A1/c1 ;
 wire \V4/V3/A3/A1/c2 ;
 wire \V4/V3/A3/A1/c3 ;
 wire \V4/V3/A3/A1/M1/c1 ;
 wire \V4/V3/A3/A1/M1/c2 ;
 wire \V4/V3/A3/A1/M1/s1 ;
 wire \V4/V3/A3/A1/M2/c1 ;
 wire \V4/V3/A3/A1/M2/c2 ;
 wire \V4/V3/A3/A1/M2/s1 ;
 wire \V4/V3/A3/A1/M3/c1 ;
 wire \V4/V3/A3/A1/M3/c2 ;
 wire \V4/V3/A3/A1/M3/s1 ;
 wire \V4/V3/A3/A1/M4/c1 ;
 wire \V4/V3/A3/A1/M4/c2 ;
 wire \V4/V3/A3/A1/M4/s1 ;
 wire \V4/V3/A3/A2/c1 ;
 wire \V4/V3/A3/A2/c2 ;
 wire \V4/V3/A3/A2/c3 ;
 wire \V4/V3/A3/A2/M1/c1 ;
 wire \V4/V3/A3/A2/M1/c2 ;
 wire \V4/V3/A3/A2/M1/s1 ;
 wire \V4/V3/A3/A2/M2/c1 ;
 wire \V4/V3/A3/A2/M2/c2 ;
 wire \V4/V3/A3/A2/M2/s1 ;
 wire \V4/V3/A3/A2/M3/c1 ;
 wire \V4/V3/A3/A2/M3/c2 ;
 wire \V4/V3/A3/A2/M3/s1 ;
 wire \V4/V3/A3/A2/M4/c1 ;
 wire \V4/V3/A3/A2/M4/c2 ;
 wire \V4/V3/A3/A2/M4/s1 ;
 wire \V4/V3/V1/c1 ;
 wire \V4/V3/V1/c2 ;
 wire \V4/V3/V1/c3 ;
 wire \V4/V3/V1/overflow ;
 wire \V4/V3/V1/A1/c1 ;
 wire \V4/V3/V1/A1/c2 ;
 wire \V4/V3/V1/A1/c3 ;
 wire \V4/V3/V1/A1/M1/c1 ;
 wire \V4/V3/V1/A1/M1/c2 ;
 wire \V4/V3/V1/A1/M1/s1 ;
 wire \V4/V3/V1/A1/M2/c1 ;
 wire \V4/V3/V1/A1/M2/c2 ;
 wire \V4/V3/V1/A1/M2/s1 ;
 wire \V4/V3/V1/A1/M3/c1 ;
 wire \V4/V3/V1/A1/M3/c2 ;
 wire \V4/V3/V1/A1/M3/s1 ;
 wire \V4/V3/V1/A1/M4/c1 ;
 wire \V4/V3/V1/A1/M4/c2 ;
 wire \V4/V3/V1/A1/M4/s1 ;
 wire \V4/V3/V1/A2/c1 ;
 wire \V4/V3/V1/A2/c2 ;
 wire \V4/V3/V1/A2/c3 ;
 wire \V4/V3/V1/A2/M1/c1 ;
 wire \V4/V3/V1/A2/M1/c2 ;
 wire \V4/V3/V1/A2/M1/s1 ;
 wire \V4/V3/V1/A2/M2/c1 ;
 wire \V4/V3/V1/A2/M2/c2 ;
 wire \V4/V3/V1/A2/M2/s1 ;
 wire \V4/V3/V1/A2/M3/c1 ;
 wire \V4/V3/V1/A2/M3/c2 ;
 wire \V4/V3/V1/A2/M3/s1 ;
 wire \V4/V3/V1/A2/M4/c1 ;
 wire \V4/V3/V1/A2/M4/c2 ;
 wire \V4/V3/V1/A2/M4/s1 ;
 wire \V4/V3/V1/A3/c1 ;
 wire \V4/V3/V1/A3/c2 ;
 wire \V4/V3/V1/A3/c3 ;
 wire \V4/V3/V1/A3/M1/c1 ;
 wire \V4/V3/V1/A3/M1/c2 ;
 wire \V4/V3/V1/A3/M1/s1 ;
 wire \V4/V3/V1/A3/M2/c1 ;
 wire \V4/V3/V1/A3/M2/c2 ;
 wire \V4/V3/V1/A3/M2/s1 ;
 wire \V4/V3/V1/A3/M3/c1 ;
 wire \V4/V3/V1/A3/M3/c2 ;
 wire \V4/V3/V1/A3/M3/s1 ;
 wire \V4/V3/V1/A3/M4/c1 ;
 wire \V4/V3/V1/A3/M4/c2 ;
 wire \V4/V3/V1/A3/M4/s1 ;
 wire \V4/V3/V1/V1/w1 ;
 wire \V4/V3/V1/V1/w2 ;
 wire \V4/V3/V1/V1/w3 ;
 wire \V4/V3/V1/V1/w4 ;
 wire \V4/V3/V1/V2/w1 ;
 wire \V4/V3/V1/V2/w2 ;
 wire \V4/V3/V1/V2/w3 ;
 wire \V4/V3/V1/V2/w4 ;
 wire \V4/V3/V1/V3/w1 ;
 wire \V4/V3/V1/V3/w2 ;
 wire \V4/V3/V1/V3/w3 ;
 wire \V4/V3/V1/V3/w4 ;
 wire \V4/V3/V1/V4/w1 ;
 wire \V4/V3/V1/V4/w2 ;
 wire \V4/V3/V1/V4/w3 ;
 wire \V4/V3/V1/V4/w4 ;
 wire \V4/V3/V2/c1 ;
 wire \V4/V3/V2/c2 ;
 wire \V4/V3/V2/c3 ;
 wire \V4/V3/V2/overflow ;
 wire \V4/V3/V2/A1/c1 ;
 wire \V4/V3/V2/A1/c2 ;
 wire \V4/V3/V2/A1/c3 ;
 wire \V4/V3/V2/A1/M1/c1 ;
 wire \V4/V3/V2/A1/M1/c2 ;
 wire \V4/V3/V2/A1/M1/s1 ;
 wire \V4/V3/V2/A1/M2/c1 ;
 wire \V4/V3/V2/A1/M2/c2 ;
 wire \V4/V3/V2/A1/M2/s1 ;
 wire \V4/V3/V2/A1/M3/c1 ;
 wire \V4/V3/V2/A1/M3/c2 ;
 wire \V4/V3/V2/A1/M3/s1 ;
 wire \V4/V3/V2/A1/M4/c1 ;
 wire \V4/V3/V2/A1/M4/c2 ;
 wire \V4/V3/V2/A1/M4/s1 ;
 wire \V4/V3/V2/A2/c1 ;
 wire \V4/V3/V2/A2/c2 ;
 wire \V4/V3/V2/A2/c3 ;
 wire \V4/V3/V2/A2/M1/c1 ;
 wire \V4/V3/V2/A2/M1/c2 ;
 wire \V4/V3/V2/A2/M1/s1 ;
 wire \V4/V3/V2/A2/M2/c1 ;
 wire \V4/V3/V2/A2/M2/c2 ;
 wire \V4/V3/V2/A2/M2/s1 ;
 wire \V4/V3/V2/A2/M3/c1 ;
 wire \V4/V3/V2/A2/M3/c2 ;
 wire \V4/V3/V2/A2/M3/s1 ;
 wire \V4/V3/V2/A2/M4/c1 ;
 wire \V4/V3/V2/A2/M4/c2 ;
 wire \V4/V3/V2/A2/M4/s1 ;
 wire \V4/V3/V2/A3/c1 ;
 wire \V4/V3/V2/A3/c2 ;
 wire \V4/V3/V2/A3/c3 ;
 wire \V4/V3/V2/A3/M1/c1 ;
 wire \V4/V3/V2/A3/M1/c2 ;
 wire \V4/V3/V2/A3/M1/s1 ;
 wire \V4/V3/V2/A3/M2/c1 ;
 wire \V4/V3/V2/A3/M2/c2 ;
 wire \V4/V3/V2/A3/M2/s1 ;
 wire \V4/V3/V2/A3/M3/c1 ;
 wire \V4/V3/V2/A3/M3/c2 ;
 wire \V4/V3/V2/A3/M3/s1 ;
 wire \V4/V3/V2/A3/M4/c1 ;
 wire \V4/V3/V2/A3/M4/c2 ;
 wire \V4/V3/V2/A3/M4/s1 ;
 wire \V4/V3/V2/V1/w1 ;
 wire \V4/V3/V2/V1/w2 ;
 wire \V4/V3/V2/V1/w3 ;
 wire \V4/V3/V2/V1/w4 ;
 wire \V4/V3/V2/V2/w1 ;
 wire \V4/V3/V2/V2/w2 ;
 wire \V4/V3/V2/V2/w3 ;
 wire \V4/V3/V2/V2/w4 ;
 wire \V4/V3/V2/V3/w1 ;
 wire \V4/V3/V2/V3/w2 ;
 wire \V4/V3/V2/V3/w3 ;
 wire \V4/V3/V2/V3/w4 ;
 wire \V4/V3/V2/V4/w1 ;
 wire \V4/V3/V2/V4/w2 ;
 wire \V4/V3/V2/V4/w3 ;
 wire \V4/V3/V2/V4/w4 ;
 wire \V4/V3/V3/c1 ;
 wire \V4/V3/V3/c2 ;
 wire \V4/V3/V3/c3 ;
 wire \V4/V3/V3/overflow ;
 wire \V4/V3/V3/A1/c1 ;
 wire \V4/V3/V3/A1/c2 ;
 wire \V4/V3/V3/A1/c3 ;
 wire \V4/V3/V3/A1/M1/c1 ;
 wire \V4/V3/V3/A1/M1/c2 ;
 wire \V4/V3/V3/A1/M1/s1 ;
 wire \V4/V3/V3/A1/M2/c1 ;
 wire \V4/V3/V3/A1/M2/c2 ;
 wire \V4/V3/V3/A1/M2/s1 ;
 wire \V4/V3/V3/A1/M3/c1 ;
 wire \V4/V3/V3/A1/M3/c2 ;
 wire \V4/V3/V3/A1/M3/s1 ;
 wire \V4/V3/V3/A1/M4/c1 ;
 wire \V4/V3/V3/A1/M4/c2 ;
 wire \V4/V3/V3/A1/M4/s1 ;
 wire \V4/V3/V3/A2/c1 ;
 wire \V4/V3/V3/A2/c2 ;
 wire \V4/V3/V3/A2/c3 ;
 wire \V4/V3/V3/A2/M1/c1 ;
 wire \V4/V3/V3/A2/M1/c2 ;
 wire \V4/V3/V3/A2/M1/s1 ;
 wire \V4/V3/V3/A2/M2/c1 ;
 wire \V4/V3/V3/A2/M2/c2 ;
 wire \V4/V3/V3/A2/M2/s1 ;
 wire \V4/V3/V3/A2/M3/c1 ;
 wire \V4/V3/V3/A2/M3/c2 ;
 wire \V4/V3/V3/A2/M3/s1 ;
 wire \V4/V3/V3/A2/M4/c1 ;
 wire \V4/V3/V3/A2/M4/c2 ;
 wire \V4/V3/V3/A2/M4/s1 ;
 wire \V4/V3/V3/A3/c1 ;
 wire \V4/V3/V3/A3/c2 ;
 wire \V4/V3/V3/A3/c3 ;
 wire \V4/V3/V3/A3/M1/c1 ;
 wire \V4/V3/V3/A3/M1/c2 ;
 wire \V4/V3/V3/A3/M1/s1 ;
 wire \V4/V3/V3/A3/M2/c1 ;
 wire \V4/V3/V3/A3/M2/c2 ;
 wire \V4/V3/V3/A3/M2/s1 ;
 wire \V4/V3/V3/A3/M3/c1 ;
 wire \V4/V3/V3/A3/M3/c2 ;
 wire \V4/V3/V3/A3/M3/s1 ;
 wire \V4/V3/V3/A3/M4/c1 ;
 wire \V4/V3/V3/A3/M4/c2 ;
 wire \V4/V3/V3/A3/M4/s1 ;
 wire \V4/V3/V3/V1/w1 ;
 wire \V4/V3/V3/V1/w2 ;
 wire \V4/V3/V3/V1/w3 ;
 wire \V4/V3/V3/V1/w4 ;
 wire \V4/V3/V3/V2/w1 ;
 wire \V4/V3/V3/V2/w2 ;
 wire \V4/V3/V3/V2/w3 ;
 wire \V4/V3/V3/V2/w4 ;
 wire \V4/V3/V3/V3/w1 ;
 wire \V4/V3/V3/V3/w2 ;
 wire \V4/V3/V3/V3/w3 ;
 wire \V4/V3/V3/V3/w4 ;
 wire \V4/V3/V3/V4/w1 ;
 wire \V4/V3/V3/V4/w2 ;
 wire \V4/V3/V3/V4/w3 ;
 wire \V4/V3/V3/V4/w4 ;
 wire \V4/V3/V4/c1 ;
 wire \V4/V3/V4/c2 ;
 wire \V4/V3/V4/c3 ;
 wire \V4/V3/V4/overflow ;
 wire \V4/V3/V4/A1/c1 ;
 wire \V4/V3/V4/A1/c2 ;
 wire \V4/V3/V4/A1/c3 ;
 wire \V4/V3/V4/A1/M1/c1 ;
 wire \V4/V3/V4/A1/M1/c2 ;
 wire \V4/V3/V4/A1/M1/s1 ;
 wire \V4/V3/V4/A1/M2/c1 ;
 wire \V4/V3/V4/A1/M2/c2 ;
 wire \V4/V3/V4/A1/M2/s1 ;
 wire \V4/V3/V4/A1/M3/c1 ;
 wire \V4/V3/V4/A1/M3/c2 ;
 wire \V4/V3/V4/A1/M3/s1 ;
 wire \V4/V3/V4/A1/M4/c1 ;
 wire \V4/V3/V4/A1/M4/c2 ;
 wire \V4/V3/V4/A1/M4/s1 ;
 wire \V4/V3/V4/A2/c1 ;
 wire \V4/V3/V4/A2/c2 ;
 wire \V4/V3/V4/A2/c3 ;
 wire \V4/V3/V4/A2/M1/c1 ;
 wire \V4/V3/V4/A2/M1/c2 ;
 wire \V4/V3/V4/A2/M1/s1 ;
 wire \V4/V3/V4/A2/M2/c1 ;
 wire \V4/V3/V4/A2/M2/c2 ;
 wire \V4/V3/V4/A2/M2/s1 ;
 wire \V4/V3/V4/A2/M3/c1 ;
 wire \V4/V3/V4/A2/M3/c2 ;
 wire \V4/V3/V4/A2/M3/s1 ;
 wire \V4/V3/V4/A2/M4/c1 ;
 wire \V4/V3/V4/A2/M4/c2 ;
 wire \V4/V3/V4/A2/M4/s1 ;
 wire \V4/V3/V4/A3/c1 ;
 wire \V4/V3/V4/A3/c2 ;
 wire \V4/V3/V4/A3/c3 ;
 wire \V4/V3/V4/A3/M1/c1 ;
 wire \V4/V3/V4/A3/M1/c2 ;
 wire \V4/V3/V4/A3/M1/s1 ;
 wire \V4/V3/V4/A3/M2/c1 ;
 wire \V4/V3/V4/A3/M2/c2 ;
 wire \V4/V3/V4/A3/M2/s1 ;
 wire \V4/V3/V4/A3/M3/c1 ;
 wire \V4/V3/V4/A3/M3/c2 ;
 wire \V4/V3/V4/A3/M3/s1 ;
 wire \V4/V3/V4/A3/M4/c1 ;
 wire \V4/V3/V4/A3/M4/c2 ;
 wire \V4/V3/V4/A3/M4/s1 ;
 wire \V4/V3/V4/V1/w1 ;
 wire \V4/V3/V4/V1/w2 ;
 wire \V4/V3/V4/V1/w3 ;
 wire \V4/V3/V4/V1/w4 ;
 wire \V4/V3/V4/V2/w1 ;
 wire \V4/V3/V4/V2/w2 ;
 wire \V4/V3/V4/V2/w3 ;
 wire \V4/V3/V4/V2/w4 ;
 wire \V4/V3/V4/V3/w1 ;
 wire \V4/V3/V4/V3/w2 ;
 wire \V4/V3/V4/V3/w3 ;
 wire \V4/V3/V4/V3/w4 ;
 wire \V4/V3/V4/V4/w1 ;
 wire \V4/V3/V4/V4/w2 ;
 wire \V4/V3/V4/V4/w3 ;
 wire \V4/V3/V4/V4/w4 ;
 wire \V4/V4/c1 ;
 wire \V4/V4/c2 ;
 wire \V4/V4/c3 ;
 wire \V4/V4/overflow ;
 wire \V4/V4/A1/c1 ;
 wire \V4/V4/A1/A1/c1 ;
 wire \V4/V4/A1/A1/c2 ;
 wire \V4/V4/A1/A1/c3 ;
 wire \V4/V4/A1/A1/M1/c1 ;
 wire \V4/V4/A1/A1/M1/c2 ;
 wire \V4/V4/A1/A1/M1/s1 ;
 wire \V4/V4/A1/A1/M2/c1 ;
 wire \V4/V4/A1/A1/M2/c2 ;
 wire \V4/V4/A1/A1/M2/s1 ;
 wire \V4/V4/A1/A1/M3/c1 ;
 wire \V4/V4/A1/A1/M3/c2 ;
 wire \V4/V4/A1/A1/M3/s1 ;
 wire \V4/V4/A1/A1/M4/c1 ;
 wire \V4/V4/A1/A1/M4/c2 ;
 wire \V4/V4/A1/A1/M4/s1 ;
 wire \V4/V4/A1/A2/c1 ;
 wire \V4/V4/A1/A2/c2 ;
 wire \V4/V4/A1/A2/c3 ;
 wire \V4/V4/A1/A2/M1/c1 ;
 wire \V4/V4/A1/A2/M1/c2 ;
 wire \V4/V4/A1/A2/M1/s1 ;
 wire \V4/V4/A1/A2/M2/c1 ;
 wire \V4/V4/A1/A2/M2/c2 ;
 wire \V4/V4/A1/A2/M2/s1 ;
 wire \V4/V4/A1/A2/M3/c1 ;
 wire \V4/V4/A1/A2/M3/c2 ;
 wire \V4/V4/A1/A2/M3/s1 ;
 wire \V4/V4/A1/A2/M4/c1 ;
 wire \V4/V4/A1/A2/M4/c2 ;
 wire \V4/V4/A1/A2/M4/s1 ;
 wire \V4/V4/A2/c1 ;
 wire \V4/V4/A2/A1/c1 ;
 wire \V4/V4/A2/A1/c2 ;
 wire \V4/V4/A2/A1/c3 ;
 wire \V4/V4/A2/A1/M1/c1 ;
 wire \V4/V4/A2/A1/M1/c2 ;
 wire \V4/V4/A2/A1/M1/s1 ;
 wire \V4/V4/A2/A1/M2/c1 ;
 wire \V4/V4/A2/A1/M2/c2 ;
 wire \V4/V4/A2/A1/M2/s1 ;
 wire \V4/V4/A2/A1/M3/c1 ;
 wire \V4/V4/A2/A1/M3/c2 ;
 wire \V4/V4/A2/A1/M3/s1 ;
 wire \V4/V4/A2/A1/M4/c1 ;
 wire \V4/V4/A2/A1/M4/c2 ;
 wire \V4/V4/A2/A1/M4/s1 ;
 wire \V4/V4/A2/A2/c1 ;
 wire \V4/V4/A2/A2/c2 ;
 wire \V4/V4/A2/A2/c3 ;
 wire \V4/V4/A2/A2/M1/c1 ;
 wire \V4/V4/A2/A2/M1/c2 ;
 wire \V4/V4/A2/A2/M1/s1 ;
 wire \V4/V4/A2/A2/M2/c1 ;
 wire \V4/V4/A2/A2/M2/c2 ;
 wire \V4/V4/A2/A2/M2/s1 ;
 wire \V4/V4/A2/A2/M3/c1 ;
 wire \V4/V4/A2/A2/M3/c2 ;
 wire \V4/V4/A2/A2/M3/s1 ;
 wire \V4/V4/A2/A2/M4/c1 ;
 wire \V4/V4/A2/A2/M4/c2 ;
 wire \V4/V4/A2/A2/M4/s1 ;
 wire \V4/V4/A3/c1 ;
 wire \V4/V4/A3/A1/c1 ;
 wire \V4/V4/A3/A1/c2 ;
 wire \V4/V4/A3/A1/c3 ;
 wire \V4/V4/A3/A1/M1/c1 ;
 wire \V4/V4/A3/A1/M1/c2 ;
 wire \V4/V4/A3/A1/M1/s1 ;
 wire \V4/V4/A3/A1/M2/c1 ;
 wire \V4/V4/A3/A1/M2/c2 ;
 wire \V4/V4/A3/A1/M2/s1 ;
 wire \V4/V4/A3/A1/M3/c1 ;
 wire \V4/V4/A3/A1/M3/c2 ;
 wire \V4/V4/A3/A1/M3/s1 ;
 wire \V4/V4/A3/A1/M4/c1 ;
 wire \V4/V4/A3/A1/M4/c2 ;
 wire \V4/V4/A3/A1/M4/s1 ;
 wire \V4/V4/A3/A2/c1 ;
 wire \V4/V4/A3/A2/c2 ;
 wire \V4/V4/A3/A2/c3 ;
 wire \V4/V4/A3/A2/M1/c1 ;
 wire \V4/V4/A3/A2/M1/c2 ;
 wire \V4/V4/A3/A2/M1/s1 ;
 wire \V4/V4/A3/A2/M2/c1 ;
 wire \V4/V4/A3/A2/M2/c2 ;
 wire \V4/V4/A3/A2/M2/s1 ;
 wire \V4/V4/A3/A2/M3/c1 ;
 wire \V4/V4/A3/A2/M3/c2 ;
 wire \V4/V4/A3/A2/M3/s1 ;
 wire \V4/V4/A3/A2/M4/c1 ;
 wire \V4/V4/A3/A2/M4/c2 ;
 wire \V4/V4/A3/A2/M4/s1 ;
 wire \V4/V4/V1/c1 ;
 wire \V4/V4/V1/c2 ;
 wire \V4/V4/V1/c3 ;
 wire \V4/V4/V1/overflow ;
 wire \V4/V4/V1/A1/c1 ;
 wire \V4/V4/V1/A1/c2 ;
 wire \V4/V4/V1/A1/c3 ;
 wire \V4/V4/V1/A1/M1/c1 ;
 wire \V4/V4/V1/A1/M1/c2 ;
 wire \V4/V4/V1/A1/M1/s1 ;
 wire \V4/V4/V1/A1/M2/c1 ;
 wire \V4/V4/V1/A1/M2/c2 ;
 wire \V4/V4/V1/A1/M2/s1 ;
 wire \V4/V4/V1/A1/M3/c1 ;
 wire \V4/V4/V1/A1/M3/c2 ;
 wire \V4/V4/V1/A1/M3/s1 ;
 wire \V4/V4/V1/A1/M4/c1 ;
 wire \V4/V4/V1/A1/M4/c2 ;
 wire \V4/V4/V1/A1/M4/s1 ;
 wire \V4/V4/V1/A2/c1 ;
 wire \V4/V4/V1/A2/c2 ;
 wire \V4/V4/V1/A2/c3 ;
 wire \V4/V4/V1/A2/M1/c1 ;
 wire \V4/V4/V1/A2/M1/c2 ;
 wire \V4/V4/V1/A2/M1/s1 ;
 wire \V4/V4/V1/A2/M2/c1 ;
 wire \V4/V4/V1/A2/M2/c2 ;
 wire \V4/V4/V1/A2/M2/s1 ;
 wire \V4/V4/V1/A2/M3/c1 ;
 wire \V4/V4/V1/A2/M3/c2 ;
 wire \V4/V4/V1/A2/M3/s1 ;
 wire \V4/V4/V1/A2/M4/c1 ;
 wire \V4/V4/V1/A2/M4/c2 ;
 wire \V4/V4/V1/A2/M4/s1 ;
 wire \V4/V4/V1/A3/c1 ;
 wire \V4/V4/V1/A3/c2 ;
 wire \V4/V4/V1/A3/c3 ;
 wire \V4/V4/V1/A3/M1/c1 ;
 wire \V4/V4/V1/A3/M1/c2 ;
 wire \V4/V4/V1/A3/M1/s1 ;
 wire \V4/V4/V1/A3/M2/c1 ;
 wire \V4/V4/V1/A3/M2/c2 ;
 wire \V4/V4/V1/A3/M2/s1 ;
 wire \V4/V4/V1/A3/M3/c1 ;
 wire \V4/V4/V1/A3/M3/c2 ;
 wire \V4/V4/V1/A3/M3/s1 ;
 wire \V4/V4/V1/A3/M4/c1 ;
 wire \V4/V4/V1/A3/M4/c2 ;
 wire \V4/V4/V1/A3/M4/s1 ;
 wire \V4/V4/V1/V1/w1 ;
 wire \V4/V4/V1/V1/w2 ;
 wire \V4/V4/V1/V1/w3 ;
 wire \V4/V4/V1/V1/w4 ;
 wire \V4/V4/V1/V2/w1 ;
 wire \V4/V4/V1/V2/w2 ;
 wire \V4/V4/V1/V2/w3 ;
 wire \V4/V4/V1/V2/w4 ;
 wire \V4/V4/V1/V3/w1 ;
 wire \V4/V4/V1/V3/w2 ;
 wire \V4/V4/V1/V3/w3 ;
 wire \V4/V4/V1/V3/w4 ;
 wire \V4/V4/V1/V4/w1 ;
 wire \V4/V4/V1/V4/w2 ;
 wire \V4/V4/V1/V4/w3 ;
 wire \V4/V4/V1/V4/w4 ;
 wire \V4/V4/V2/c1 ;
 wire \V4/V4/V2/c2 ;
 wire \V4/V4/V2/c3 ;
 wire \V4/V4/V2/overflow ;
 wire \V4/V4/V2/A1/c1 ;
 wire \V4/V4/V2/A1/c2 ;
 wire \V4/V4/V2/A1/c3 ;
 wire \V4/V4/V2/A1/M1/c1 ;
 wire \V4/V4/V2/A1/M1/c2 ;
 wire \V4/V4/V2/A1/M1/s1 ;
 wire \V4/V4/V2/A1/M2/c1 ;
 wire \V4/V4/V2/A1/M2/c2 ;
 wire \V4/V4/V2/A1/M2/s1 ;
 wire \V4/V4/V2/A1/M3/c1 ;
 wire \V4/V4/V2/A1/M3/c2 ;
 wire \V4/V4/V2/A1/M3/s1 ;
 wire \V4/V4/V2/A1/M4/c1 ;
 wire \V4/V4/V2/A1/M4/c2 ;
 wire \V4/V4/V2/A1/M4/s1 ;
 wire \V4/V4/V2/A2/c1 ;
 wire \V4/V4/V2/A2/c2 ;
 wire \V4/V4/V2/A2/c3 ;
 wire \V4/V4/V2/A2/M1/c1 ;
 wire \V4/V4/V2/A2/M1/c2 ;
 wire \V4/V4/V2/A2/M1/s1 ;
 wire \V4/V4/V2/A2/M2/c1 ;
 wire \V4/V4/V2/A2/M2/c2 ;
 wire \V4/V4/V2/A2/M2/s1 ;
 wire \V4/V4/V2/A2/M3/c1 ;
 wire \V4/V4/V2/A2/M3/c2 ;
 wire \V4/V4/V2/A2/M3/s1 ;
 wire \V4/V4/V2/A2/M4/c1 ;
 wire \V4/V4/V2/A2/M4/c2 ;
 wire \V4/V4/V2/A2/M4/s1 ;
 wire \V4/V4/V2/A3/c1 ;
 wire \V4/V4/V2/A3/c2 ;
 wire \V4/V4/V2/A3/c3 ;
 wire \V4/V4/V2/A3/M1/c1 ;
 wire \V4/V4/V2/A3/M1/c2 ;
 wire \V4/V4/V2/A3/M1/s1 ;
 wire \V4/V4/V2/A3/M2/c1 ;
 wire \V4/V4/V2/A3/M2/c2 ;
 wire \V4/V4/V2/A3/M2/s1 ;
 wire \V4/V4/V2/A3/M3/c1 ;
 wire \V4/V4/V2/A3/M3/c2 ;
 wire \V4/V4/V2/A3/M3/s1 ;
 wire \V4/V4/V2/A3/M4/c1 ;
 wire \V4/V4/V2/A3/M4/c2 ;
 wire \V4/V4/V2/A3/M4/s1 ;
 wire \V4/V4/V2/V1/w1 ;
 wire \V4/V4/V2/V1/w2 ;
 wire \V4/V4/V2/V1/w3 ;
 wire \V4/V4/V2/V1/w4 ;
 wire \V4/V4/V2/V2/w1 ;
 wire \V4/V4/V2/V2/w2 ;
 wire \V4/V4/V2/V2/w3 ;
 wire \V4/V4/V2/V2/w4 ;
 wire \V4/V4/V2/V3/w1 ;
 wire \V4/V4/V2/V3/w2 ;
 wire \V4/V4/V2/V3/w3 ;
 wire \V4/V4/V2/V3/w4 ;
 wire \V4/V4/V2/V4/w1 ;
 wire \V4/V4/V2/V4/w2 ;
 wire \V4/V4/V2/V4/w3 ;
 wire \V4/V4/V2/V4/w4 ;
 wire \V4/V4/V3/c1 ;
 wire \V4/V4/V3/c2 ;
 wire \V4/V4/V3/c3 ;
 wire \V4/V4/V3/overflow ;
 wire \V4/V4/V3/A1/c1 ;
 wire \V4/V4/V3/A1/c2 ;
 wire \V4/V4/V3/A1/c3 ;
 wire \V4/V4/V3/A1/M1/c1 ;
 wire \V4/V4/V3/A1/M1/c2 ;
 wire \V4/V4/V3/A1/M1/s1 ;
 wire \V4/V4/V3/A1/M2/c1 ;
 wire \V4/V4/V3/A1/M2/c2 ;
 wire \V4/V4/V3/A1/M2/s1 ;
 wire \V4/V4/V3/A1/M3/c1 ;
 wire \V4/V4/V3/A1/M3/c2 ;
 wire \V4/V4/V3/A1/M3/s1 ;
 wire \V4/V4/V3/A1/M4/c1 ;
 wire \V4/V4/V3/A1/M4/c2 ;
 wire \V4/V4/V3/A1/M4/s1 ;
 wire \V4/V4/V3/A2/c1 ;
 wire \V4/V4/V3/A2/c2 ;
 wire \V4/V4/V3/A2/c3 ;
 wire \V4/V4/V3/A2/M1/c1 ;
 wire \V4/V4/V3/A2/M1/c2 ;
 wire \V4/V4/V3/A2/M1/s1 ;
 wire \V4/V4/V3/A2/M2/c1 ;
 wire \V4/V4/V3/A2/M2/c2 ;
 wire \V4/V4/V3/A2/M2/s1 ;
 wire \V4/V4/V3/A2/M3/c1 ;
 wire \V4/V4/V3/A2/M3/c2 ;
 wire \V4/V4/V3/A2/M3/s1 ;
 wire \V4/V4/V3/A2/M4/c1 ;
 wire \V4/V4/V3/A2/M4/c2 ;
 wire \V4/V4/V3/A2/M4/s1 ;
 wire \V4/V4/V3/A3/c1 ;
 wire \V4/V4/V3/A3/c2 ;
 wire \V4/V4/V3/A3/c3 ;
 wire \V4/V4/V3/A3/M1/c1 ;
 wire \V4/V4/V3/A3/M1/c2 ;
 wire \V4/V4/V3/A3/M1/s1 ;
 wire \V4/V4/V3/A3/M2/c1 ;
 wire \V4/V4/V3/A3/M2/c2 ;
 wire \V4/V4/V3/A3/M2/s1 ;
 wire \V4/V4/V3/A3/M3/c1 ;
 wire \V4/V4/V3/A3/M3/c2 ;
 wire \V4/V4/V3/A3/M3/s1 ;
 wire \V4/V4/V3/A3/M4/c1 ;
 wire \V4/V4/V3/A3/M4/c2 ;
 wire \V4/V4/V3/A3/M4/s1 ;
 wire \V4/V4/V3/V1/w1 ;
 wire \V4/V4/V3/V1/w2 ;
 wire \V4/V4/V3/V1/w3 ;
 wire \V4/V4/V3/V1/w4 ;
 wire \V4/V4/V3/V2/w1 ;
 wire \V4/V4/V3/V2/w2 ;
 wire \V4/V4/V3/V2/w3 ;
 wire \V4/V4/V3/V2/w4 ;
 wire \V4/V4/V3/V3/w1 ;
 wire \V4/V4/V3/V3/w2 ;
 wire \V4/V4/V3/V3/w3 ;
 wire \V4/V4/V3/V3/w4 ;
 wire \V4/V4/V3/V4/w1 ;
 wire \V4/V4/V3/V4/w2 ;
 wire \V4/V4/V3/V4/w3 ;
 wire \V4/V4/V3/V4/w4 ;
 wire \V4/V4/V4/c1 ;
 wire \V4/V4/V4/c2 ;
 wire \V4/V4/V4/c3 ;
 wire \V4/V4/V4/overflow ;
 wire \V4/V4/V4/A1/c1 ;
 wire \V4/V4/V4/A1/c2 ;
 wire \V4/V4/V4/A1/c3 ;
 wire \V4/V4/V4/A1/M1/c1 ;
 wire \V4/V4/V4/A1/M1/c2 ;
 wire \V4/V4/V4/A1/M1/s1 ;
 wire \V4/V4/V4/A1/M2/c1 ;
 wire \V4/V4/V4/A1/M2/c2 ;
 wire \V4/V4/V4/A1/M2/s1 ;
 wire \V4/V4/V4/A1/M3/c1 ;
 wire \V4/V4/V4/A1/M3/c2 ;
 wire \V4/V4/V4/A1/M3/s1 ;
 wire \V4/V4/V4/A1/M4/c1 ;
 wire \V4/V4/V4/A1/M4/c2 ;
 wire \V4/V4/V4/A1/M4/s1 ;
 wire \V4/V4/V4/A2/c1 ;
 wire \V4/V4/V4/A2/c2 ;
 wire \V4/V4/V4/A2/c3 ;
 wire \V4/V4/V4/A2/M1/c1 ;
 wire \V4/V4/V4/A2/M1/c2 ;
 wire \V4/V4/V4/A2/M1/s1 ;
 wire \V4/V4/V4/A2/M2/c1 ;
 wire \V4/V4/V4/A2/M2/c2 ;
 wire \V4/V4/V4/A2/M2/s1 ;
 wire \V4/V4/V4/A2/M3/c1 ;
 wire \V4/V4/V4/A2/M3/c2 ;
 wire \V4/V4/V4/A2/M3/s1 ;
 wire \V4/V4/V4/A2/M4/c1 ;
 wire \V4/V4/V4/A2/M4/c2 ;
 wire \V4/V4/V4/A2/M4/s1 ;
 wire \V4/V4/V4/A3/c1 ;
 wire \V4/V4/V4/A3/c2 ;
 wire \V4/V4/V4/A3/c3 ;
 wire \V4/V4/V4/A3/M1/c1 ;
 wire \V4/V4/V4/A3/M1/c2 ;
 wire \V4/V4/V4/A3/M1/s1 ;
 wire \V4/V4/V4/A3/M2/c1 ;
 wire \V4/V4/V4/A3/M2/c2 ;
 wire \V4/V4/V4/A3/M2/s1 ;
 wire \V4/V4/V4/A3/M3/c1 ;
 wire \V4/V4/V4/A3/M3/c2 ;
 wire \V4/V4/V4/A3/M3/s1 ;
 wire \V4/V4/V4/A3/M4/c1 ;
 wire \V4/V4/V4/A3/M4/c2 ;
 wire \V4/V4/V4/A3/M4/s1 ;
 wire \V4/V4/V4/V1/w1 ;
 wire \V4/V4/V4/V1/w2 ;
 wire \V4/V4/V4/V1/w3 ;
 wire \V4/V4/V4/V1/w4 ;
 wire \V4/V4/V4/V2/w1 ;
 wire \V4/V4/V4/V2/w2 ;
 wire \V4/V4/V4/V2/w3 ;
 wire \V4/V4/V4/V2/w4 ;
 wire \V4/V4/V4/V3/w1 ;
 wire \V4/V4/V4/V3/w2 ;
 wire \V4/V4/V4/V3/w3 ;
 wire \V4/V4/V4/V3/w4 ;
 wire \V4/V4/V4/V4/w1 ;
 wire \V4/V4/V4/V4/w2 ;
 wire \V4/V4/V4/V4/w3 ;
 wire \V4/V4/V4/V4/w4 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire [3:0] \V1/V1/V1/s1 ;
 wire [3:0] \V1/V1/V1/s2 ;
 wire [3:0] \V1/V1/V1/v1 ;
 wire [3:0] \V1/V1/V1/v2 ;
 wire [3:0] \V1/V1/V1/v3 ;
 wire [3:0] \V1/V1/V1/v4 ;
 wire [3:0] \V1/V1/V2/s1 ;
 wire [3:0] \V1/V1/V2/s2 ;
 wire [3:0] \V1/V1/V2/v1 ;
 wire [3:0] \V1/V1/V2/v2 ;
 wire [3:0] \V1/V1/V2/v3 ;
 wire [3:0] \V1/V1/V2/v4 ;
 wire [3:0] \V1/V1/V3/s1 ;
 wire [3:0] \V1/V1/V3/s2 ;
 wire [3:0] \V1/V1/V3/v1 ;
 wire [3:0] \V1/V1/V3/v2 ;
 wire [3:0] \V1/V1/V3/v3 ;
 wire [3:0] \V1/V1/V3/v4 ;
 wire [3:0] \V1/V1/V4/s1 ;
 wire [3:0] \V1/V1/V4/s2 ;
 wire [3:0] \V1/V1/V4/v1 ;
 wire [3:0] \V1/V1/V4/v2 ;
 wire [3:0] \V1/V1/V4/v3 ;
 wire [3:0] \V1/V1/V4/v4 ;
 wire [7:0] \V1/V1/s1 ;
 wire [7:0] \V1/V1/s2 ;
 wire [7:0] \V1/V1/v1 ;
 wire [7:0] \V1/V1/v2 ;
 wire [7:0] \V1/V1/v3 ;
 wire [7:0] \V1/V1/v4 ;
 wire [3:0] \V1/V2/V1/s1 ;
 wire [3:0] \V1/V2/V1/s2 ;
 wire [3:0] \V1/V2/V1/v1 ;
 wire [3:0] \V1/V2/V1/v2 ;
 wire [3:0] \V1/V2/V1/v3 ;
 wire [3:0] \V1/V2/V1/v4 ;
 wire [3:0] \V1/V2/V2/s1 ;
 wire [3:0] \V1/V2/V2/s2 ;
 wire [3:0] \V1/V2/V2/v1 ;
 wire [3:0] \V1/V2/V2/v2 ;
 wire [3:0] \V1/V2/V2/v3 ;
 wire [3:0] \V1/V2/V2/v4 ;
 wire [3:0] \V1/V2/V3/s1 ;
 wire [3:0] \V1/V2/V3/s2 ;
 wire [3:0] \V1/V2/V3/v1 ;
 wire [3:0] \V1/V2/V3/v2 ;
 wire [3:0] \V1/V2/V3/v3 ;
 wire [3:0] \V1/V2/V3/v4 ;
 wire [3:0] \V1/V2/V4/s1 ;
 wire [3:0] \V1/V2/V4/s2 ;
 wire [3:0] \V1/V2/V4/v1 ;
 wire [3:0] \V1/V2/V4/v2 ;
 wire [3:0] \V1/V2/V4/v3 ;
 wire [3:0] \V1/V2/V4/v4 ;
 wire [7:0] \V1/V2/s1 ;
 wire [7:0] \V1/V2/s2 ;
 wire [7:0] \V1/V2/v1 ;
 wire [7:0] \V1/V2/v2 ;
 wire [7:0] \V1/V2/v3 ;
 wire [7:0] \V1/V2/v4 ;
 wire [3:0] \V1/V3/V1/s1 ;
 wire [3:0] \V1/V3/V1/s2 ;
 wire [3:0] \V1/V3/V1/v1 ;
 wire [3:0] \V1/V3/V1/v2 ;
 wire [3:0] \V1/V3/V1/v3 ;
 wire [3:0] \V1/V3/V1/v4 ;
 wire [3:0] \V1/V3/V2/s1 ;
 wire [3:0] \V1/V3/V2/s2 ;
 wire [3:0] \V1/V3/V2/v1 ;
 wire [3:0] \V1/V3/V2/v2 ;
 wire [3:0] \V1/V3/V2/v3 ;
 wire [3:0] \V1/V3/V2/v4 ;
 wire [3:0] \V1/V3/V3/s1 ;
 wire [3:0] \V1/V3/V3/s2 ;
 wire [3:0] \V1/V3/V3/v1 ;
 wire [3:0] \V1/V3/V3/v2 ;
 wire [3:0] \V1/V3/V3/v3 ;
 wire [3:0] \V1/V3/V3/v4 ;
 wire [3:0] \V1/V3/V4/s1 ;
 wire [3:0] \V1/V3/V4/s2 ;
 wire [3:0] \V1/V3/V4/v1 ;
 wire [3:0] \V1/V3/V4/v2 ;
 wire [3:0] \V1/V3/V4/v3 ;
 wire [3:0] \V1/V3/V4/v4 ;
 wire [7:0] \V1/V3/s1 ;
 wire [7:0] \V1/V3/s2 ;
 wire [7:0] \V1/V3/v1 ;
 wire [7:0] \V1/V3/v2 ;
 wire [7:0] \V1/V3/v3 ;
 wire [7:0] \V1/V3/v4 ;
 wire [3:0] \V1/V4/V1/s1 ;
 wire [3:0] \V1/V4/V1/s2 ;
 wire [3:0] \V1/V4/V1/v1 ;
 wire [3:0] \V1/V4/V1/v2 ;
 wire [3:0] \V1/V4/V1/v3 ;
 wire [3:0] \V1/V4/V1/v4 ;
 wire [3:0] \V1/V4/V2/s1 ;
 wire [3:0] \V1/V4/V2/s2 ;
 wire [3:0] \V1/V4/V2/v1 ;
 wire [3:0] \V1/V4/V2/v2 ;
 wire [3:0] \V1/V4/V2/v3 ;
 wire [3:0] \V1/V4/V2/v4 ;
 wire [3:0] \V1/V4/V3/s1 ;
 wire [3:0] \V1/V4/V3/s2 ;
 wire [3:0] \V1/V4/V3/v1 ;
 wire [3:0] \V1/V4/V3/v2 ;
 wire [3:0] \V1/V4/V3/v3 ;
 wire [3:0] \V1/V4/V3/v4 ;
 wire [3:0] \V1/V4/V4/s1 ;
 wire [3:0] \V1/V4/V4/s2 ;
 wire [3:0] \V1/V4/V4/v1 ;
 wire [3:0] \V1/V4/V4/v2 ;
 wire [3:0] \V1/V4/V4/v3 ;
 wire [3:0] \V1/V4/V4/v4 ;
 wire [7:0] \V1/V4/s1 ;
 wire [7:0] \V1/V4/s2 ;
 wire [7:0] \V1/V4/v1 ;
 wire [7:0] \V1/V4/v2 ;
 wire [7:0] \V1/V4/v3 ;
 wire [7:0] \V1/V4/v4 ;
 wire [15:0] \V1/s1 ;
 wire [15:0] \V1/s2 ;
 wire [15:0] \V1/v1 ;
 wire [15:0] \V1/v2 ;
 wire [15:0] \V1/v3 ;
 wire [15:0] \V1/v4 ;
 wire [3:0] \V2/V1/V1/s1 ;
 wire [3:0] \V2/V1/V1/s2 ;
 wire [3:0] \V2/V1/V1/v1 ;
 wire [3:0] \V2/V1/V1/v2 ;
 wire [3:0] \V2/V1/V1/v3 ;
 wire [3:0] \V2/V1/V1/v4 ;
 wire [3:0] \V2/V1/V2/s1 ;
 wire [3:0] \V2/V1/V2/s2 ;
 wire [3:0] \V2/V1/V2/v1 ;
 wire [3:0] \V2/V1/V2/v2 ;
 wire [3:0] \V2/V1/V2/v3 ;
 wire [3:0] \V2/V1/V2/v4 ;
 wire [3:0] \V2/V1/V3/s1 ;
 wire [3:0] \V2/V1/V3/s2 ;
 wire [3:0] \V2/V1/V3/v1 ;
 wire [3:0] \V2/V1/V3/v2 ;
 wire [3:0] \V2/V1/V3/v3 ;
 wire [3:0] \V2/V1/V3/v4 ;
 wire [3:0] \V2/V1/V4/s1 ;
 wire [3:0] \V2/V1/V4/s2 ;
 wire [3:0] \V2/V1/V4/v1 ;
 wire [3:0] \V2/V1/V4/v2 ;
 wire [3:0] \V2/V1/V4/v3 ;
 wire [3:0] \V2/V1/V4/v4 ;
 wire [7:0] \V2/V1/s1 ;
 wire [7:0] \V2/V1/s2 ;
 wire [7:0] \V2/V1/v1 ;
 wire [7:0] \V2/V1/v2 ;
 wire [7:0] \V2/V1/v3 ;
 wire [7:0] \V2/V1/v4 ;
 wire [3:0] \V2/V2/V1/s1 ;
 wire [3:0] \V2/V2/V1/s2 ;
 wire [3:0] \V2/V2/V1/v1 ;
 wire [3:0] \V2/V2/V1/v2 ;
 wire [3:0] \V2/V2/V1/v3 ;
 wire [3:0] \V2/V2/V1/v4 ;
 wire [3:0] \V2/V2/V2/s1 ;
 wire [3:0] \V2/V2/V2/s2 ;
 wire [3:0] \V2/V2/V2/v1 ;
 wire [3:0] \V2/V2/V2/v2 ;
 wire [3:0] \V2/V2/V2/v3 ;
 wire [3:0] \V2/V2/V2/v4 ;
 wire [3:0] \V2/V2/V3/s1 ;
 wire [3:0] \V2/V2/V3/s2 ;
 wire [3:0] \V2/V2/V3/v1 ;
 wire [3:0] \V2/V2/V3/v2 ;
 wire [3:0] \V2/V2/V3/v3 ;
 wire [3:0] \V2/V2/V3/v4 ;
 wire [3:0] \V2/V2/V4/s1 ;
 wire [3:0] \V2/V2/V4/s2 ;
 wire [3:0] \V2/V2/V4/v1 ;
 wire [3:0] \V2/V2/V4/v2 ;
 wire [3:0] \V2/V2/V4/v3 ;
 wire [3:0] \V2/V2/V4/v4 ;
 wire [7:0] \V2/V2/s1 ;
 wire [7:0] \V2/V2/s2 ;
 wire [7:0] \V2/V2/v1 ;
 wire [7:0] \V2/V2/v2 ;
 wire [7:0] \V2/V2/v3 ;
 wire [7:0] \V2/V2/v4 ;
 wire [3:0] \V2/V3/V1/s1 ;
 wire [3:0] \V2/V3/V1/s2 ;
 wire [3:0] \V2/V3/V1/v1 ;
 wire [3:0] \V2/V3/V1/v2 ;
 wire [3:0] \V2/V3/V1/v3 ;
 wire [3:0] \V2/V3/V1/v4 ;
 wire [3:0] \V2/V3/V2/s1 ;
 wire [3:0] \V2/V3/V2/s2 ;
 wire [3:0] \V2/V3/V2/v1 ;
 wire [3:0] \V2/V3/V2/v2 ;
 wire [3:0] \V2/V3/V2/v3 ;
 wire [3:0] \V2/V3/V2/v4 ;
 wire [3:0] \V2/V3/V3/s1 ;
 wire [3:0] \V2/V3/V3/s2 ;
 wire [3:0] \V2/V3/V3/v1 ;
 wire [3:0] \V2/V3/V3/v2 ;
 wire [3:0] \V2/V3/V3/v3 ;
 wire [3:0] \V2/V3/V3/v4 ;
 wire [3:0] \V2/V3/V4/s1 ;
 wire [3:0] \V2/V3/V4/s2 ;
 wire [3:0] \V2/V3/V4/v1 ;
 wire [3:0] \V2/V3/V4/v2 ;
 wire [3:0] \V2/V3/V4/v3 ;
 wire [3:0] \V2/V3/V4/v4 ;
 wire [7:0] \V2/V3/s1 ;
 wire [7:0] \V2/V3/s2 ;
 wire [7:0] \V2/V3/v1 ;
 wire [7:0] \V2/V3/v2 ;
 wire [7:0] \V2/V3/v3 ;
 wire [7:0] \V2/V3/v4 ;
 wire [3:0] \V2/V4/V1/s1 ;
 wire [3:0] \V2/V4/V1/s2 ;
 wire [3:0] \V2/V4/V1/v1 ;
 wire [3:0] \V2/V4/V1/v2 ;
 wire [3:0] \V2/V4/V1/v3 ;
 wire [3:0] \V2/V4/V1/v4 ;
 wire [3:0] \V2/V4/V2/s1 ;
 wire [3:0] \V2/V4/V2/s2 ;
 wire [3:0] \V2/V4/V2/v1 ;
 wire [3:0] \V2/V4/V2/v2 ;
 wire [3:0] \V2/V4/V2/v3 ;
 wire [3:0] \V2/V4/V2/v4 ;
 wire [3:0] \V2/V4/V3/s1 ;
 wire [3:0] \V2/V4/V3/s2 ;
 wire [3:0] \V2/V4/V3/v1 ;
 wire [3:0] \V2/V4/V3/v2 ;
 wire [3:0] \V2/V4/V3/v3 ;
 wire [3:0] \V2/V4/V3/v4 ;
 wire [3:0] \V2/V4/V4/s1 ;
 wire [3:0] \V2/V4/V4/s2 ;
 wire [3:0] \V2/V4/V4/v1 ;
 wire [3:0] \V2/V4/V4/v2 ;
 wire [3:0] \V2/V4/V4/v3 ;
 wire [3:0] \V2/V4/V4/v4 ;
 wire [7:0] \V2/V4/s1 ;
 wire [7:0] \V2/V4/s2 ;
 wire [7:0] \V2/V4/v1 ;
 wire [7:0] \V2/V4/v2 ;
 wire [7:0] \V2/V4/v3 ;
 wire [7:0] \V2/V4/v4 ;
 wire [15:0] \V2/s1 ;
 wire [15:0] \V2/s2 ;
 wire [15:0] \V2/v1 ;
 wire [15:0] \V2/v2 ;
 wire [15:0] \V2/v3 ;
 wire [15:0] \V2/v4 ;
 wire [3:0] \V3/V1/V1/s1 ;
 wire [3:0] \V3/V1/V1/s2 ;
 wire [3:0] \V3/V1/V1/v1 ;
 wire [3:0] \V3/V1/V1/v2 ;
 wire [3:0] \V3/V1/V1/v3 ;
 wire [3:0] \V3/V1/V1/v4 ;
 wire [3:0] \V3/V1/V2/s1 ;
 wire [3:0] \V3/V1/V2/s2 ;
 wire [3:0] \V3/V1/V2/v1 ;
 wire [3:0] \V3/V1/V2/v2 ;
 wire [3:0] \V3/V1/V2/v3 ;
 wire [3:0] \V3/V1/V2/v4 ;
 wire [3:0] \V3/V1/V3/s1 ;
 wire [3:0] \V3/V1/V3/s2 ;
 wire [3:0] \V3/V1/V3/v1 ;
 wire [3:0] \V3/V1/V3/v2 ;
 wire [3:0] \V3/V1/V3/v3 ;
 wire [3:0] \V3/V1/V3/v4 ;
 wire [3:0] \V3/V1/V4/s1 ;
 wire [3:0] \V3/V1/V4/s2 ;
 wire [3:0] \V3/V1/V4/v1 ;
 wire [3:0] \V3/V1/V4/v2 ;
 wire [3:0] \V3/V1/V4/v3 ;
 wire [3:0] \V3/V1/V4/v4 ;
 wire [7:0] \V3/V1/s1 ;
 wire [7:0] \V3/V1/s2 ;
 wire [7:0] \V3/V1/v1 ;
 wire [7:0] \V3/V1/v2 ;
 wire [7:0] \V3/V1/v3 ;
 wire [7:0] \V3/V1/v4 ;
 wire [3:0] \V3/V2/V1/s1 ;
 wire [3:0] \V3/V2/V1/s2 ;
 wire [3:0] \V3/V2/V1/v1 ;
 wire [3:0] \V3/V2/V1/v2 ;
 wire [3:0] \V3/V2/V1/v3 ;
 wire [3:0] \V3/V2/V1/v4 ;
 wire [3:0] \V3/V2/V2/s1 ;
 wire [3:0] \V3/V2/V2/s2 ;
 wire [3:0] \V3/V2/V2/v1 ;
 wire [3:0] \V3/V2/V2/v2 ;
 wire [3:0] \V3/V2/V2/v3 ;
 wire [3:0] \V3/V2/V2/v4 ;
 wire [3:0] \V3/V2/V3/s1 ;
 wire [3:0] \V3/V2/V3/s2 ;
 wire [3:0] \V3/V2/V3/v1 ;
 wire [3:0] \V3/V2/V3/v2 ;
 wire [3:0] \V3/V2/V3/v3 ;
 wire [3:0] \V3/V2/V3/v4 ;
 wire [3:0] \V3/V2/V4/s1 ;
 wire [3:0] \V3/V2/V4/s2 ;
 wire [3:0] \V3/V2/V4/v1 ;
 wire [3:0] \V3/V2/V4/v2 ;
 wire [3:0] \V3/V2/V4/v3 ;
 wire [3:0] \V3/V2/V4/v4 ;
 wire [7:0] \V3/V2/s1 ;
 wire [7:0] \V3/V2/s2 ;
 wire [7:0] \V3/V2/v1 ;
 wire [7:0] \V3/V2/v2 ;
 wire [7:0] \V3/V2/v3 ;
 wire [7:0] \V3/V2/v4 ;
 wire [3:0] \V3/V3/V1/s1 ;
 wire [3:0] \V3/V3/V1/s2 ;
 wire [3:0] \V3/V3/V1/v1 ;
 wire [3:0] \V3/V3/V1/v2 ;
 wire [3:0] \V3/V3/V1/v3 ;
 wire [3:0] \V3/V3/V1/v4 ;
 wire [3:0] \V3/V3/V2/s1 ;
 wire [3:0] \V3/V3/V2/s2 ;
 wire [3:0] \V3/V3/V2/v1 ;
 wire [3:0] \V3/V3/V2/v2 ;
 wire [3:0] \V3/V3/V2/v3 ;
 wire [3:0] \V3/V3/V2/v4 ;
 wire [3:0] \V3/V3/V3/s1 ;
 wire [3:0] \V3/V3/V3/s2 ;
 wire [3:0] \V3/V3/V3/v1 ;
 wire [3:0] \V3/V3/V3/v2 ;
 wire [3:0] \V3/V3/V3/v3 ;
 wire [3:0] \V3/V3/V3/v4 ;
 wire [3:0] \V3/V3/V4/s1 ;
 wire [3:0] \V3/V3/V4/s2 ;
 wire [3:0] \V3/V3/V4/v1 ;
 wire [3:0] \V3/V3/V4/v2 ;
 wire [3:0] \V3/V3/V4/v3 ;
 wire [3:0] \V3/V3/V4/v4 ;
 wire [7:0] \V3/V3/s1 ;
 wire [7:0] \V3/V3/s2 ;
 wire [7:0] \V3/V3/v1 ;
 wire [7:0] \V3/V3/v2 ;
 wire [7:0] \V3/V3/v3 ;
 wire [7:0] \V3/V3/v4 ;
 wire [3:0] \V3/V4/V1/s1 ;
 wire [3:0] \V3/V4/V1/s2 ;
 wire [3:0] \V3/V4/V1/v1 ;
 wire [3:0] \V3/V4/V1/v2 ;
 wire [3:0] \V3/V4/V1/v3 ;
 wire [3:0] \V3/V4/V1/v4 ;
 wire [3:0] \V3/V4/V2/s1 ;
 wire [3:0] \V3/V4/V2/s2 ;
 wire [3:0] \V3/V4/V2/v1 ;
 wire [3:0] \V3/V4/V2/v2 ;
 wire [3:0] \V3/V4/V2/v3 ;
 wire [3:0] \V3/V4/V2/v4 ;
 wire [3:0] \V3/V4/V3/s1 ;
 wire [3:0] \V3/V4/V3/s2 ;
 wire [3:0] \V3/V4/V3/v1 ;
 wire [3:0] \V3/V4/V3/v2 ;
 wire [3:0] \V3/V4/V3/v3 ;
 wire [3:0] \V3/V4/V3/v4 ;
 wire [3:0] \V3/V4/V4/s1 ;
 wire [3:0] \V3/V4/V4/s2 ;
 wire [3:0] \V3/V4/V4/v1 ;
 wire [3:0] \V3/V4/V4/v2 ;
 wire [3:0] \V3/V4/V4/v3 ;
 wire [3:0] \V3/V4/V4/v4 ;
 wire [7:0] \V3/V4/s1 ;
 wire [7:0] \V3/V4/s2 ;
 wire [7:0] \V3/V4/v1 ;
 wire [7:0] \V3/V4/v2 ;
 wire [7:0] \V3/V4/v3 ;
 wire [7:0] \V3/V4/v4 ;
 wire [15:0] \V3/s1 ;
 wire [15:0] \V3/s2 ;
 wire [15:0] \V3/v1 ;
 wire [15:0] \V3/v2 ;
 wire [15:0] \V3/v3 ;
 wire [15:0] \V3/v4 ;
 wire [3:0] \V4/V1/V1/s1 ;
 wire [3:0] \V4/V1/V1/s2 ;
 wire [3:0] \V4/V1/V1/v1 ;
 wire [3:0] \V4/V1/V1/v2 ;
 wire [3:0] \V4/V1/V1/v3 ;
 wire [3:0] \V4/V1/V1/v4 ;
 wire [3:0] \V4/V1/V2/s1 ;
 wire [3:0] \V4/V1/V2/s2 ;
 wire [3:0] \V4/V1/V2/v1 ;
 wire [3:0] \V4/V1/V2/v2 ;
 wire [3:0] \V4/V1/V2/v3 ;
 wire [3:0] \V4/V1/V2/v4 ;
 wire [3:0] \V4/V1/V3/s1 ;
 wire [3:0] \V4/V1/V3/s2 ;
 wire [3:0] \V4/V1/V3/v1 ;
 wire [3:0] \V4/V1/V3/v2 ;
 wire [3:0] \V4/V1/V3/v3 ;
 wire [3:0] \V4/V1/V3/v4 ;
 wire [3:0] \V4/V1/V4/s1 ;
 wire [3:0] \V4/V1/V4/s2 ;
 wire [3:0] \V4/V1/V4/v1 ;
 wire [3:0] \V4/V1/V4/v2 ;
 wire [3:0] \V4/V1/V4/v3 ;
 wire [3:0] \V4/V1/V4/v4 ;
 wire [7:0] \V4/V1/s1 ;
 wire [7:0] \V4/V1/s2 ;
 wire [7:0] \V4/V1/v1 ;
 wire [7:0] \V4/V1/v2 ;
 wire [7:0] \V4/V1/v3 ;
 wire [7:0] \V4/V1/v4 ;
 wire [3:0] \V4/V2/V1/s1 ;
 wire [3:0] \V4/V2/V1/s2 ;
 wire [3:0] \V4/V2/V1/v1 ;
 wire [3:0] \V4/V2/V1/v2 ;
 wire [3:0] \V4/V2/V1/v3 ;
 wire [3:0] \V4/V2/V1/v4 ;
 wire [3:0] \V4/V2/V2/s1 ;
 wire [3:0] \V4/V2/V2/s2 ;
 wire [3:0] \V4/V2/V2/v1 ;
 wire [3:0] \V4/V2/V2/v2 ;
 wire [3:0] \V4/V2/V2/v3 ;
 wire [3:0] \V4/V2/V2/v4 ;
 wire [3:0] \V4/V2/V3/s1 ;
 wire [3:0] \V4/V2/V3/s2 ;
 wire [3:0] \V4/V2/V3/v1 ;
 wire [3:0] \V4/V2/V3/v2 ;
 wire [3:0] \V4/V2/V3/v3 ;
 wire [3:0] \V4/V2/V3/v4 ;
 wire [3:0] \V4/V2/V4/s1 ;
 wire [3:0] \V4/V2/V4/s2 ;
 wire [3:0] \V4/V2/V4/v1 ;
 wire [3:0] \V4/V2/V4/v2 ;
 wire [3:0] \V4/V2/V4/v3 ;
 wire [3:0] \V4/V2/V4/v4 ;
 wire [7:0] \V4/V2/s1 ;
 wire [7:0] \V4/V2/s2 ;
 wire [7:0] \V4/V2/v1 ;
 wire [7:0] \V4/V2/v2 ;
 wire [7:0] \V4/V2/v3 ;
 wire [7:0] \V4/V2/v4 ;
 wire [3:0] \V4/V3/V1/s1 ;
 wire [3:0] \V4/V3/V1/s2 ;
 wire [3:0] \V4/V3/V1/v1 ;
 wire [3:0] \V4/V3/V1/v2 ;
 wire [3:0] \V4/V3/V1/v3 ;
 wire [3:0] \V4/V3/V1/v4 ;
 wire [3:0] \V4/V3/V2/s1 ;
 wire [3:0] \V4/V3/V2/s2 ;
 wire [3:0] \V4/V3/V2/v1 ;
 wire [3:0] \V4/V3/V2/v2 ;
 wire [3:0] \V4/V3/V2/v3 ;
 wire [3:0] \V4/V3/V2/v4 ;
 wire [3:0] \V4/V3/V3/s1 ;
 wire [3:0] \V4/V3/V3/s2 ;
 wire [3:0] \V4/V3/V3/v1 ;
 wire [3:0] \V4/V3/V3/v2 ;
 wire [3:0] \V4/V3/V3/v3 ;
 wire [3:0] \V4/V3/V3/v4 ;
 wire [3:0] \V4/V3/V4/s1 ;
 wire [3:0] \V4/V3/V4/s2 ;
 wire [3:0] \V4/V3/V4/v1 ;
 wire [3:0] \V4/V3/V4/v2 ;
 wire [3:0] \V4/V3/V4/v3 ;
 wire [3:0] \V4/V3/V4/v4 ;
 wire [7:0] \V4/V3/s1 ;
 wire [7:0] \V4/V3/s2 ;
 wire [7:0] \V4/V3/v1 ;
 wire [7:0] \V4/V3/v2 ;
 wire [7:0] \V4/V3/v3 ;
 wire [7:0] \V4/V3/v4 ;
 wire [3:0] \V4/V4/V1/s1 ;
 wire [3:0] \V4/V4/V1/s2 ;
 wire [3:0] \V4/V4/V1/v1 ;
 wire [3:0] \V4/V4/V1/v2 ;
 wire [3:0] \V4/V4/V1/v3 ;
 wire [3:0] \V4/V4/V1/v4 ;
 wire [3:0] \V4/V4/V2/s1 ;
 wire [3:0] \V4/V4/V2/s2 ;
 wire [3:0] \V4/V4/V2/v1 ;
 wire [3:0] \V4/V4/V2/v2 ;
 wire [3:0] \V4/V4/V2/v3 ;
 wire [3:0] \V4/V4/V2/v4 ;
 wire [3:0] \V4/V4/V3/s1 ;
 wire [3:0] \V4/V4/V3/s2 ;
 wire [3:0] \V4/V4/V3/v1 ;
 wire [3:0] \V4/V4/V3/v2 ;
 wire [3:0] \V4/V4/V3/v3 ;
 wire [3:0] \V4/V4/V3/v4 ;
 wire [3:0] \V4/V4/V4/s1 ;
 wire [3:0] \V4/V4/V4/s2 ;
 wire [3:0] \V4/V4/V4/v1 ;
 wire [3:0] \V4/V4/V4/v2 ;
 wire [3:0] \V4/V4/V4/v3 ;
 wire [3:0] \V4/V4/V4/v4 ;
 wire [7:0] \V4/V4/s1 ;
 wire [7:0] \V4/V4/s2 ;
 wire [7:0] \V4/V4/v1 ;
 wire [7:0] \V4/V4/v2 ;
 wire [7:0] \V4/V4/v3 ;
 wire [7:0] \V4/V4/v4 ;
 wire [15:0] \V4/s1 ;
 wire [15:0] \V4/s2 ;
 wire [15:0] \V4/v1 ;
 wire [15:0] \V4/v2 ;
 wire [15:0] \V4/v3 ;
 wire [15:0] \V4/v4 ;
 wire [31:0] s1;
 wire [31:0] s2;
 wire [31:0] v1;
 wire [31:0] v2;
 wire [31:0] v3;
 wire [31:0] v4;

 AND2_X1 \A1/A1/A1/A1/M1/M1/_0_  (.A1(v2[0]),
    .A2(v3[0]),
    .ZN(\A1/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M1/M1/_1_  (.A(v2[0]),
    .B(v3[0]),
    .Z(\A1/A1/A1/A1/M1/s1 ));
 AND2_X1 \A1/A1/A1/A1/M1/M2/_0_  (.A1(\A1/A1/A1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\A1/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M1/M2/_1_  (.A(\A1/A1/A1/A1/M1/s1 ),
    .B(net3),
    .Z(s1[0]));
 OR2_X1 \A1/A1/A1/A1/M1/_0_  (.A1(\A1/A1/A1/A1/M1/c1 ),
    .A2(\A1/A1/A1/A1/M1/c2 ),
    .ZN(\A1/A1/A1/A1/c1 ));
 AND2_X1 \A1/A1/A1/A1/M2/M1/_0_  (.A1(v2[1]),
    .A2(v3[1]),
    .ZN(\A1/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M2/M1/_1_  (.A(v2[1]),
    .B(v3[1]),
    .Z(\A1/A1/A1/A1/M2/s1 ));
 AND2_X1 \A1/A1/A1/A1/M2/M2/_0_  (.A1(\A1/A1/A1/A1/M2/s1 ),
    .A2(\A1/A1/A1/A1/c1 ),
    .ZN(\A1/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M2/M2/_1_  (.A(\A1/A1/A1/A1/M2/s1 ),
    .B(\A1/A1/A1/A1/c1 ),
    .Z(s1[1]));
 OR2_X1 \A1/A1/A1/A1/M2/_0_  (.A1(\A1/A1/A1/A1/M2/c1 ),
    .A2(\A1/A1/A1/A1/M2/c2 ),
    .ZN(\A1/A1/A1/A1/c2 ));
 AND2_X1 \A1/A1/A1/A1/M3/M1/_0_  (.A1(v2[2]),
    .A2(v3[2]),
    .ZN(\A1/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M3/M1/_1_  (.A(v2[2]),
    .B(v3[2]),
    .Z(\A1/A1/A1/A1/M3/s1 ));
 AND2_X1 \A1/A1/A1/A1/M3/M2/_0_  (.A1(\A1/A1/A1/A1/M3/s1 ),
    .A2(\A1/A1/A1/A1/c2 ),
    .ZN(\A1/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M3/M2/_1_  (.A(\A1/A1/A1/A1/M3/s1 ),
    .B(\A1/A1/A1/A1/c2 ),
    .Z(s1[2]));
 OR2_X1 \A1/A1/A1/A1/M3/_0_  (.A1(\A1/A1/A1/A1/M3/c1 ),
    .A2(\A1/A1/A1/A1/M3/c2 ),
    .ZN(\A1/A1/A1/A1/c3 ));
 AND2_X1 \A1/A1/A1/A1/M4/M1/_0_  (.A1(v2[3]),
    .A2(v3[3]),
    .ZN(\A1/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A1/A1/A1/A1/M4/M1/_1_  (.A(v2[3]),
    .B(v3[3]),
    .Z(\A1/A1/A1/A1/M4/s1 ));
 AND2_X1 \A1/A1/A1/A1/M4/M2/_0_  (.A1(\A1/A1/A1/A1/M4/s1 ),
    .A2(\A1/A1/A1/A1/c3 ),
    .ZN(\A1/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A1/A1/A1/A1/M4/M2/_1_  (.A(\A1/A1/A1/A1/M4/s1 ),
    .B(\A1/A1/A1/A1/c3 ),
    .Z(s1[3]));
 OR2_X1 \A1/A1/A1/A1/M4/_0_  (.A1(\A1/A1/A1/A1/M4/c1 ),
    .A2(\A1/A1/A1/A1/M4/c2 ),
    .ZN(\A1/A1/A1/c1 ));
 AND2_X1 \A1/A1/A1/A2/M1/M1/_0_  (.A1(v2[4]),
    .A2(v3[4]),
    .ZN(\A1/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M1/M1/_1_  (.A(v2[4]),
    .B(v3[4]),
    .Z(\A1/A1/A1/A2/M1/s1 ));
 AND2_X1 \A1/A1/A1/A2/M1/M2/_0_  (.A1(\A1/A1/A1/A2/M1/s1 ),
    .A2(\A1/A1/A1/c1 ),
    .ZN(\A1/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M1/M2/_1_  (.A(\A1/A1/A1/A2/M1/s1 ),
    .B(\A1/A1/A1/c1 ),
    .Z(s1[4]));
 OR2_X1 \A1/A1/A1/A2/M1/_0_  (.A1(\A1/A1/A1/A2/M1/c1 ),
    .A2(\A1/A1/A1/A2/M1/c2 ),
    .ZN(\A1/A1/A1/A2/c1 ));
 AND2_X1 \A1/A1/A1/A2/M2/M1/_0_  (.A1(v2[5]),
    .A2(v3[5]),
    .ZN(\A1/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M2/M1/_1_  (.A(v2[5]),
    .B(v3[5]),
    .Z(\A1/A1/A1/A2/M2/s1 ));
 AND2_X1 \A1/A1/A1/A2/M2/M2/_0_  (.A1(\A1/A1/A1/A2/M2/s1 ),
    .A2(\A1/A1/A1/A2/c1 ),
    .ZN(\A1/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M2/M2/_1_  (.A(\A1/A1/A1/A2/M2/s1 ),
    .B(\A1/A1/A1/A2/c1 ),
    .Z(s1[5]));
 OR2_X1 \A1/A1/A1/A2/M2/_0_  (.A1(\A1/A1/A1/A2/M2/c1 ),
    .A2(\A1/A1/A1/A2/M2/c2 ),
    .ZN(\A1/A1/A1/A2/c2 ));
 AND2_X1 \A1/A1/A1/A2/M3/M1/_0_  (.A1(v2[6]),
    .A2(v3[6]),
    .ZN(\A1/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M3/M1/_1_  (.A(v2[6]),
    .B(v3[6]),
    .Z(\A1/A1/A1/A2/M3/s1 ));
 AND2_X1 \A1/A1/A1/A2/M3/M2/_0_  (.A1(\A1/A1/A1/A2/M3/s1 ),
    .A2(\A1/A1/A1/A2/c2 ),
    .ZN(\A1/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M3/M2/_1_  (.A(\A1/A1/A1/A2/M3/s1 ),
    .B(\A1/A1/A1/A2/c2 ),
    .Z(s1[6]));
 OR2_X1 \A1/A1/A1/A2/M3/_0_  (.A1(\A1/A1/A1/A2/M3/c1 ),
    .A2(\A1/A1/A1/A2/M3/c2 ),
    .ZN(\A1/A1/A1/A2/c3 ));
 AND2_X1 \A1/A1/A1/A2/M4/M1/_0_  (.A1(v2[7]),
    .A2(v3[7]),
    .ZN(\A1/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A1/A1/A1/A2/M4/M1/_1_  (.A(v2[7]),
    .B(v3[7]),
    .Z(\A1/A1/A1/A2/M4/s1 ));
 AND2_X1 \A1/A1/A1/A2/M4/M2/_0_  (.A1(\A1/A1/A1/A2/M4/s1 ),
    .A2(\A1/A1/A1/A2/c3 ),
    .ZN(\A1/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A1/A1/A1/A2/M4/M2/_1_  (.A(\A1/A1/A1/A2/M4/s1 ),
    .B(\A1/A1/A1/A2/c3 ),
    .Z(s1[7]));
 OR2_X2 \A1/A1/A1/A2/M4/_0_  (.A1(\A1/A1/A1/A2/M4/c1 ),
    .A2(\A1/A1/A1/A2/M4/c2 ),
    .ZN(\A1/A1/c1 ));
 AND2_X1 \A1/A1/A2/A1/M1/M1/_0_  (.A1(v2[8]),
    .A2(v3[8]),
    .ZN(\A1/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M1/M1/_1_  (.A(v2[8]),
    .B(v3[8]),
    .Z(\A1/A1/A2/A1/M1/s1 ));
 AND2_X1 \A1/A1/A2/A1/M1/M2/_0_  (.A1(\A1/A1/A2/A1/M1/s1 ),
    .A2(\A1/A1/c1 ),
    .ZN(\A1/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M1/M2/_1_  (.A(\A1/A1/A2/A1/M1/s1 ),
    .B(\A1/A1/c1 ),
    .Z(s1[8]));
 OR2_X1 \A1/A1/A2/A1/M1/_0_  (.A1(\A1/A1/A2/A1/M1/c1 ),
    .A2(\A1/A1/A2/A1/M1/c2 ),
    .ZN(\A1/A1/A2/A1/c1 ));
 AND2_X1 \A1/A1/A2/A1/M2/M1/_0_  (.A1(v2[9]),
    .A2(v3[9]),
    .ZN(\A1/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M2/M1/_1_  (.A(v2[9]),
    .B(v3[9]),
    .Z(\A1/A1/A2/A1/M2/s1 ));
 AND2_X1 \A1/A1/A2/A1/M2/M2/_0_  (.A1(\A1/A1/A2/A1/M2/s1 ),
    .A2(\A1/A1/A2/A1/c1 ),
    .ZN(\A1/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M2/M2/_1_  (.A(\A1/A1/A2/A1/M2/s1 ),
    .B(\A1/A1/A2/A1/c1 ),
    .Z(s1[9]));
 OR2_X1 \A1/A1/A2/A1/M2/_0_  (.A1(\A1/A1/A2/A1/M2/c1 ),
    .A2(\A1/A1/A2/A1/M2/c2 ),
    .ZN(\A1/A1/A2/A1/c2 ));
 AND2_X1 \A1/A1/A2/A1/M3/M1/_0_  (.A1(v2[10]),
    .A2(v3[10]),
    .ZN(\A1/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M3/M1/_1_  (.A(v2[10]),
    .B(v3[10]),
    .Z(\A1/A1/A2/A1/M3/s1 ));
 AND2_X1 \A1/A1/A2/A1/M3/M2/_0_  (.A1(\A1/A1/A2/A1/M3/s1 ),
    .A2(\A1/A1/A2/A1/c2 ),
    .ZN(\A1/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M3/M2/_1_  (.A(\A1/A1/A2/A1/M3/s1 ),
    .B(\A1/A1/A2/A1/c2 ),
    .Z(s1[10]));
 OR2_X1 \A1/A1/A2/A1/M3/_0_  (.A1(\A1/A1/A2/A1/M3/c1 ),
    .A2(\A1/A1/A2/A1/M3/c2 ),
    .ZN(\A1/A1/A2/A1/c3 ));
 AND2_X1 \A1/A1/A2/A1/M4/M1/_0_  (.A1(v2[11]),
    .A2(v3[11]),
    .ZN(\A1/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A1/A1/A2/A1/M4/M1/_1_  (.A(v2[11]),
    .B(v3[11]),
    .Z(\A1/A1/A2/A1/M4/s1 ));
 AND2_X1 \A1/A1/A2/A1/M4/M2/_0_  (.A1(\A1/A1/A2/A1/M4/s1 ),
    .A2(\A1/A1/A2/A1/c3 ),
    .ZN(\A1/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A1/A1/A2/A1/M4/M2/_1_  (.A(\A1/A1/A2/A1/M4/s1 ),
    .B(\A1/A1/A2/A1/c3 ),
    .Z(s1[11]));
 OR2_X1 \A1/A1/A2/A1/M4/_0_  (.A1(\A1/A1/A2/A1/M4/c1 ),
    .A2(\A1/A1/A2/A1/M4/c2 ),
    .ZN(\A1/A1/A2/c1 ));
 AND2_X1 \A1/A1/A2/A2/M1/M1/_0_  (.A1(v2[12]),
    .A2(v3[12]),
    .ZN(\A1/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M1/M1/_1_  (.A(v2[12]),
    .B(v3[12]),
    .Z(\A1/A1/A2/A2/M1/s1 ));
 AND2_X1 \A1/A1/A2/A2/M1/M2/_0_  (.A1(\A1/A1/A2/A2/M1/s1 ),
    .A2(\A1/A1/A2/c1 ),
    .ZN(\A1/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M1/M2/_1_  (.A(\A1/A1/A2/A2/M1/s1 ),
    .B(\A1/A1/A2/c1 ),
    .Z(s1[12]));
 OR2_X1 \A1/A1/A2/A2/M1/_0_  (.A1(\A1/A1/A2/A2/M1/c1 ),
    .A2(\A1/A1/A2/A2/M1/c2 ),
    .ZN(\A1/A1/A2/A2/c1 ));
 AND2_X1 \A1/A1/A2/A2/M2/M1/_0_  (.A1(v2[13]),
    .A2(v3[13]),
    .ZN(\A1/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M2/M1/_1_  (.A(v2[13]),
    .B(v3[13]),
    .Z(\A1/A1/A2/A2/M2/s1 ));
 AND2_X1 \A1/A1/A2/A2/M2/M2/_0_  (.A1(\A1/A1/A2/A2/M2/s1 ),
    .A2(\A1/A1/A2/A2/c1 ),
    .ZN(\A1/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M2/M2/_1_  (.A(\A1/A1/A2/A2/M2/s1 ),
    .B(\A1/A1/A2/A2/c1 ),
    .Z(s1[13]));
 OR2_X1 \A1/A1/A2/A2/M2/_0_  (.A1(\A1/A1/A2/A2/M2/c1 ),
    .A2(\A1/A1/A2/A2/M2/c2 ),
    .ZN(\A1/A1/A2/A2/c2 ));
 AND2_X1 \A1/A1/A2/A2/M3/M1/_0_  (.A1(v2[14]),
    .A2(v3[14]),
    .ZN(\A1/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M3/M1/_1_  (.A(v2[14]),
    .B(v3[14]),
    .Z(\A1/A1/A2/A2/M3/s1 ));
 AND2_X1 \A1/A1/A2/A2/M3/M2/_0_  (.A1(\A1/A1/A2/A2/M3/s1 ),
    .A2(\A1/A1/A2/A2/c2 ),
    .ZN(\A1/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M3/M2/_1_  (.A(\A1/A1/A2/A2/M3/s1 ),
    .B(\A1/A1/A2/A2/c2 ),
    .Z(s1[14]));
 OR2_X1 \A1/A1/A2/A2/M3/_0_  (.A1(\A1/A1/A2/A2/M3/c1 ),
    .A2(\A1/A1/A2/A2/M3/c2 ),
    .ZN(\A1/A1/A2/A2/c3 ));
 AND2_X1 \A1/A1/A2/A2/M4/M1/_0_  (.A1(v2[15]),
    .A2(v3[15]),
    .ZN(\A1/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A1/A1/A2/A2/M4/M1/_1_  (.A(v2[15]),
    .B(v3[15]),
    .Z(\A1/A1/A2/A2/M4/s1 ));
 AND2_X1 \A1/A1/A2/A2/M4/M2/_0_  (.A1(\A1/A1/A2/A2/M4/s1 ),
    .A2(\A1/A1/A2/A2/c3 ),
    .ZN(\A1/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A1/A1/A2/A2/M4/M2/_1_  (.A(\A1/A1/A2/A2/M4/s1 ),
    .B(\A1/A1/A2/A2/c3 ),
    .Z(s1[15]));
 OR2_X1 \A1/A1/A2/A2/M4/_0_  (.A1(\A1/A1/A2/A2/M4/c1 ),
    .A2(\A1/A1/A2/A2/M4/c2 ),
    .ZN(\A1/c1 ));
 AND2_X1 \A1/A2/A1/A1/M1/M1/_0_  (.A1(v2[16]),
    .A2(v3[16]),
    .ZN(\A1/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M1/M1/_1_  (.A(v2[16]),
    .B(v3[16]),
    .Z(\A1/A2/A1/A1/M1/s1 ));
 AND2_X1 \A1/A2/A1/A1/M1/M2/_0_  (.A1(\A1/A2/A1/A1/M1/s1 ),
    .A2(net7),
    .ZN(\A1/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M1/M2/_1_  (.A(\A1/A2/A1/A1/M1/s1 ),
    .B(net2),
    .Z(s1[16]));
 OR2_X1 \A1/A2/A1/A1/M1/_0_  (.A1(\A1/A2/A1/A1/M1/c1 ),
    .A2(\A1/A2/A1/A1/M1/c2 ),
    .ZN(\A1/A2/A1/A1/c1 ));
 AND2_X1 \A1/A2/A1/A1/M2/M1/_0_  (.A1(v2[17]),
    .A2(v3[17]),
    .ZN(\A1/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M2/M1/_1_  (.A(v2[17]),
    .B(v3[17]),
    .Z(\A1/A2/A1/A1/M2/s1 ));
 AND2_X1 \A1/A2/A1/A1/M2/M2/_0_  (.A1(\A1/A2/A1/A1/M2/s1 ),
    .A2(\A1/A2/A1/A1/c1 ),
    .ZN(\A1/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M2/M2/_1_  (.A(\A1/A2/A1/A1/M2/s1 ),
    .B(\A1/A2/A1/A1/c1 ),
    .Z(s1[17]));
 OR2_X1 \A1/A2/A1/A1/M2/_0_  (.A1(\A1/A2/A1/A1/M2/c1 ),
    .A2(\A1/A2/A1/A1/M2/c2 ),
    .ZN(\A1/A2/A1/A1/c2 ));
 AND2_X1 \A1/A2/A1/A1/M3/M1/_0_  (.A1(v2[18]),
    .A2(v3[18]),
    .ZN(\A1/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M3/M1/_1_  (.A(v2[18]),
    .B(v3[18]),
    .Z(\A1/A2/A1/A1/M3/s1 ));
 AND2_X1 \A1/A2/A1/A1/M3/M2/_0_  (.A1(\A1/A2/A1/A1/M3/s1 ),
    .A2(\A1/A2/A1/A1/c2 ),
    .ZN(\A1/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M3/M2/_1_  (.A(\A1/A2/A1/A1/M3/s1 ),
    .B(\A1/A2/A1/A1/c2 ),
    .Z(s1[18]));
 OR2_X1 \A1/A2/A1/A1/M3/_0_  (.A1(\A1/A2/A1/A1/M3/c1 ),
    .A2(\A1/A2/A1/A1/M3/c2 ),
    .ZN(\A1/A2/A1/A1/c3 ));
 AND2_X1 \A1/A2/A1/A1/M4/M1/_0_  (.A1(v2[19]),
    .A2(v3[19]),
    .ZN(\A1/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A1/A2/A1/A1/M4/M1/_1_  (.A(v2[19]),
    .B(v3[19]),
    .Z(\A1/A2/A1/A1/M4/s1 ));
 AND2_X1 \A1/A2/A1/A1/M4/M2/_0_  (.A1(\A1/A2/A1/A1/M4/s1 ),
    .A2(\A1/A2/A1/A1/c3 ),
    .ZN(\A1/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A1/A2/A1/A1/M4/M2/_1_  (.A(\A1/A2/A1/A1/M4/s1 ),
    .B(\A1/A2/A1/A1/c3 ),
    .Z(s1[19]));
 OR2_X1 \A1/A2/A1/A1/M4/_0_  (.A1(\A1/A2/A1/A1/M4/c1 ),
    .A2(\A1/A2/A1/A1/M4/c2 ),
    .ZN(\A1/A2/A1/c1 ));
 AND2_X1 \A1/A2/A1/A2/M1/M1/_0_  (.A1(v2[20]),
    .A2(v3[20]),
    .ZN(\A1/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M1/M1/_1_  (.A(v2[20]),
    .B(v3[20]),
    .Z(\A1/A2/A1/A2/M1/s1 ));
 AND2_X1 \A1/A2/A1/A2/M1/M2/_0_  (.A1(\A1/A2/A1/A2/M1/s1 ),
    .A2(\A1/A2/A1/c1 ),
    .ZN(\A1/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M1/M2/_1_  (.A(\A1/A2/A1/A2/M1/s1 ),
    .B(\A1/A2/A1/c1 ),
    .Z(s1[20]));
 OR2_X1 \A1/A2/A1/A2/M1/_0_  (.A1(\A1/A2/A1/A2/M1/c1 ),
    .A2(\A1/A2/A1/A2/M1/c2 ),
    .ZN(\A1/A2/A1/A2/c1 ));
 AND2_X1 \A1/A2/A1/A2/M2/M1/_0_  (.A1(v2[21]),
    .A2(v3[21]),
    .ZN(\A1/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M2/M1/_1_  (.A(v2[21]),
    .B(v3[21]),
    .Z(\A1/A2/A1/A2/M2/s1 ));
 AND2_X1 \A1/A2/A1/A2/M2/M2/_0_  (.A1(\A1/A2/A1/A2/M2/s1 ),
    .A2(\A1/A2/A1/A2/c1 ),
    .ZN(\A1/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M2/M2/_1_  (.A(\A1/A2/A1/A2/M2/s1 ),
    .B(\A1/A2/A1/A2/c1 ),
    .Z(s1[21]));
 OR2_X1 \A1/A2/A1/A2/M2/_0_  (.A1(\A1/A2/A1/A2/M2/c1 ),
    .A2(\A1/A2/A1/A2/M2/c2 ),
    .ZN(\A1/A2/A1/A2/c2 ));
 AND2_X1 \A1/A2/A1/A2/M3/M1/_0_  (.A1(v2[22]),
    .A2(v3[22]),
    .ZN(\A1/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M3/M1/_1_  (.A(v2[22]),
    .B(v3[22]),
    .Z(\A1/A2/A1/A2/M3/s1 ));
 AND2_X1 \A1/A2/A1/A2/M3/M2/_0_  (.A1(\A1/A2/A1/A2/M3/s1 ),
    .A2(\A1/A2/A1/A2/c2 ),
    .ZN(\A1/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M3/M2/_1_  (.A(\A1/A2/A1/A2/M3/s1 ),
    .B(\A1/A2/A1/A2/c2 ),
    .Z(s1[22]));
 OR2_X1 \A1/A2/A1/A2/M3/_0_  (.A1(\A1/A2/A1/A2/M3/c1 ),
    .A2(\A1/A2/A1/A2/M3/c2 ),
    .ZN(\A1/A2/A1/A2/c3 ));
 AND2_X1 \A1/A2/A1/A2/M4/M1/_0_  (.A1(v2[23]),
    .A2(v3[23]),
    .ZN(\A1/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A1/A2/A1/A2/M4/M1/_1_  (.A(v2[23]),
    .B(v3[23]),
    .Z(\A1/A2/A1/A2/M4/s1 ));
 AND2_X1 \A1/A2/A1/A2/M4/M2/_0_  (.A1(\A1/A2/A1/A2/M4/s1 ),
    .A2(\A1/A2/A1/A2/c3 ),
    .ZN(\A1/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A1/A2/A1/A2/M4/M2/_1_  (.A(\A1/A2/A1/A2/M4/s1 ),
    .B(\A1/A2/A1/A2/c3 ),
    .Z(s1[23]));
 OR2_X1 \A1/A2/A1/A2/M4/_0_  (.A1(\A1/A2/A1/A2/M4/c1 ),
    .A2(\A1/A2/A1/A2/M4/c2 ),
    .ZN(\A1/A2/c1 ));
 AND2_X1 \A1/A2/A2/A1/M1/M1/_0_  (.A1(v2[24]),
    .A2(v3[24]),
    .ZN(\A1/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M1/M1/_1_  (.A(v2[24]),
    .B(v3[24]),
    .Z(\A1/A2/A2/A1/M1/s1 ));
 AND2_X1 \A1/A2/A2/A1/M1/M2/_0_  (.A1(\A1/A2/A2/A1/M1/s1 ),
    .A2(\A1/A2/c1 ),
    .ZN(\A1/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M1/M2/_1_  (.A(\A1/A2/A2/A1/M1/s1 ),
    .B(\A1/A2/c1 ),
    .Z(s1[24]));
 OR2_X1 \A1/A2/A2/A1/M1/_0_  (.A1(\A1/A2/A2/A1/M1/c1 ),
    .A2(\A1/A2/A2/A1/M1/c2 ),
    .ZN(\A1/A2/A2/A1/c1 ));
 AND2_X1 \A1/A2/A2/A1/M2/M1/_0_  (.A1(v2[25]),
    .A2(v3[25]),
    .ZN(\A1/A2/A2/A1/M2/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M2/M1/_1_  (.A(v2[25]),
    .B(v3[25]),
    .Z(\A1/A2/A2/A1/M2/s1 ));
 AND2_X1 \A1/A2/A2/A1/M2/M2/_0_  (.A1(\A1/A2/A2/A1/M2/s1 ),
    .A2(\A1/A2/A2/A1/c1 ),
    .ZN(\A1/A2/A2/A1/M2/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M2/M2/_1_  (.A(\A1/A2/A2/A1/M2/s1 ),
    .B(\A1/A2/A2/A1/c1 ),
    .Z(s1[25]));
 OR2_X1 \A1/A2/A2/A1/M2/_0_  (.A1(\A1/A2/A2/A1/M2/c1 ),
    .A2(\A1/A2/A2/A1/M2/c2 ),
    .ZN(\A1/A2/A2/A1/c2 ));
 AND2_X1 \A1/A2/A2/A1/M3/M1/_0_  (.A1(v2[26]),
    .A2(v3[26]),
    .ZN(\A1/A2/A2/A1/M3/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M3/M1/_1_  (.A(v2[26]),
    .B(v3[26]),
    .Z(\A1/A2/A2/A1/M3/s1 ));
 AND2_X1 \A1/A2/A2/A1/M3/M2/_0_  (.A1(\A1/A2/A2/A1/M3/s1 ),
    .A2(\A1/A2/A2/A1/c2 ),
    .ZN(\A1/A2/A2/A1/M3/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M3/M2/_1_  (.A(\A1/A2/A2/A1/M3/s1 ),
    .B(\A1/A2/A2/A1/c2 ),
    .Z(s1[26]));
 OR2_X1 \A1/A2/A2/A1/M3/_0_  (.A1(\A1/A2/A2/A1/M3/c1 ),
    .A2(\A1/A2/A2/A1/M3/c2 ),
    .ZN(\A1/A2/A2/A1/c3 ));
 AND2_X1 \A1/A2/A2/A1/M4/M1/_0_  (.A1(v2[27]),
    .A2(v3[27]),
    .ZN(\A1/A2/A2/A1/M4/c1 ));
 XOR2_X2 \A1/A2/A2/A1/M4/M1/_1_  (.A(v2[27]),
    .B(v3[27]),
    .Z(\A1/A2/A2/A1/M4/s1 ));
 AND2_X1 \A1/A2/A2/A1/M4/M2/_0_  (.A1(\A1/A2/A2/A1/M4/s1 ),
    .A2(\A1/A2/A2/A1/c3 ),
    .ZN(\A1/A2/A2/A1/M4/c2 ));
 XOR2_X2 \A1/A2/A2/A1/M4/M2/_1_  (.A(\A1/A2/A2/A1/M4/s1 ),
    .B(\A1/A2/A2/A1/c3 ),
    .Z(s1[27]));
 OR2_X1 \A1/A2/A2/A1/M4/_0_  (.A1(\A1/A2/A2/A1/M4/c1 ),
    .A2(\A1/A2/A2/A1/M4/c2 ),
    .ZN(\A1/A2/A2/c1 ));
 AND2_X1 \A1/A2/A2/A2/M1/M1/_0_  (.A1(v2[28]),
    .A2(v3[28]),
    .ZN(\A1/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M1/M1/_1_  (.A(v2[28]),
    .B(v3[28]),
    .Z(\A1/A2/A2/A2/M1/s1 ));
 AND2_X1 \A1/A2/A2/A2/M1/M2/_0_  (.A1(\A1/A2/A2/A2/M1/s1 ),
    .A2(\A1/A2/A2/c1 ),
    .ZN(\A1/A2/A2/A2/M1/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M1/M2/_1_  (.A(\A1/A2/A2/A2/M1/s1 ),
    .B(\A1/A2/A2/c1 ),
    .Z(s1[28]));
 OR2_X1 \A1/A2/A2/A2/M1/_0_  (.A1(\A1/A2/A2/A2/M1/c1 ),
    .A2(\A1/A2/A2/A2/M1/c2 ),
    .ZN(\A1/A2/A2/A2/c1 ));
 AND2_X1 \A1/A2/A2/A2/M2/M1/_0_  (.A1(v2[29]),
    .A2(v3[29]),
    .ZN(\A1/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M2/M1/_1_  (.A(v2[29]),
    .B(v3[29]),
    .Z(\A1/A2/A2/A2/M2/s1 ));
 AND2_X1 \A1/A2/A2/A2/M2/M2/_0_  (.A1(\A1/A2/A2/A2/M2/s1 ),
    .A2(\A1/A2/A2/A2/c1 ),
    .ZN(\A1/A2/A2/A2/M2/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M2/M2/_1_  (.A(\A1/A2/A2/A2/M2/s1 ),
    .B(\A1/A2/A2/A2/c1 ),
    .Z(s1[29]));
 OR2_X1 \A1/A2/A2/A2/M2/_0_  (.A1(\A1/A2/A2/A2/M2/c1 ),
    .A2(\A1/A2/A2/A2/M2/c2 ),
    .ZN(\A1/A2/A2/A2/c2 ));
 AND2_X1 \A1/A2/A2/A2/M3/M1/_0_  (.A1(v2[30]),
    .A2(v3[30]),
    .ZN(\A1/A2/A2/A2/M3/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M3/M1/_1_  (.A(v2[30]),
    .B(v3[30]),
    .Z(\A1/A2/A2/A2/M3/s1 ));
 AND2_X1 \A1/A2/A2/A2/M3/M2/_0_  (.A1(\A1/A2/A2/A2/M3/s1 ),
    .A2(\A1/A2/A2/A2/c2 ),
    .ZN(\A1/A2/A2/A2/M3/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M3/M2/_1_  (.A(\A1/A2/A2/A2/M3/s1 ),
    .B(\A1/A2/A2/A2/c2 ),
    .Z(s1[30]));
 OR2_X1 \A1/A2/A2/A2/M3/_0_  (.A1(\A1/A2/A2/A2/M3/c1 ),
    .A2(\A1/A2/A2/A2/M3/c2 ),
    .ZN(\A1/A2/A2/A2/c3 ));
 AND2_X1 \A1/A2/A2/A2/M4/M1/_0_  (.A1(v2[31]),
    .A2(v3[31]),
    .ZN(\A1/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A1/A2/A2/A2/M4/M1/_1_  (.A(v2[31]),
    .B(v3[31]),
    .Z(\A1/A2/A2/A2/M4/s1 ));
 AND2_X1 \A1/A2/A2/A2/M4/M2/_0_  (.A1(\A1/A2/A2/A2/M4/s1 ),
    .A2(\A1/A2/A2/A2/c3 ),
    .ZN(\A1/A2/A2/A2/M4/c2 ));
 XOR2_X2 \A1/A2/A2/A2/M4/M2/_1_  (.A(\A1/A2/A2/A2/M4/s1 ),
    .B(\A1/A2/A2/A2/c3 ),
    .Z(s1[31]));
 OR2_X1 \A1/A2/A2/A2/M4/_0_  (.A1(\A1/A2/A2/A2/M4/c1 ),
    .A2(\A1/A2/A2/A2/M4/c2 ),
    .ZN(c1));
 AND2_X1 \A2/A1/A1/A1/M1/M1/_0_  (.A1(s1[0]),
    .A2(v1[16]),
    .ZN(\A2/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M1/M1/_1_  (.A(s1[0]),
    .B(v1[16]),
    .Z(\A2/A1/A1/A1/M1/s1 ));
 AND2_X1 \A2/A1/A1/A1/M1/M2/_0_  (.A1(\A2/A1/A1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\A2/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M1/M2/_1_  (.A(\A2/A1/A1/A1/M1/s1 ),
    .B(net3),
    .Z(s2[0]));
 OR2_X1 \A2/A1/A1/A1/M1/_0_  (.A1(\A2/A1/A1/A1/M1/c1 ),
    .A2(\A2/A1/A1/A1/M1/c2 ),
    .ZN(\A2/A1/A1/A1/c1 ));
 AND2_X1 \A2/A1/A1/A1/M2/M1/_0_  (.A1(s1[1]),
    .A2(v1[17]),
    .ZN(\A2/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M2/M1/_1_  (.A(s1[1]),
    .B(v1[17]),
    .Z(\A2/A1/A1/A1/M2/s1 ));
 AND2_X1 \A2/A1/A1/A1/M2/M2/_0_  (.A1(\A2/A1/A1/A1/M2/s1 ),
    .A2(\A2/A1/A1/A1/c1 ),
    .ZN(\A2/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M2/M2/_1_  (.A(\A2/A1/A1/A1/M2/s1 ),
    .B(\A2/A1/A1/A1/c1 ),
    .Z(s2[1]));
 OR2_X1 \A2/A1/A1/A1/M2/_0_  (.A1(\A2/A1/A1/A1/M2/c1 ),
    .A2(\A2/A1/A1/A1/M2/c2 ),
    .ZN(\A2/A1/A1/A1/c2 ));
 AND2_X1 \A2/A1/A1/A1/M3/M1/_0_  (.A1(s1[2]),
    .A2(v1[18]),
    .ZN(\A2/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M3/M1/_1_  (.A(s1[2]),
    .B(v1[18]),
    .Z(\A2/A1/A1/A1/M3/s1 ));
 AND2_X1 \A2/A1/A1/A1/M3/M2/_0_  (.A1(\A2/A1/A1/A1/M3/s1 ),
    .A2(\A2/A1/A1/A1/c2 ),
    .ZN(\A2/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M3/M2/_1_  (.A(\A2/A1/A1/A1/M3/s1 ),
    .B(\A2/A1/A1/A1/c2 ),
    .Z(s2[2]));
 OR2_X1 \A2/A1/A1/A1/M3/_0_  (.A1(\A2/A1/A1/A1/M3/c1 ),
    .A2(\A2/A1/A1/A1/M3/c2 ),
    .ZN(\A2/A1/A1/A1/c3 ));
 AND2_X1 \A2/A1/A1/A1/M4/M1/_0_  (.A1(s1[3]),
    .A2(v1[19]),
    .ZN(\A2/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A2/A1/A1/A1/M4/M1/_1_  (.A(s1[3]),
    .B(v1[19]),
    .Z(\A2/A1/A1/A1/M4/s1 ));
 AND2_X1 \A2/A1/A1/A1/M4/M2/_0_  (.A1(\A2/A1/A1/A1/M4/s1 ),
    .A2(\A2/A1/A1/A1/c3 ),
    .ZN(\A2/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A2/A1/A1/A1/M4/M2/_1_  (.A(\A2/A1/A1/A1/M4/s1 ),
    .B(\A2/A1/A1/A1/c3 ),
    .Z(s2[3]));
 OR2_X1 \A2/A1/A1/A1/M4/_0_  (.A1(\A2/A1/A1/A1/M4/c1 ),
    .A2(\A2/A1/A1/A1/M4/c2 ),
    .ZN(\A2/A1/A1/c1 ));
 AND2_X1 \A2/A1/A1/A2/M1/M1/_0_  (.A1(s1[4]),
    .A2(v1[20]),
    .ZN(\A2/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M1/M1/_1_  (.A(s1[4]),
    .B(v1[20]),
    .Z(\A2/A1/A1/A2/M1/s1 ));
 AND2_X1 \A2/A1/A1/A2/M1/M2/_0_  (.A1(\A2/A1/A1/A2/M1/s1 ),
    .A2(\A2/A1/A1/c1 ),
    .ZN(\A2/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M1/M2/_1_  (.A(\A2/A1/A1/A2/M1/s1 ),
    .B(\A2/A1/A1/c1 ),
    .Z(s2[4]));
 OR2_X1 \A2/A1/A1/A2/M1/_0_  (.A1(\A2/A1/A1/A2/M1/c1 ),
    .A2(\A2/A1/A1/A2/M1/c2 ),
    .ZN(\A2/A1/A1/A2/c1 ));
 AND2_X1 \A2/A1/A1/A2/M2/M1/_0_  (.A1(s1[5]),
    .A2(v1[21]),
    .ZN(\A2/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M2/M1/_1_  (.A(s1[5]),
    .B(v1[21]),
    .Z(\A2/A1/A1/A2/M2/s1 ));
 AND2_X1 \A2/A1/A1/A2/M2/M2/_0_  (.A1(\A2/A1/A1/A2/M2/s1 ),
    .A2(\A2/A1/A1/A2/c1 ),
    .ZN(\A2/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M2/M2/_1_  (.A(\A2/A1/A1/A2/M2/s1 ),
    .B(\A2/A1/A1/A2/c1 ),
    .Z(s2[5]));
 OR2_X1 \A2/A1/A1/A2/M2/_0_  (.A1(\A2/A1/A1/A2/M2/c1 ),
    .A2(\A2/A1/A1/A2/M2/c2 ),
    .ZN(\A2/A1/A1/A2/c2 ));
 AND2_X1 \A2/A1/A1/A2/M3/M1/_0_  (.A1(s1[6]),
    .A2(v1[22]),
    .ZN(\A2/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M3/M1/_1_  (.A(s1[6]),
    .B(v1[22]),
    .Z(\A2/A1/A1/A2/M3/s1 ));
 AND2_X1 \A2/A1/A1/A2/M3/M2/_0_  (.A1(\A2/A1/A1/A2/M3/s1 ),
    .A2(\A2/A1/A1/A2/c2 ),
    .ZN(\A2/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M3/M2/_1_  (.A(\A2/A1/A1/A2/M3/s1 ),
    .B(\A2/A1/A1/A2/c2 ),
    .Z(s2[6]));
 OR2_X1 \A2/A1/A1/A2/M3/_0_  (.A1(\A2/A1/A1/A2/M3/c1 ),
    .A2(\A2/A1/A1/A2/M3/c2 ),
    .ZN(\A2/A1/A1/A2/c3 ));
 AND2_X1 \A2/A1/A1/A2/M4/M1/_0_  (.A1(s1[7]),
    .A2(v1[23]),
    .ZN(\A2/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A2/A1/A1/A2/M4/M1/_1_  (.A(s1[7]),
    .B(v1[23]),
    .Z(\A2/A1/A1/A2/M4/s1 ));
 AND2_X1 \A2/A1/A1/A2/M4/M2/_0_  (.A1(\A2/A1/A1/A2/M4/s1 ),
    .A2(\A2/A1/A1/A2/c3 ),
    .ZN(\A2/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A2/A1/A1/A2/M4/M2/_1_  (.A(\A2/A1/A1/A2/M4/s1 ),
    .B(\A2/A1/A1/A2/c3 ),
    .Z(s2[7]));
 OR2_X2 \A2/A1/A1/A2/M4/_0_  (.A1(\A2/A1/A1/A2/M4/c1 ),
    .A2(\A2/A1/A1/A2/M4/c2 ),
    .ZN(\A2/A1/c1 ));
 AND2_X1 \A2/A1/A2/A1/M1/M1/_0_  (.A1(s1[8]),
    .A2(v1[24]),
    .ZN(\A2/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M1/M1/_1_  (.A(s1[8]),
    .B(v1[24]),
    .Z(\A2/A1/A2/A1/M1/s1 ));
 AND2_X1 \A2/A1/A2/A1/M1/M2/_0_  (.A1(\A2/A1/A2/A1/M1/s1 ),
    .A2(\A2/A1/c1 ),
    .ZN(\A2/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M1/M2/_1_  (.A(\A2/A1/A2/A1/M1/s1 ),
    .B(\A2/A1/c1 ),
    .Z(s2[8]));
 OR2_X1 \A2/A1/A2/A1/M1/_0_  (.A1(\A2/A1/A2/A1/M1/c1 ),
    .A2(\A2/A1/A2/A1/M1/c2 ),
    .ZN(\A2/A1/A2/A1/c1 ));
 AND2_X1 \A2/A1/A2/A1/M2/M1/_0_  (.A1(s1[9]),
    .A2(v1[25]),
    .ZN(\A2/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M2/M1/_1_  (.A(s1[9]),
    .B(v1[25]),
    .Z(\A2/A1/A2/A1/M2/s1 ));
 AND2_X1 \A2/A1/A2/A1/M2/M2/_0_  (.A1(\A2/A1/A2/A1/M2/s1 ),
    .A2(\A2/A1/A2/A1/c1 ),
    .ZN(\A2/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M2/M2/_1_  (.A(\A2/A1/A2/A1/M2/s1 ),
    .B(\A2/A1/A2/A1/c1 ),
    .Z(s2[9]));
 OR2_X1 \A2/A1/A2/A1/M2/_0_  (.A1(\A2/A1/A2/A1/M2/c1 ),
    .A2(\A2/A1/A2/A1/M2/c2 ),
    .ZN(\A2/A1/A2/A1/c2 ));
 AND2_X1 \A2/A1/A2/A1/M3/M1/_0_  (.A1(s1[10]),
    .A2(v1[26]),
    .ZN(\A2/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M3/M1/_1_  (.A(s1[10]),
    .B(v1[26]),
    .Z(\A2/A1/A2/A1/M3/s1 ));
 AND2_X1 \A2/A1/A2/A1/M3/M2/_0_  (.A1(\A2/A1/A2/A1/M3/s1 ),
    .A2(\A2/A1/A2/A1/c2 ),
    .ZN(\A2/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M3/M2/_1_  (.A(\A2/A1/A2/A1/M3/s1 ),
    .B(\A2/A1/A2/A1/c2 ),
    .Z(s2[10]));
 OR2_X1 \A2/A1/A2/A1/M3/_0_  (.A1(\A2/A1/A2/A1/M3/c1 ),
    .A2(\A2/A1/A2/A1/M3/c2 ),
    .ZN(\A2/A1/A2/A1/c3 ));
 AND2_X1 \A2/A1/A2/A1/M4/M1/_0_  (.A1(s1[11]),
    .A2(v1[27]),
    .ZN(\A2/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A2/A1/A2/A1/M4/M1/_1_  (.A(s1[11]),
    .B(v1[27]),
    .Z(\A2/A1/A2/A1/M4/s1 ));
 AND2_X1 \A2/A1/A2/A1/M4/M2/_0_  (.A1(\A2/A1/A2/A1/M4/s1 ),
    .A2(\A2/A1/A2/A1/c3 ),
    .ZN(\A2/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A2/A1/A2/A1/M4/M2/_1_  (.A(\A2/A1/A2/A1/M4/s1 ),
    .B(\A2/A1/A2/A1/c3 ),
    .Z(s2[11]));
 OR2_X1 \A2/A1/A2/A1/M4/_0_  (.A1(\A2/A1/A2/A1/M4/c1 ),
    .A2(\A2/A1/A2/A1/M4/c2 ),
    .ZN(\A2/A1/A2/c1 ));
 AND2_X1 \A2/A1/A2/A2/M1/M1/_0_  (.A1(s1[12]),
    .A2(v1[28]),
    .ZN(\A2/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M1/M1/_1_  (.A(s1[12]),
    .B(v1[28]),
    .Z(\A2/A1/A2/A2/M1/s1 ));
 AND2_X1 \A2/A1/A2/A2/M1/M2/_0_  (.A1(\A2/A1/A2/A2/M1/s1 ),
    .A2(\A2/A1/A2/c1 ),
    .ZN(\A2/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M1/M2/_1_  (.A(\A2/A1/A2/A2/M1/s1 ),
    .B(\A2/A1/A2/c1 ),
    .Z(s2[12]));
 OR2_X1 \A2/A1/A2/A2/M1/_0_  (.A1(\A2/A1/A2/A2/M1/c1 ),
    .A2(\A2/A1/A2/A2/M1/c2 ),
    .ZN(\A2/A1/A2/A2/c1 ));
 AND2_X1 \A2/A1/A2/A2/M2/M1/_0_  (.A1(s1[13]),
    .A2(v1[29]),
    .ZN(\A2/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M2/M1/_1_  (.A(s1[13]),
    .B(v1[29]),
    .Z(\A2/A1/A2/A2/M2/s1 ));
 AND2_X1 \A2/A1/A2/A2/M2/M2/_0_  (.A1(\A2/A1/A2/A2/M2/s1 ),
    .A2(\A2/A1/A2/A2/c1 ),
    .ZN(\A2/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M2/M2/_1_  (.A(\A2/A1/A2/A2/M2/s1 ),
    .B(\A2/A1/A2/A2/c1 ),
    .Z(s2[13]));
 OR2_X1 \A2/A1/A2/A2/M2/_0_  (.A1(\A2/A1/A2/A2/M2/c1 ),
    .A2(\A2/A1/A2/A2/M2/c2 ),
    .ZN(\A2/A1/A2/A2/c2 ));
 AND2_X1 \A2/A1/A2/A2/M3/M1/_0_  (.A1(s1[14]),
    .A2(v1[30]),
    .ZN(\A2/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M3/M1/_1_  (.A(s1[14]),
    .B(v1[30]),
    .Z(\A2/A1/A2/A2/M3/s1 ));
 AND2_X1 \A2/A1/A2/A2/M3/M2/_0_  (.A1(\A2/A1/A2/A2/M3/s1 ),
    .A2(\A2/A1/A2/A2/c2 ),
    .ZN(\A2/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M3/M2/_1_  (.A(\A2/A1/A2/A2/M3/s1 ),
    .B(\A2/A1/A2/A2/c2 ),
    .Z(s2[14]));
 OR2_X1 \A2/A1/A2/A2/M3/_0_  (.A1(\A2/A1/A2/A2/M3/c1 ),
    .A2(\A2/A1/A2/A2/M3/c2 ),
    .ZN(\A2/A1/A2/A2/c3 ));
 AND2_X1 \A2/A1/A2/A2/M4/M1/_0_  (.A1(s1[15]),
    .A2(v1[31]),
    .ZN(\A2/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A2/A1/A2/A2/M4/M1/_1_  (.A(s1[15]),
    .B(v1[31]),
    .Z(\A2/A1/A2/A2/M4/s1 ));
 AND2_X1 \A2/A1/A2/A2/M4/M2/_0_  (.A1(\A2/A1/A2/A2/M4/s1 ),
    .A2(\A2/A1/A2/A2/c3 ),
    .ZN(\A2/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A2/A1/A2/A2/M4/M2/_1_  (.A(\A2/A1/A2/A2/M4/s1 ),
    .B(\A2/A1/A2/A2/c3 ),
    .Z(s2[15]));
 OR2_X1 \A2/A1/A2/A2/M4/_0_  (.A1(\A2/A1/A2/A2/M4/c1 ),
    .A2(\A2/A1/A2/A2/M4/c2 ),
    .ZN(\A2/c1 ));
 AND2_X1 \A2/A2/A1/A1/M1/M1/_0_  (.A1(s1[16]),
    .A2(net2),
    .ZN(\A2/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M1/M1/_1_  (.A(s1[16]),
    .B(net2),
    .Z(\A2/A2/A1/A1/M1/s1 ));
 AND2_X1 \A2/A2/A1/A1/M1/M2/_0_  (.A1(\A2/A2/A1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\A2/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M1/M2/_1_  (.A(\A2/A2/A1/A1/M1/s1 ),
    .B(net2),
    .Z(s2[16]));
 OR2_X1 \A2/A2/A1/A1/M1/_0_  (.A1(\A2/A2/A1/A1/M1/c1 ),
    .A2(\A2/A2/A1/A1/M1/c2 ),
    .ZN(\A2/A2/A1/A1/c1 ));
 AND2_X1 \A2/A2/A1/A1/M2/M1/_0_  (.A1(s1[17]),
    .A2(net2),
    .ZN(\A2/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M2/M1/_1_  (.A(s1[17]),
    .B(net2),
    .Z(\A2/A2/A1/A1/M2/s1 ));
 AND2_X1 \A2/A2/A1/A1/M2/M2/_0_  (.A1(\A2/A2/A1/A1/M2/s1 ),
    .A2(\A2/A2/A1/A1/c1 ),
    .ZN(\A2/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M2/M2/_1_  (.A(\A2/A2/A1/A1/M2/s1 ),
    .B(\A2/A2/A1/A1/c1 ),
    .Z(s2[17]));
 OR2_X1 \A2/A2/A1/A1/M2/_0_  (.A1(\A2/A2/A1/A1/M2/c1 ),
    .A2(\A2/A2/A1/A1/M2/c2 ),
    .ZN(\A2/A2/A1/A1/c2 ));
 AND2_X1 \A2/A2/A1/A1/M3/M1/_0_  (.A1(s1[18]),
    .A2(net7),
    .ZN(\A2/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M3/M1/_1_  (.A(s1[18]),
    .B(net2),
    .Z(\A2/A2/A1/A1/M3/s1 ));
 AND2_X1 \A2/A2/A1/A1/M3/M2/_0_  (.A1(\A2/A2/A1/A1/M3/s1 ),
    .A2(\A2/A2/A1/A1/c2 ),
    .ZN(\A2/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M3/M2/_1_  (.A(\A2/A2/A1/A1/M3/s1 ),
    .B(\A2/A2/A1/A1/c2 ),
    .Z(s2[18]));
 OR2_X1 \A2/A2/A1/A1/M3/_0_  (.A1(\A2/A2/A1/A1/M3/c1 ),
    .A2(\A2/A2/A1/A1/M3/c2 ),
    .ZN(\A2/A2/A1/A1/c3 ));
 AND2_X1 \A2/A2/A1/A1/M4/M1/_0_  (.A1(s1[19]),
    .A2(net9),
    .ZN(\A2/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A2/A2/A1/A1/M4/M1/_1_  (.A(s1[19]),
    .B(net9),
    .Z(\A2/A2/A1/A1/M4/s1 ));
 AND2_X1 \A2/A2/A1/A1/M4/M2/_0_  (.A1(\A2/A2/A1/A1/M4/s1 ),
    .A2(\A2/A2/A1/A1/c3 ),
    .ZN(\A2/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A2/A2/A1/A1/M4/M2/_1_  (.A(\A2/A2/A1/A1/M4/s1 ),
    .B(\A2/A2/A1/A1/c3 ),
    .Z(s2[19]));
 OR2_X1 \A2/A2/A1/A1/M4/_0_  (.A1(\A2/A2/A1/A1/M4/c1 ),
    .A2(\A2/A2/A1/A1/M4/c2 ),
    .ZN(\A2/A2/A1/c1 ));
 AND2_X1 \A2/A2/A1/A2/M1/M1/_0_  (.A1(s1[20]),
    .A2(net9),
    .ZN(\A2/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M1/M1/_1_  (.A(s1[20]),
    .B(net9),
    .Z(\A2/A2/A1/A2/M1/s1 ));
 AND2_X1 \A2/A2/A1/A2/M1/M2/_0_  (.A1(\A2/A2/A1/A2/M1/s1 ),
    .A2(\A2/A2/A1/c1 ),
    .ZN(\A2/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M1/M2/_1_  (.A(\A2/A2/A1/A2/M1/s1 ),
    .B(\A2/A2/A1/c1 ),
    .Z(s2[20]));
 OR2_X1 \A2/A2/A1/A2/M1/_0_  (.A1(\A2/A2/A1/A2/M1/c1 ),
    .A2(\A2/A2/A1/A2/M1/c2 ),
    .ZN(\A2/A2/A1/A2/c1 ));
 AND2_X1 \A2/A2/A1/A2/M2/M1/_0_  (.A1(s1[21]),
    .A2(net9),
    .ZN(\A2/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M2/M1/_1_  (.A(s1[21]),
    .B(net9),
    .Z(\A2/A2/A1/A2/M2/s1 ));
 AND2_X1 \A2/A2/A1/A2/M2/M2/_0_  (.A1(\A2/A2/A1/A2/M2/s1 ),
    .A2(\A2/A2/A1/A2/c1 ),
    .ZN(\A2/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M2/M2/_1_  (.A(\A2/A2/A1/A2/M2/s1 ),
    .B(\A2/A2/A1/A2/c1 ),
    .Z(s2[21]));
 OR2_X1 \A2/A2/A1/A2/M2/_0_  (.A1(\A2/A2/A1/A2/M2/c1 ),
    .A2(\A2/A2/A1/A2/M2/c2 ),
    .ZN(\A2/A2/A1/A2/c2 ));
 AND2_X1 \A2/A2/A1/A2/M3/M1/_0_  (.A1(s1[22]),
    .A2(net9),
    .ZN(\A2/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M3/M1/_1_  (.A(s1[22]),
    .B(net9),
    .Z(\A2/A2/A1/A2/M3/s1 ));
 AND2_X1 \A2/A2/A1/A2/M3/M2/_0_  (.A1(\A2/A2/A1/A2/M3/s1 ),
    .A2(\A2/A2/A1/A2/c2 ),
    .ZN(\A2/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M3/M2/_1_  (.A(\A2/A2/A1/A2/M3/s1 ),
    .B(\A2/A2/A1/A2/c2 ),
    .Z(s2[22]));
 OR2_X1 \A2/A2/A1/A2/M3/_0_  (.A1(\A2/A2/A1/A2/M3/c1 ),
    .A2(\A2/A2/A1/A2/M3/c2 ),
    .ZN(\A2/A2/A1/A2/c3 ));
 AND2_X1 \A2/A2/A1/A2/M4/M1/_0_  (.A1(s1[23]),
    .A2(net9),
    .ZN(\A2/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A2/A2/A1/A2/M4/M1/_1_  (.A(s1[23]),
    .B(net9),
    .Z(\A2/A2/A1/A2/M4/s1 ));
 AND2_X1 \A2/A2/A1/A2/M4/M2/_0_  (.A1(\A2/A2/A1/A2/M4/s1 ),
    .A2(\A2/A2/A1/A2/c3 ),
    .ZN(\A2/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A2/A2/A1/A2/M4/M2/_1_  (.A(\A2/A2/A1/A2/M4/s1 ),
    .B(\A2/A2/A1/A2/c3 ),
    .Z(s2[23]));
 OR2_X1 \A2/A2/A1/A2/M4/_0_  (.A1(\A2/A2/A1/A2/M4/c1 ),
    .A2(\A2/A2/A1/A2/M4/c2 ),
    .ZN(\A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A1/M1/M1/_0_  (.A1(s1[24]),
    .A2(net9),
    .ZN(\A2/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M1/M1/_1_  (.A(s1[24]),
    .B(net9),
    .Z(\A2/A2/A2/A1/M1/s1 ));
 AND2_X1 \A2/A2/A2/A1/M1/M2/_0_  (.A1(\A2/A2/A2/A1/M1/s1 ),
    .A2(\A2/A2/c1 ),
    .ZN(\A2/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M1/M2/_1_  (.A(\A2/A2/A2/A1/M1/s1 ),
    .B(\A2/A2/c1 ),
    .Z(s2[24]));
 OR2_X1 \A2/A2/A2/A1/M1/_0_  (.A1(\A2/A2/A2/A1/M1/c1 ),
    .A2(\A2/A2/A2/A1/M1/c2 ),
    .ZN(\A2/A2/A2/A1/c1 ));
 AND2_X1 \A2/A2/A2/A1/M2/M1/_0_  (.A1(s1[25]),
    .A2(net9),
    .ZN(\A2/A2/A2/A1/M2/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M2/M1/_1_  (.A(s1[25]),
    .B(net9),
    .Z(\A2/A2/A2/A1/M2/s1 ));
 AND2_X1 \A2/A2/A2/A1/M2/M2/_0_  (.A1(\A2/A2/A2/A1/M2/s1 ),
    .A2(\A2/A2/A2/A1/c1 ),
    .ZN(\A2/A2/A2/A1/M2/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M2/M2/_1_  (.A(\A2/A2/A2/A1/M2/s1 ),
    .B(\A2/A2/A2/A1/c1 ),
    .Z(s2[25]));
 OR2_X1 \A2/A2/A2/A1/M2/_0_  (.A1(\A2/A2/A2/A1/M2/c1 ),
    .A2(\A2/A2/A2/A1/M2/c2 ),
    .ZN(\A2/A2/A2/A1/c2 ));
 AND2_X1 \A2/A2/A2/A1/M3/M1/_0_  (.A1(s1[26]),
    .A2(net9),
    .ZN(\A2/A2/A2/A1/M3/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M3/M1/_1_  (.A(s1[26]),
    .B(net9),
    .Z(\A2/A2/A2/A1/M3/s1 ));
 AND2_X1 \A2/A2/A2/A1/M3/M2/_0_  (.A1(\A2/A2/A2/A1/M3/s1 ),
    .A2(\A2/A2/A2/A1/c2 ),
    .ZN(\A2/A2/A2/A1/M3/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M3/M2/_1_  (.A(\A2/A2/A2/A1/M3/s1 ),
    .B(\A2/A2/A2/A1/c2 ),
    .Z(s2[26]));
 OR2_X1 \A2/A2/A2/A1/M3/_0_  (.A1(\A2/A2/A2/A1/M3/c1 ),
    .A2(\A2/A2/A2/A1/M3/c2 ),
    .ZN(\A2/A2/A2/A1/c3 ));
 AND2_X1 \A2/A2/A2/A1/M4/M1/_0_  (.A1(s1[27]),
    .A2(net9),
    .ZN(\A2/A2/A2/A1/M4/c1 ));
 XOR2_X2 \A2/A2/A2/A1/M4/M1/_1_  (.A(s1[27]),
    .B(net9),
    .Z(\A2/A2/A2/A1/M4/s1 ));
 AND2_X1 \A2/A2/A2/A1/M4/M2/_0_  (.A1(\A2/A2/A2/A1/M4/s1 ),
    .A2(\A2/A2/A2/A1/c3 ),
    .ZN(\A2/A2/A2/A1/M4/c2 ));
 XOR2_X2 \A2/A2/A2/A1/M4/M2/_1_  (.A(\A2/A2/A2/A1/M4/s1 ),
    .B(\A2/A2/A2/A1/c3 ),
    .Z(s2[27]));
 OR2_X1 \A2/A2/A2/A1/M4/_0_  (.A1(\A2/A2/A2/A1/M4/c1 ),
    .A2(\A2/A2/A2/A1/M4/c2 ),
    .ZN(\A2/A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A2/M1/M1/_0_  (.A1(s1[28]),
    .A2(net9),
    .ZN(\A2/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M1/M1/_1_  (.A(s1[28]),
    .B(net9),
    .Z(\A2/A2/A2/A2/M1/s1 ));
 AND2_X1 \A2/A2/A2/A2/M1/M2/_0_  (.A1(\A2/A2/A2/A2/M1/s1 ),
    .A2(\A2/A2/A2/c1 ),
    .ZN(\A2/A2/A2/A2/M1/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M1/M2/_1_  (.A(\A2/A2/A2/A2/M1/s1 ),
    .B(\A2/A2/A2/c1 ),
    .Z(s2[28]));
 OR2_X1 \A2/A2/A2/A2/M1/_0_  (.A1(\A2/A2/A2/A2/M1/c1 ),
    .A2(\A2/A2/A2/A2/M1/c2 ),
    .ZN(\A2/A2/A2/A2/c1 ));
 AND2_X1 \A2/A2/A2/A2/M2/M1/_0_  (.A1(s1[29]),
    .A2(net9),
    .ZN(\A2/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M2/M1/_1_  (.A(s1[29]),
    .B(net9),
    .Z(\A2/A2/A2/A2/M2/s1 ));
 AND2_X1 \A2/A2/A2/A2/M2/M2/_0_  (.A1(\A2/A2/A2/A2/M2/s1 ),
    .A2(\A2/A2/A2/A2/c1 ),
    .ZN(\A2/A2/A2/A2/M2/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M2/M2/_1_  (.A(\A2/A2/A2/A2/M2/s1 ),
    .B(\A2/A2/A2/A2/c1 ),
    .Z(s2[29]));
 OR2_X1 \A2/A2/A2/A2/M2/_0_  (.A1(\A2/A2/A2/A2/M2/c1 ),
    .A2(\A2/A2/A2/A2/M2/c2 ),
    .ZN(\A2/A2/A2/A2/c2 ));
 AND2_X1 \A2/A2/A2/A2/M3/M1/_0_  (.A1(s1[30]),
    .A2(net9),
    .ZN(\A2/A2/A2/A2/M3/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M3/M1/_1_  (.A(s1[30]),
    .B(net9),
    .Z(\A2/A2/A2/A2/M3/s1 ));
 AND2_X1 \A2/A2/A2/A2/M3/M2/_0_  (.A1(\A2/A2/A2/A2/M3/s1 ),
    .A2(\A2/A2/A2/A2/c2 ),
    .ZN(\A2/A2/A2/A2/M3/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M3/M2/_1_  (.A(\A2/A2/A2/A2/M3/s1 ),
    .B(\A2/A2/A2/A2/c2 ),
    .Z(s2[30]));
 OR2_X1 \A2/A2/A2/A2/M3/_0_  (.A1(\A2/A2/A2/A2/M3/c1 ),
    .A2(\A2/A2/A2/A2/M3/c2 ),
    .ZN(\A2/A2/A2/A2/c3 ));
 AND2_X1 \A2/A2/A2/A2/M4/M1/_0_  (.A1(s1[31]),
    .A2(net9),
    .ZN(\A2/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A2/A2/A2/A2/M4/M1/_1_  (.A(s1[31]),
    .B(net9),
    .Z(\A2/A2/A2/A2/M4/s1 ));
 AND2_X1 \A2/A2/A2/A2/M4/M2/_0_  (.A1(\A2/A2/A2/A2/M4/s1 ),
    .A2(\A2/A2/A2/A2/c3 ),
    .ZN(\A2/A2/A2/A2/M4/c2 ));
 XOR2_X2 \A2/A2/A2/A2/M4/M2/_1_  (.A(\A2/A2/A2/A2/M4/s1 ),
    .B(\A2/A2/A2/A2/c3 ),
    .Z(s2[31]));
 OR2_X1 \A2/A2/A2/A2/M4/_0_  (.A1(\A2/A2/A2/A2/M4/c1 ),
    .A2(\A2/A2/A2/A2/M4/c2 ),
    .ZN(c2));
 AND2_X1 \A3/A1/A1/A1/M1/M1/_0_  (.A1(v4[0]),
    .A2(s2[16]),
    .ZN(\A3/A1/A1/A1/M1/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M1/M1/_1_  (.A(v4[0]),
    .B(s2[16]),
    .Z(\A3/A1/A1/A1/M1/s1 ));
 AND2_X1 \A3/A1/A1/A1/M1/M2/_0_  (.A1(\A3/A1/A1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\A3/A1/A1/A1/M1/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M1/M2/_1_  (.A(\A3/A1/A1/A1/M1/s1 ),
    .B(net2),
    .Z(Prod[32]));
 OR2_X1 \A3/A1/A1/A1/M1/_0_  (.A1(\A3/A1/A1/A1/M1/c1 ),
    .A2(\A3/A1/A1/A1/M1/c2 ),
    .ZN(\A3/A1/A1/A1/c1 ));
 AND2_X1 \A3/A1/A1/A1/M2/M1/_0_  (.A1(v4[1]),
    .A2(s2[17]),
    .ZN(\A3/A1/A1/A1/M2/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M2/M1/_1_  (.A(v4[1]),
    .B(s2[17]),
    .Z(\A3/A1/A1/A1/M2/s1 ));
 AND2_X1 \A3/A1/A1/A1/M2/M2/_0_  (.A1(\A3/A1/A1/A1/M2/s1 ),
    .A2(\A3/A1/A1/A1/c1 ),
    .ZN(\A3/A1/A1/A1/M2/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M2/M2/_1_  (.A(\A3/A1/A1/A1/M2/s1 ),
    .B(\A3/A1/A1/A1/c1 ),
    .Z(Prod[33]));
 OR2_X1 \A3/A1/A1/A1/M2/_0_  (.A1(\A3/A1/A1/A1/M2/c1 ),
    .A2(\A3/A1/A1/A1/M2/c2 ),
    .ZN(\A3/A1/A1/A1/c2 ));
 AND2_X1 \A3/A1/A1/A1/M3/M1/_0_  (.A1(v4[2]),
    .A2(s2[18]),
    .ZN(\A3/A1/A1/A1/M3/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M3/M1/_1_  (.A(v4[2]),
    .B(s2[18]),
    .Z(\A3/A1/A1/A1/M3/s1 ));
 AND2_X1 \A3/A1/A1/A1/M3/M2/_0_  (.A1(\A3/A1/A1/A1/M3/s1 ),
    .A2(\A3/A1/A1/A1/c2 ),
    .ZN(\A3/A1/A1/A1/M3/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M3/M2/_1_  (.A(\A3/A1/A1/A1/M3/s1 ),
    .B(\A3/A1/A1/A1/c2 ),
    .Z(Prod[34]));
 OR2_X1 \A3/A1/A1/A1/M3/_0_  (.A1(\A3/A1/A1/A1/M3/c1 ),
    .A2(\A3/A1/A1/A1/M3/c2 ),
    .ZN(\A3/A1/A1/A1/c3 ));
 AND2_X1 \A3/A1/A1/A1/M4/M1/_0_  (.A1(v4[3]),
    .A2(s2[19]),
    .ZN(\A3/A1/A1/A1/M4/c1 ));
 XOR2_X2 \A3/A1/A1/A1/M4/M1/_1_  (.A(v4[3]),
    .B(s2[19]),
    .Z(\A3/A1/A1/A1/M4/s1 ));
 AND2_X1 \A3/A1/A1/A1/M4/M2/_0_  (.A1(\A3/A1/A1/A1/M4/s1 ),
    .A2(\A3/A1/A1/A1/c3 ),
    .ZN(\A3/A1/A1/A1/M4/c2 ));
 XOR2_X2 \A3/A1/A1/A1/M4/M2/_1_  (.A(\A3/A1/A1/A1/M4/s1 ),
    .B(\A3/A1/A1/A1/c3 ),
    .Z(Prod[35]));
 OR2_X1 \A3/A1/A1/A1/M4/_0_  (.A1(\A3/A1/A1/A1/M4/c1 ),
    .A2(\A3/A1/A1/A1/M4/c2 ),
    .ZN(\A3/A1/A1/c1 ));
 AND2_X1 \A3/A1/A1/A2/M1/M1/_0_  (.A1(v4[4]),
    .A2(s2[20]),
    .ZN(\A3/A1/A1/A2/M1/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M1/M1/_1_  (.A(v4[4]),
    .B(s2[20]),
    .Z(\A3/A1/A1/A2/M1/s1 ));
 AND2_X1 \A3/A1/A1/A2/M1/M2/_0_  (.A1(\A3/A1/A1/A2/M1/s1 ),
    .A2(\A3/A1/A1/c1 ),
    .ZN(\A3/A1/A1/A2/M1/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M1/M2/_1_  (.A(\A3/A1/A1/A2/M1/s1 ),
    .B(\A3/A1/A1/c1 ),
    .Z(Prod[36]));
 OR2_X1 \A3/A1/A1/A2/M1/_0_  (.A1(\A3/A1/A1/A2/M1/c1 ),
    .A2(\A3/A1/A1/A2/M1/c2 ),
    .ZN(\A3/A1/A1/A2/c1 ));
 AND2_X1 \A3/A1/A1/A2/M2/M1/_0_  (.A1(v4[5]),
    .A2(s2[21]),
    .ZN(\A3/A1/A1/A2/M2/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M2/M1/_1_  (.A(v4[5]),
    .B(s2[21]),
    .Z(\A3/A1/A1/A2/M2/s1 ));
 AND2_X1 \A3/A1/A1/A2/M2/M2/_0_  (.A1(\A3/A1/A1/A2/M2/s1 ),
    .A2(\A3/A1/A1/A2/c1 ),
    .ZN(\A3/A1/A1/A2/M2/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M2/M2/_1_  (.A(\A3/A1/A1/A2/M2/s1 ),
    .B(\A3/A1/A1/A2/c1 ),
    .Z(Prod[37]));
 OR2_X1 \A3/A1/A1/A2/M2/_0_  (.A1(\A3/A1/A1/A2/M2/c1 ),
    .A2(\A3/A1/A1/A2/M2/c2 ),
    .ZN(\A3/A1/A1/A2/c2 ));
 AND2_X1 \A3/A1/A1/A2/M3/M1/_0_  (.A1(v4[6]),
    .A2(s2[22]),
    .ZN(\A3/A1/A1/A2/M3/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M3/M1/_1_  (.A(v4[6]),
    .B(s2[22]),
    .Z(\A3/A1/A1/A2/M3/s1 ));
 AND2_X1 \A3/A1/A1/A2/M3/M2/_0_  (.A1(\A3/A1/A1/A2/M3/s1 ),
    .A2(\A3/A1/A1/A2/c2 ),
    .ZN(\A3/A1/A1/A2/M3/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M3/M2/_1_  (.A(\A3/A1/A1/A2/M3/s1 ),
    .B(\A3/A1/A1/A2/c2 ),
    .Z(Prod[38]));
 OR2_X1 \A3/A1/A1/A2/M3/_0_  (.A1(\A3/A1/A1/A2/M3/c1 ),
    .A2(\A3/A1/A1/A2/M3/c2 ),
    .ZN(\A3/A1/A1/A2/c3 ));
 AND2_X1 \A3/A1/A1/A2/M4/M1/_0_  (.A1(v4[7]),
    .A2(s2[23]),
    .ZN(\A3/A1/A1/A2/M4/c1 ));
 XOR2_X2 \A3/A1/A1/A2/M4/M1/_1_  (.A(v4[7]),
    .B(s2[23]),
    .Z(\A3/A1/A1/A2/M4/s1 ));
 AND2_X1 \A3/A1/A1/A2/M4/M2/_0_  (.A1(\A3/A1/A1/A2/M4/s1 ),
    .A2(\A3/A1/A1/A2/c3 ),
    .ZN(\A3/A1/A1/A2/M4/c2 ));
 XOR2_X2 \A3/A1/A1/A2/M4/M2/_1_  (.A(\A3/A1/A1/A2/M4/s1 ),
    .B(\A3/A1/A1/A2/c3 ),
    .Z(Prod[39]));
 OR2_X1 \A3/A1/A1/A2/M4/_0_  (.A1(\A3/A1/A1/A2/M4/c1 ),
    .A2(\A3/A1/A1/A2/M4/c2 ),
    .ZN(\A3/A1/c1 ));
 AND2_X1 \A3/A1/A2/A1/M1/M1/_0_  (.A1(v4[8]),
    .A2(s2[24]),
    .ZN(\A3/A1/A2/A1/M1/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M1/M1/_1_  (.A(v4[8]),
    .B(s2[24]),
    .Z(\A3/A1/A2/A1/M1/s1 ));
 AND2_X1 \A3/A1/A2/A1/M1/M2/_0_  (.A1(\A3/A1/A2/A1/M1/s1 ),
    .A2(\A3/A1/c1 ),
    .ZN(\A3/A1/A2/A1/M1/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M1/M2/_1_  (.A(\A3/A1/A2/A1/M1/s1 ),
    .B(\A3/A1/c1 ),
    .Z(Prod[40]));
 OR2_X1 \A3/A1/A2/A1/M1/_0_  (.A1(\A3/A1/A2/A1/M1/c1 ),
    .A2(\A3/A1/A2/A1/M1/c2 ),
    .ZN(\A3/A1/A2/A1/c1 ));
 AND2_X1 \A3/A1/A2/A1/M2/M1/_0_  (.A1(v4[9]),
    .A2(s2[25]),
    .ZN(\A3/A1/A2/A1/M2/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M2/M1/_1_  (.A(v4[9]),
    .B(s2[25]),
    .Z(\A3/A1/A2/A1/M2/s1 ));
 AND2_X1 \A3/A1/A2/A1/M2/M2/_0_  (.A1(\A3/A1/A2/A1/M2/s1 ),
    .A2(\A3/A1/A2/A1/c1 ),
    .ZN(\A3/A1/A2/A1/M2/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M2/M2/_1_  (.A(\A3/A1/A2/A1/M2/s1 ),
    .B(\A3/A1/A2/A1/c1 ),
    .Z(Prod[41]));
 OR2_X1 \A3/A1/A2/A1/M2/_0_  (.A1(\A3/A1/A2/A1/M2/c1 ),
    .A2(\A3/A1/A2/A1/M2/c2 ),
    .ZN(\A3/A1/A2/A1/c2 ));
 AND2_X1 \A3/A1/A2/A1/M3/M1/_0_  (.A1(v4[10]),
    .A2(s2[26]),
    .ZN(\A3/A1/A2/A1/M3/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M3/M1/_1_  (.A(v4[10]),
    .B(s2[26]),
    .Z(\A3/A1/A2/A1/M3/s1 ));
 AND2_X1 \A3/A1/A2/A1/M3/M2/_0_  (.A1(\A3/A1/A2/A1/M3/s1 ),
    .A2(\A3/A1/A2/A1/c2 ),
    .ZN(\A3/A1/A2/A1/M3/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M3/M2/_1_  (.A(\A3/A1/A2/A1/M3/s1 ),
    .B(\A3/A1/A2/A1/c2 ),
    .Z(Prod[42]));
 OR2_X1 \A3/A1/A2/A1/M3/_0_  (.A1(\A3/A1/A2/A1/M3/c1 ),
    .A2(\A3/A1/A2/A1/M3/c2 ),
    .ZN(\A3/A1/A2/A1/c3 ));
 AND2_X1 \A3/A1/A2/A1/M4/M1/_0_  (.A1(v4[11]),
    .A2(s2[27]),
    .ZN(\A3/A1/A2/A1/M4/c1 ));
 XOR2_X2 \A3/A1/A2/A1/M4/M1/_1_  (.A(v4[11]),
    .B(s2[27]),
    .Z(\A3/A1/A2/A1/M4/s1 ));
 AND2_X1 \A3/A1/A2/A1/M4/M2/_0_  (.A1(\A3/A1/A2/A1/M4/s1 ),
    .A2(\A3/A1/A2/A1/c3 ),
    .ZN(\A3/A1/A2/A1/M4/c2 ));
 XOR2_X2 \A3/A1/A2/A1/M4/M2/_1_  (.A(\A3/A1/A2/A1/M4/s1 ),
    .B(\A3/A1/A2/A1/c3 ),
    .Z(Prod[43]));
 OR2_X1 \A3/A1/A2/A1/M4/_0_  (.A1(\A3/A1/A2/A1/M4/c1 ),
    .A2(\A3/A1/A2/A1/M4/c2 ),
    .ZN(\A3/A1/A2/c1 ));
 AND2_X1 \A3/A1/A2/A2/M1/M1/_0_  (.A1(v4[12]),
    .A2(s2[28]),
    .ZN(\A3/A1/A2/A2/M1/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M1/M1/_1_  (.A(v4[12]),
    .B(s2[28]),
    .Z(\A3/A1/A2/A2/M1/s1 ));
 AND2_X1 \A3/A1/A2/A2/M1/M2/_0_  (.A1(\A3/A1/A2/A2/M1/s1 ),
    .A2(\A3/A1/A2/c1 ),
    .ZN(\A3/A1/A2/A2/M1/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M1/M2/_1_  (.A(\A3/A1/A2/A2/M1/s1 ),
    .B(\A3/A1/A2/c1 ),
    .Z(Prod[44]));
 OR2_X1 \A3/A1/A2/A2/M1/_0_  (.A1(\A3/A1/A2/A2/M1/c1 ),
    .A2(\A3/A1/A2/A2/M1/c2 ),
    .ZN(\A3/A1/A2/A2/c1 ));
 AND2_X1 \A3/A1/A2/A2/M2/M1/_0_  (.A1(v4[13]),
    .A2(s2[29]),
    .ZN(\A3/A1/A2/A2/M2/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M2/M1/_1_  (.A(v4[13]),
    .B(s2[29]),
    .Z(\A3/A1/A2/A2/M2/s1 ));
 AND2_X1 \A3/A1/A2/A2/M2/M2/_0_  (.A1(\A3/A1/A2/A2/M2/s1 ),
    .A2(\A3/A1/A2/A2/c1 ),
    .ZN(\A3/A1/A2/A2/M2/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M2/M2/_1_  (.A(\A3/A1/A2/A2/M2/s1 ),
    .B(\A3/A1/A2/A2/c1 ),
    .Z(Prod[45]));
 OR2_X1 \A3/A1/A2/A2/M2/_0_  (.A1(\A3/A1/A2/A2/M2/c1 ),
    .A2(\A3/A1/A2/A2/M2/c2 ),
    .ZN(\A3/A1/A2/A2/c2 ));
 AND2_X1 \A3/A1/A2/A2/M3/M1/_0_  (.A1(v4[14]),
    .A2(s2[30]),
    .ZN(\A3/A1/A2/A2/M3/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M3/M1/_1_  (.A(v4[14]),
    .B(s2[30]),
    .Z(\A3/A1/A2/A2/M3/s1 ));
 AND2_X1 \A3/A1/A2/A2/M3/M2/_0_  (.A1(\A3/A1/A2/A2/M3/s1 ),
    .A2(\A3/A1/A2/A2/c2 ),
    .ZN(\A3/A1/A2/A2/M3/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M3/M2/_1_  (.A(\A3/A1/A2/A2/M3/s1 ),
    .B(\A3/A1/A2/A2/c2 ),
    .Z(Prod[46]));
 OR2_X1 \A3/A1/A2/A2/M3/_0_  (.A1(\A3/A1/A2/A2/M3/c1 ),
    .A2(\A3/A1/A2/A2/M3/c2 ),
    .ZN(\A3/A1/A2/A2/c3 ));
 AND2_X1 \A3/A1/A2/A2/M4/M1/_0_  (.A1(v4[15]),
    .A2(s2[31]),
    .ZN(\A3/A1/A2/A2/M4/c1 ));
 XOR2_X2 \A3/A1/A2/A2/M4/M1/_1_  (.A(v4[15]),
    .B(s2[31]),
    .Z(\A3/A1/A2/A2/M4/s1 ));
 AND2_X1 \A3/A1/A2/A2/M4/M2/_0_  (.A1(\A3/A1/A2/A2/M4/s1 ),
    .A2(\A3/A1/A2/A2/c3 ),
    .ZN(\A3/A1/A2/A2/M4/c2 ));
 XOR2_X2 \A3/A1/A2/A2/M4/M2/_1_  (.A(\A3/A1/A2/A2/M4/s1 ),
    .B(\A3/A1/A2/A2/c3 ),
    .Z(Prod[47]));
 OR2_X1 \A3/A1/A2/A2/M4/_0_  (.A1(\A3/A1/A2/A2/M4/c1 ),
    .A2(\A3/A1/A2/A2/M4/c2 ),
    .ZN(\A3/c1 ));
 AND2_X1 \A3/A2/A1/A1/M1/M1/_0_  (.A1(v4[16]),
    .A2(c3),
    .ZN(\A3/A2/A1/A1/M1/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M1/M1/_1_  (.A(v4[16]),
    .B(c3),
    .Z(\A3/A2/A1/A1/M1/s1 ));
 AND2_X1 \A3/A2/A1/A1/M1/M2/_0_  (.A1(\A3/A2/A1/A1/M1/s1 ),
    .A2(net1),
    .ZN(\A3/A2/A1/A1/M1/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M1/M2/_1_  (.A(\A3/A2/A1/A1/M1/s1 ),
    .B(net1),
    .Z(Prod[48]));
 OR2_X1 \A3/A2/A1/A1/M1/_0_  (.A1(\A3/A2/A1/A1/M1/c1 ),
    .A2(\A3/A2/A1/A1/M1/c2 ),
    .ZN(\A3/A2/A1/A1/c1 ));
 AND2_X1 \A3/A2/A1/A1/M2/M1/_0_  (.A1(v4[17]),
    .A2(net1),
    .ZN(\A3/A2/A1/A1/M2/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M2/M1/_1_  (.A(v4[17]),
    .B(net1),
    .Z(\A3/A2/A1/A1/M2/s1 ));
 AND2_X1 \A3/A2/A1/A1/M2/M2/_0_  (.A1(\A3/A2/A1/A1/M2/s1 ),
    .A2(\A3/A2/A1/A1/c1 ),
    .ZN(\A3/A2/A1/A1/M2/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M2/M2/_1_  (.A(\A3/A2/A1/A1/M2/s1 ),
    .B(\A3/A2/A1/A1/c1 ),
    .Z(Prod[49]));
 OR2_X1 \A3/A2/A1/A1/M2/_0_  (.A1(\A3/A2/A1/A1/M2/c1 ),
    .A2(\A3/A2/A1/A1/M2/c2 ),
    .ZN(\A3/A2/A1/A1/c2 ));
 AND2_X1 \A3/A2/A1/A1/M3/M1/_0_  (.A1(v4[18]),
    .A2(net1),
    .ZN(\A3/A2/A1/A1/M3/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M3/M1/_1_  (.A(v4[18]),
    .B(net1),
    .Z(\A3/A2/A1/A1/M3/s1 ));
 AND2_X1 \A3/A2/A1/A1/M3/M2/_0_  (.A1(\A3/A2/A1/A1/M3/s1 ),
    .A2(\A3/A2/A1/A1/c2 ),
    .ZN(\A3/A2/A1/A1/M3/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M3/M2/_1_  (.A(\A3/A2/A1/A1/M3/s1 ),
    .B(\A3/A2/A1/A1/c2 ),
    .Z(Prod[50]));
 OR2_X1 \A3/A2/A1/A1/M3/_0_  (.A1(\A3/A2/A1/A1/M3/c1 ),
    .A2(\A3/A2/A1/A1/M3/c2 ),
    .ZN(\A3/A2/A1/A1/c3 ));
 AND2_X1 \A3/A2/A1/A1/M4/M1/_0_  (.A1(v4[19]),
    .A2(net1),
    .ZN(\A3/A2/A1/A1/M4/c1 ));
 XOR2_X2 \A3/A2/A1/A1/M4/M1/_1_  (.A(v4[19]),
    .B(net1),
    .Z(\A3/A2/A1/A1/M4/s1 ));
 AND2_X1 \A3/A2/A1/A1/M4/M2/_0_  (.A1(\A3/A2/A1/A1/M4/s1 ),
    .A2(\A3/A2/A1/A1/c3 ),
    .ZN(\A3/A2/A1/A1/M4/c2 ));
 XOR2_X2 \A3/A2/A1/A1/M4/M2/_1_  (.A(\A3/A2/A1/A1/M4/s1 ),
    .B(\A3/A2/A1/A1/c3 ),
    .Z(Prod[51]));
 OR2_X1 \A3/A2/A1/A1/M4/_0_  (.A1(\A3/A2/A1/A1/M4/c1 ),
    .A2(\A3/A2/A1/A1/M4/c2 ),
    .ZN(\A3/A2/A1/c1 ));
 AND2_X1 \A3/A2/A1/A2/M1/M1/_0_  (.A1(v4[20]),
    .A2(net10),
    .ZN(\A3/A2/A1/A2/M1/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M1/M1/_1_  (.A(v4[20]),
    .B(net10),
    .Z(\A3/A2/A1/A2/M1/s1 ));
 AND2_X1 \A3/A2/A1/A2/M1/M2/_0_  (.A1(\A3/A2/A1/A2/M1/s1 ),
    .A2(\A3/A2/A1/c1 ),
    .ZN(\A3/A2/A1/A2/M1/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M1/M2/_1_  (.A(\A3/A2/A1/A2/M1/s1 ),
    .B(\A3/A2/A1/c1 ),
    .Z(Prod[52]));
 OR2_X1 \A3/A2/A1/A2/M1/_0_  (.A1(\A3/A2/A1/A2/M1/c1 ),
    .A2(\A3/A2/A1/A2/M1/c2 ),
    .ZN(\A3/A2/A1/A2/c1 ));
 AND2_X1 \A3/A2/A1/A2/M2/M1/_0_  (.A1(v4[21]),
    .A2(net10),
    .ZN(\A3/A2/A1/A2/M2/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M2/M1/_1_  (.A(v4[21]),
    .B(net10),
    .Z(\A3/A2/A1/A2/M2/s1 ));
 AND2_X1 \A3/A2/A1/A2/M2/M2/_0_  (.A1(\A3/A2/A1/A2/M2/s1 ),
    .A2(\A3/A2/A1/A2/c1 ),
    .ZN(\A3/A2/A1/A2/M2/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M2/M2/_1_  (.A(\A3/A2/A1/A2/M2/s1 ),
    .B(\A3/A2/A1/A2/c1 ),
    .Z(Prod[53]));
 OR2_X1 \A3/A2/A1/A2/M2/_0_  (.A1(\A3/A2/A1/A2/M2/c1 ),
    .A2(\A3/A2/A1/A2/M2/c2 ),
    .ZN(\A3/A2/A1/A2/c2 ));
 AND2_X1 \A3/A2/A1/A2/M3/M1/_0_  (.A1(v4[22]),
    .A2(net10),
    .ZN(\A3/A2/A1/A2/M3/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M3/M1/_1_  (.A(v4[22]),
    .B(net10),
    .Z(\A3/A2/A1/A2/M3/s1 ));
 AND2_X1 \A3/A2/A1/A2/M3/M2/_0_  (.A1(\A3/A2/A1/A2/M3/s1 ),
    .A2(\A3/A2/A1/A2/c2 ),
    .ZN(\A3/A2/A1/A2/M3/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M3/M2/_1_  (.A(\A3/A2/A1/A2/M3/s1 ),
    .B(\A3/A2/A1/A2/c2 ),
    .Z(Prod[54]));
 OR2_X1 \A3/A2/A1/A2/M3/_0_  (.A1(\A3/A2/A1/A2/M3/c1 ),
    .A2(\A3/A2/A1/A2/M3/c2 ),
    .ZN(\A3/A2/A1/A2/c3 ));
 AND2_X1 \A3/A2/A1/A2/M4/M1/_0_  (.A1(v4[23]),
    .A2(net10),
    .ZN(\A3/A2/A1/A2/M4/c1 ));
 XOR2_X2 \A3/A2/A1/A2/M4/M1/_1_  (.A(v4[23]),
    .B(net10),
    .Z(\A3/A2/A1/A2/M4/s1 ));
 AND2_X1 \A3/A2/A1/A2/M4/M2/_0_  (.A1(\A3/A2/A1/A2/M4/s1 ),
    .A2(\A3/A2/A1/A2/c3 ),
    .ZN(\A3/A2/A1/A2/M4/c2 ));
 XOR2_X2 \A3/A2/A1/A2/M4/M2/_1_  (.A(\A3/A2/A1/A2/M4/s1 ),
    .B(\A3/A2/A1/A2/c3 ),
    .Z(Prod[55]));
 OR2_X1 \A3/A2/A1/A2/M4/_0_  (.A1(\A3/A2/A1/A2/M4/c1 ),
    .A2(\A3/A2/A1/A2/M4/c2 ),
    .ZN(\A3/A2/c1 ));
 AND2_X1 \A3/A2/A2/A1/M1/M1/_0_  (.A1(v4[24]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M1/c1 ));
 XOR2_X2 \A3/A2/A2/A1/M1/M1/_1_  (.A(v4[24]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M1/s1 ));
 AND2_X1 \A3/A2/A2/A1/M1/M2/_0_  (.A1(\A3/A2/A2/A1/M1/s1 ),
    .A2(\A3/A2/c1 ),
    .ZN(\A3/A2/A2/A1/M1/c2 ));
 XOR2_X2 \A3/A2/A2/A1/M1/M2/_1_  (.A(\A3/A2/A2/A1/M1/s1 ),
    .B(\A3/A2/c1 ),
    .Z(Prod[56]));
 OR2_X1 \A3/A2/A2/A1/M1/_0_  (.A1(\A3/A2/A2/A1/M1/c1 ),
    .A2(\A3/A2/A2/A1/M1/c2 ),
    .ZN(\A3/A2/A2/A1/c1 ));
 AND2_X1 \A3/A2/A2/A1/M2/M1/_0_  (.A1(v4[25]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M2/c1 ));
 XOR2_X2 \A3/A2/A2/A1/M2/M1/_1_  (.A(v4[25]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M2/s1 ));
 AND2_X1 \A3/A2/A2/A1/M2/M2/_0_  (.A1(\A3/A2/A2/A1/M2/s1 ),
    .A2(\A3/A2/A2/A1/c1 ),
    .ZN(\A3/A2/A2/A1/M2/c2 ));
 XOR2_X2 \A3/A2/A2/A1/M2/M2/_1_  (.A(\A3/A2/A2/A1/M2/s1 ),
    .B(\A3/A2/A2/A1/c1 ),
    .Z(Prod[57]));
 OR2_X1 \A3/A2/A2/A1/M2/_0_  (.A1(\A3/A2/A2/A1/M2/c1 ),
    .A2(\A3/A2/A2/A1/M2/c2 ),
    .ZN(\A3/A2/A2/A1/c2 ));
 AND2_X1 \A3/A2/A2/A1/M3/M1/_0_  (.A1(v4[26]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M3/c1 ));
 XOR2_X2 \A3/A2/A2/A1/M3/M1/_1_  (.A(v4[26]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M3/s1 ));
 AND2_X1 \A3/A2/A2/A1/M3/M2/_0_  (.A1(\A3/A2/A2/A1/M3/s1 ),
    .A2(\A3/A2/A2/A1/c2 ),
    .ZN(\A3/A2/A2/A1/M3/c2 ));
 XOR2_X2 \A3/A2/A2/A1/M3/M2/_1_  (.A(\A3/A2/A2/A1/M3/s1 ),
    .B(\A3/A2/A2/A1/c2 ),
    .Z(Prod[58]));
 OR2_X1 \A3/A2/A2/A1/M3/_0_  (.A1(\A3/A2/A2/A1/M3/c1 ),
    .A2(\A3/A2/A2/A1/M3/c2 ),
    .ZN(\A3/A2/A2/A1/c3 ));
 AND2_X1 \A3/A2/A2/A1/M4/M1/_0_  (.A1(v4[27]),
    .A2(ground),
    .ZN(\A3/A2/A2/A1/M4/c1 ));
 XOR2_X2 \A3/A2/A2/A1/M4/M1/_1_  (.A(v4[27]),
    .B(ground),
    .Z(\A3/A2/A2/A1/M4/s1 ));
 AND2_X1 \A3/A2/A2/A1/M4/M2/_0_  (.A1(\A3/A2/A2/A1/M4/s1 ),
    .A2(\A3/A2/A2/A1/c3 ),
    .ZN(\A3/A2/A2/A1/M4/c2 ));
 XOR2_X2 \A3/A2/A2/A1/M4/M2/_1_  (.A(\A3/A2/A2/A1/M4/s1 ),
    .B(\A3/A2/A2/A1/c3 ),
    .Z(Prod[59]));
 OR2_X1 \A3/A2/A2/A1/M4/_0_  (.A1(\A3/A2/A2/A1/M4/c1 ),
    .A2(\A3/A2/A2/A1/M4/c2 ),
    .ZN(\A3/A2/A2/c1 ));
 AND2_X1 \A3/A2/A2/A2/M1/M1/_0_  (.A1(v4[28]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M1/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M1/M1/_1_  (.A(v4[28]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M1/s1 ));
 AND2_X1 \A3/A2/A2/A2/M1/M2/_0_  (.A1(\A3/A2/A2/A2/M1/s1 ),
    .A2(\A3/A2/A2/c1 ),
    .ZN(\A3/A2/A2/A2/M1/c2 ));
 XOR2_X2 \A3/A2/A2/A2/M1/M2/_1_  (.A(\A3/A2/A2/A2/M1/s1 ),
    .B(\A3/A2/A2/c1 ),
    .Z(Prod[60]));
 OR2_X1 \A3/A2/A2/A2/M1/_0_  (.A1(\A3/A2/A2/A2/M1/c1 ),
    .A2(\A3/A2/A2/A2/M1/c2 ),
    .ZN(\A3/A2/A2/A2/c1 ));
 AND2_X1 \A3/A2/A2/A2/M2/M1/_0_  (.A1(v4[29]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M2/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M2/M1/_1_  (.A(v4[29]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M2/s1 ));
 AND2_X1 \A3/A2/A2/A2/M2/M2/_0_  (.A1(\A3/A2/A2/A2/M2/s1 ),
    .A2(\A3/A2/A2/A2/c1 ),
    .ZN(\A3/A2/A2/A2/M2/c2 ));
 XOR2_X2 \A3/A2/A2/A2/M2/M2/_1_  (.A(\A3/A2/A2/A2/M2/s1 ),
    .B(\A3/A2/A2/A2/c1 ),
    .Z(Prod[61]));
 OR2_X1 \A3/A2/A2/A2/M2/_0_  (.A1(\A3/A2/A2/A2/M2/c1 ),
    .A2(\A3/A2/A2/A2/M2/c2 ),
    .ZN(\A3/A2/A2/A2/c2 ));
 AND2_X1 \A3/A2/A2/A2/M3/M1/_0_  (.A1(v4[30]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M3/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M3/M1/_1_  (.A(v4[30]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M3/s1 ));
 AND2_X1 \A3/A2/A2/A2/M3/M2/_0_  (.A1(\A3/A2/A2/A2/M3/s1 ),
    .A2(\A3/A2/A2/A2/c2 ),
    .ZN(\A3/A2/A2/A2/M3/c2 ));
 XOR2_X2 \A3/A2/A2/A2/M3/M2/_1_  (.A(\A3/A2/A2/A2/M3/s1 ),
    .B(\A3/A2/A2/A2/c2 ),
    .Z(Prod[62]));
 OR2_X4 \A3/A2/A2/A2/M3/_0_  (.A1(\A3/A2/A2/A2/M3/c1 ),
    .A2(\A3/A2/A2/A2/M3/c2 ),
    .ZN(\A3/A2/A2/A2/c3 ));
 AND2_X1 \A3/A2/A2/A2/M4/M1/_0_  (.A1(v4[31]),
    .A2(ground),
    .ZN(\A3/A2/A2/A2/M4/c1 ));
 XOR2_X2 \A3/A2/A2/A2/M4/M1/_1_  (.A(v4[31]),
    .B(ground),
    .Z(\A3/A2/A2/A2/M4/s1 ));
 AND2_X1 \A3/A2/A2/A2/M4/M2/_0_  (.A1(\A3/A2/A2/A2/M4/s1 ),
    .A2(\A3/A2/A2/A2/c3 ),
    .ZN(\A3/A2/A2/A2/M4/c2 ));
 XOR2_X1 \A3/A2/A2/A2/M4/M2/_1_  (.A(\A3/A2/A2/A2/M4/s1 ),
    .B(\A3/A2/A2/A2/c3 ),
    .Z(Prod[63]));
 OR2_X1 \A3/A2/A2/A2/M4/_0_  (.A1(\A3/A2/A2/A2/M4/c1 ),
    .A2(\A3/A2/A2/A2/M4/c2 ),
    .ZN(overflow));
 AND2_X1 \V1/A1/A1/A1/M1/M1/_0_  (.A1(\V1/v2 [0]),
    .A2(\V1/v3 [0]),
    .ZN(\V1/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M1/M1/_1_  (.A(\V1/v2 [0]),
    .B(\V1/v3 [0]),
    .Z(\V1/A1/A1/A1/M1/s1 ));
 AND2_X1 \V1/A1/A1/A1/M1/M2/_0_  (.A1(\V1/A1/A1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M1/M2/_1_  (.A(\V1/A1/A1/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/s1 [0]));
 OR2_X1 \V1/A1/A1/A1/M1/_0_  (.A1(\V1/A1/A1/A1/M1/c1 ),
    .A2(\V1/A1/A1/A1/M1/c2 ),
    .ZN(\V1/A1/A1/A1/c1 ));
 AND2_X1 \V1/A1/A1/A1/M2/M1/_0_  (.A1(\V1/v2 [1]),
    .A2(\V1/v3 [1]),
    .ZN(\V1/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M2/M1/_1_  (.A(\V1/v2 [1]),
    .B(\V1/v3 [1]),
    .Z(\V1/A1/A1/A1/M2/s1 ));
 AND2_X1 \V1/A1/A1/A1/M2/M2/_0_  (.A1(\V1/A1/A1/A1/M2/s1 ),
    .A2(\V1/A1/A1/A1/c1 ),
    .ZN(\V1/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M2/M2/_1_  (.A(\V1/A1/A1/A1/M2/s1 ),
    .B(\V1/A1/A1/A1/c1 ),
    .Z(\V1/s1 [1]));
 OR2_X1 \V1/A1/A1/A1/M2/_0_  (.A1(\V1/A1/A1/A1/M2/c1 ),
    .A2(\V1/A1/A1/A1/M2/c2 ),
    .ZN(\V1/A1/A1/A1/c2 ));
 AND2_X1 \V1/A1/A1/A1/M3/M1/_0_  (.A1(\V1/v2 [2]),
    .A2(\V1/v3 [2]),
    .ZN(\V1/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M3/M1/_1_  (.A(\V1/v2 [2]),
    .B(\V1/v3 [2]),
    .Z(\V1/A1/A1/A1/M3/s1 ));
 AND2_X1 \V1/A1/A1/A1/M3/M2/_0_  (.A1(\V1/A1/A1/A1/M3/s1 ),
    .A2(\V1/A1/A1/A1/c2 ),
    .ZN(\V1/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M3/M2/_1_  (.A(\V1/A1/A1/A1/M3/s1 ),
    .B(\V1/A1/A1/A1/c2 ),
    .Z(\V1/s1 [2]));
 OR2_X1 \V1/A1/A1/A1/M3/_0_  (.A1(\V1/A1/A1/A1/M3/c1 ),
    .A2(\V1/A1/A1/A1/M3/c2 ),
    .ZN(\V1/A1/A1/A1/c3 ));
 AND2_X1 \V1/A1/A1/A1/M4/M1/_0_  (.A1(\V1/v2 [3]),
    .A2(\V1/v3 [3]),
    .ZN(\V1/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A1/A1/A1/M4/M1/_1_  (.A(\V1/v2 [3]),
    .B(\V1/v3 [3]),
    .Z(\V1/A1/A1/A1/M4/s1 ));
 AND2_X1 \V1/A1/A1/A1/M4/M2/_0_  (.A1(\V1/A1/A1/A1/M4/s1 ),
    .A2(\V1/A1/A1/A1/c3 ),
    .ZN(\V1/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A1/A1/A1/M4/M2/_1_  (.A(\V1/A1/A1/A1/M4/s1 ),
    .B(\V1/A1/A1/A1/c3 ),
    .Z(\V1/s1 [3]));
 OR2_X1 \V1/A1/A1/A1/M4/_0_  (.A1(\V1/A1/A1/A1/M4/c1 ),
    .A2(\V1/A1/A1/A1/M4/c2 ),
    .ZN(\V1/A1/A1/c1 ));
 AND2_X1 \V1/A1/A1/A2/M1/M1/_0_  (.A1(\V1/v2 [4]),
    .A2(\V1/v3 [4]),
    .ZN(\V1/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M1/M1/_1_  (.A(\V1/v2 [4]),
    .B(\V1/v3 [4]),
    .Z(\V1/A1/A1/A2/M1/s1 ));
 AND2_X1 \V1/A1/A1/A2/M1/M2/_0_  (.A1(\V1/A1/A1/A2/M1/s1 ),
    .A2(\V1/A1/A1/c1 ),
    .ZN(\V1/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M1/M2/_1_  (.A(\V1/A1/A1/A2/M1/s1 ),
    .B(\V1/A1/A1/c1 ),
    .Z(\V1/s1 [4]));
 OR2_X1 \V1/A1/A1/A2/M1/_0_  (.A1(\V1/A1/A1/A2/M1/c1 ),
    .A2(\V1/A1/A1/A2/M1/c2 ),
    .ZN(\V1/A1/A1/A2/c1 ));
 AND2_X1 \V1/A1/A1/A2/M2/M1/_0_  (.A1(\V1/v2 [5]),
    .A2(\V1/v3 [5]),
    .ZN(\V1/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M2/M1/_1_  (.A(\V1/v2 [5]),
    .B(\V1/v3 [5]),
    .Z(\V1/A1/A1/A2/M2/s1 ));
 AND2_X1 \V1/A1/A1/A2/M2/M2/_0_  (.A1(\V1/A1/A1/A2/M2/s1 ),
    .A2(\V1/A1/A1/A2/c1 ),
    .ZN(\V1/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M2/M2/_1_  (.A(\V1/A1/A1/A2/M2/s1 ),
    .B(\V1/A1/A1/A2/c1 ),
    .Z(\V1/s1 [5]));
 OR2_X1 \V1/A1/A1/A2/M2/_0_  (.A1(\V1/A1/A1/A2/M2/c1 ),
    .A2(\V1/A1/A1/A2/M2/c2 ),
    .ZN(\V1/A1/A1/A2/c2 ));
 AND2_X1 \V1/A1/A1/A2/M3/M1/_0_  (.A1(\V1/v2 [6]),
    .A2(\V1/v3 [6]),
    .ZN(\V1/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M3/M1/_1_  (.A(\V1/v2 [6]),
    .B(\V1/v3 [6]),
    .Z(\V1/A1/A1/A2/M3/s1 ));
 AND2_X1 \V1/A1/A1/A2/M3/M2/_0_  (.A1(\V1/A1/A1/A2/M3/s1 ),
    .A2(\V1/A1/A1/A2/c2 ),
    .ZN(\V1/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M3/M2/_1_  (.A(\V1/A1/A1/A2/M3/s1 ),
    .B(\V1/A1/A1/A2/c2 ),
    .Z(\V1/s1 [6]));
 OR2_X1 \V1/A1/A1/A2/M3/_0_  (.A1(\V1/A1/A1/A2/M3/c1 ),
    .A2(\V1/A1/A1/A2/M3/c2 ),
    .ZN(\V1/A1/A1/A2/c3 ));
 AND2_X1 \V1/A1/A1/A2/M4/M1/_0_  (.A1(\V1/v2 [7]),
    .A2(\V1/v3 [7]),
    .ZN(\V1/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A1/A1/A2/M4/M1/_1_  (.A(\V1/v2 [7]),
    .B(\V1/v3 [7]),
    .Z(\V1/A1/A1/A2/M4/s1 ));
 AND2_X1 \V1/A1/A1/A2/M4/M2/_0_  (.A1(\V1/A1/A1/A2/M4/s1 ),
    .A2(\V1/A1/A1/A2/c3 ),
    .ZN(\V1/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A1/A1/A2/M4/M2/_1_  (.A(\V1/A1/A1/A2/M4/s1 ),
    .B(\V1/A1/A1/A2/c3 ),
    .Z(\V1/s1 [7]));
 OR2_X1 \V1/A1/A1/A2/M4/_0_  (.A1(\V1/A1/A1/A2/M4/c1 ),
    .A2(\V1/A1/A1/A2/M4/c2 ),
    .ZN(\V1/A1/c1 ));
 AND2_X1 \V1/A1/A2/A1/M1/M1/_0_  (.A1(\V1/v2 [8]),
    .A2(\V1/v3 [8]),
    .ZN(\V1/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M1/M1/_1_  (.A(\V1/v2 [8]),
    .B(\V1/v3 [8]),
    .Z(\V1/A1/A2/A1/M1/s1 ));
 AND2_X1 \V1/A1/A2/A1/M1/M2/_0_  (.A1(\V1/A1/A2/A1/M1/s1 ),
    .A2(\V1/A1/c1 ),
    .ZN(\V1/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M1/M2/_1_  (.A(\V1/A1/A2/A1/M1/s1 ),
    .B(\V1/A1/c1 ),
    .Z(\V1/s1 [8]));
 OR2_X1 \V1/A1/A2/A1/M1/_0_  (.A1(\V1/A1/A2/A1/M1/c1 ),
    .A2(\V1/A1/A2/A1/M1/c2 ),
    .ZN(\V1/A1/A2/A1/c1 ));
 AND2_X1 \V1/A1/A2/A1/M2/M1/_0_  (.A1(\V1/v2 [9]),
    .A2(\V1/v3 [9]),
    .ZN(\V1/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M2/M1/_1_  (.A(\V1/v2 [9]),
    .B(\V1/v3 [9]),
    .Z(\V1/A1/A2/A1/M2/s1 ));
 AND2_X1 \V1/A1/A2/A1/M2/M2/_0_  (.A1(\V1/A1/A2/A1/M2/s1 ),
    .A2(\V1/A1/A2/A1/c1 ),
    .ZN(\V1/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M2/M2/_1_  (.A(\V1/A1/A2/A1/M2/s1 ),
    .B(\V1/A1/A2/A1/c1 ),
    .Z(\V1/s1 [9]));
 OR2_X1 \V1/A1/A2/A1/M2/_0_  (.A1(\V1/A1/A2/A1/M2/c1 ),
    .A2(\V1/A1/A2/A1/M2/c2 ),
    .ZN(\V1/A1/A2/A1/c2 ));
 AND2_X1 \V1/A1/A2/A1/M3/M1/_0_  (.A1(\V1/v2 [10]),
    .A2(\V1/v3 [10]),
    .ZN(\V1/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M3/M1/_1_  (.A(\V1/v2 [10]),
    .B(\V1/v3 [10]),
    .Z(\V1/A1/A2/A1/M3/s1 ));
 AND2_X1 \V1/A1/A2/A1/M3/M2/_0_  (.A1(\V1/A1/A2/A1/M3/s1 ),
    .A2(\V1/A1/A2/A1/c2 ),
    .ZN(\V1/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M3/M2/_1_  (.A(\V1/A1/A2/A1/M3/s1 ),
    .B(\V1/A1/A2/A1/c2 ),
    .Z(\V1/s1 [10]));
 OR2_X1 \V1/A1/A2/A1/M3/_0_  (.A1(\V1/A1/A2/A1/M3/c1 ),
    .A2(\V1/A1/A2/A1/M3/c2 ),
    .ZN(\V1/A1/A2/A1/c3 ));
 AND2_X1 \V1/A1/A2/A1/M4/M1/_0_  (.A1(\V1/v2 [11]),
    .A2(\V1/v3 [11]),
    .ZN(\V1/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A1/A2/A1/M4/M1/_1_  (.A(\V1/v2 [11]),
    .B(\V1/v3 [11]),
    .Z(\V1/A1/A2/A1/M4/s1 ));
 AND2_X1 \V1/A1/A2/A1/M4/M2/_0_  (.A1(\V1/A1/A2/A1/M4/s1 ),
    .A2(\V1/A1/A2/A1/c3 ),
    .ZN(\V1/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A1/A2/A1/M4/M2/_1_  (.A(\V1/A1/A2/A1/M4/s1 ),
    .B(\V1/A1/A2/A1/c3 ),
    .Z(\V1/s1 [11]));
 OR2_X1 \V1/A1/A2/A1/M4/_0_  (.A1(\V1/A1/A2/A1/M4/c1 ),
    .A2(\V1/A1/A2/A1/M4/c2 ),
    .ZN(\V1/A1/A2/c1 ));
 AND2_X1 \V1/A1/A2/A2/M1/M1/_0_  (.A1(\V1/v2 [12]),
    .A2(\V1/v3 [12]),
    .ZN(\V1/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M1/M1/_1_  (.A(\V1/v2 [12]),
    .B(\V1/v3 [12]),
    .Z(\V1/A1/A2/A2/M1/s1 ));
 AND2_X1 \V1/A1/A2/A2/M1/M2/_0_  (.A1(\V1/A1/A2/A2/M1/s1 ),
    .A2(\V1/A1/A2/c1 ),
    .ZN(\V1/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M1/M2/_1_  (.A(\V1/A1/A2/A2/M1/s1 ),
    .B(\V1/A1/A2/c1 ),
    .Z(\V1/s1 [12]));
 OR2_X1 \V1/A1/A2/A2/M1/_0_  (.A1(\V1/A1/A2/A2/M1/c1 ),
    .A2(\V1/A1/A2/A2/M1/c2 ),
    .ZN(\V1/A1/A2/A2/c1 ));
 AND2_X1 \V1/A1/A2/A2/M2/M1/_0_  (.A1(\V1/v2 [13]),
    .A2(\V1/v3 [13]),
    .ZN(\V1/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M2/M1/_1_  (.A(\V1/v2 [13]),
    .B(\V1/v3 [13]),
    .Z(\V1/A1/A2/A2/M2/s1 ));
 AND2_X1 \V1/A1/A2/A2/M2/M2/_0_  (.A1(\V1/A1/A2/A2/M2/s1 ),
    .A2(\V1/A1/A2/A2/c1 ),
    .ZN(\V1/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M2/M2/_1_  (.A(\V1/A1/A2/A2/M2/s1 ),
    .B(\V1/A1/A2/A2/c1 ),
    .Z(\V1/s1 [13]));
 OR2_X1 \V1/A1/A2/A2/M2/_0_  (.A1(\V1/A1/A2/A2/M2/c1 ),
    .A2(\V1/A1/A2/A2/M2/c2 ),
    .ZN(\V1/A1/A2/A2/c2 ));
 AND2_X1 \V1/A1/A2/A2/M3/M1/_0_  (.A1(\V1/v2 [14]),
    .A2(\V1/v3 [14]),
    .ZN(\V1/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M3/M1/_1_  (.A(\V1/v2 [14]),
    .B(\V1/v3 [14]),
    .Z(\V1/A1/A2/A2/M3/s1 ));
 AND2_X1 \V1/A1/A2/A2/M3/M2/_0_  (.A1(\V1/A1/A2/A2/M3/s1 ),
    .A2(\V1/A1/A2/A2/c2 ),
    .ZN(\V1/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M3/M2/_1_  (.A(\V1/A1/A2/A2/M3/s1 ),
    .B(\V1/A1/A2/A2/c2 ),
    .Z(\V1/s1 [14]));
 OR2_X1 \V1/A1/A2/A2/M3/_0_  (.A1(\V1/A1/A2/A2/M3/c1 ),
    .A2(\V1/A1/A2/A2/M3/c2 ),
    .ZN(\V1/A1/A2/A2/c3 ));
 AND2_X1 \V1/A1/A2/A2/M4/M1/_0_  (.A1(\V1/v2 [15]),
    .A2(\V1/v3 [15]),
    .ZN(\V1/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A1/A2/A2/M4/M1/_1_  (.A(\V1/v2 [15]),
    .B(\V1/v3 [15]),
    .Z(\V1/A1/A2/A2/M4/s1 ));
 AND2_X1 \V1/A1/A2/A2/M4/M2/_0_  (.A1(\V1/A1/A2/A2/M4/s1 ),
    .A2(\V1/A1/A2/A2/c3 ),
    .ZN(\V1/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A1/A2/A2/M4/M2/_1_  (.A(\V1/A1/A2/A2/M4/s1 ),
    .B(\V1/A1/A2/A2/c3 ),
    .Z(\V1/s1 [15]));
 OR2_X1 \V1/A1/A2/A2/M4/_0_  (.A1(\V1/A1/A2/A2/M4/c1 ),
    .A2(\V1/A1/A2/A2/M4/c2 ),
    .ZN(\V1/c1 ));
 AND2_X1 \V1/A2/A1/A1/M1/M1/_0_  (.A1(\V1/s1 [0]),
    .A2(\V1/v1 [8]),
    .ZN(\V1/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M1/M1/_1_  (.A(\V1/s1 [0]),
    .B(\V1/v1 [8]),
    .Z(\V1/A2/A1/A1/M1/s1 ));
 AND2_X1 \V1/A2/A1/A1/M1/M2/_0_  (.A1(\V1/A2/A1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M1/M2/_1_  (.A(\V1/A2/A1/A1/M1/s1 ),
    .B(net4),
    .Z(v1[8]));
 OR2_X1 \V1/A2/A1/A1/M1/_0_  (.A1(\V1/A2/A1/A1/M1/c1 ),
    .A2(\V1/A2/A1/A1/M1/c2 ),
    .ZN(\V1/A2/A1/A1/c1 ));
 AND2_X1 \V1/A2/A1/A1/M2/M1/_0_  (.A1(\V1/s1 [1]),
    .A2(\V1/v1 [9]),
    .ZN(\V1/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M2/M1/_1_  (.A(\V1/s1 [1]),
    .B(\V1/v1 [9]),
    .Z(\V1/A2/A1/A1/M2/s1 ));
 AND2_X1 \V1/A2/A1/A1/M2/M2/_0_  (.A1(\V1/A2/A1/A1/M2/s1 ),
    .A2(\V1/A2/A1/A1/c1 ),
    .ZN(\V1/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M2/M2/_1_  (.A(\V1/A2/A1/A1/M2/s1 ),
    .B(\V1/A2/A1/A1/c1 ),
    .Z(v1[9]));
 OR2_X1 \V1/A2/A1/A1/M2/_0_  (.A1(\V1/A2/A1/A1/M2/c1 ),
    .A2(\V1/A2/A1/A1/M2/c2 ),
    .ZN(\V1/A2/A1/A1/c2 ));
 AND2_X1 \V1/A2/A1/A1/M3/M1/_0_  (.A1(\V1/s1 [2]),
    .A2(\V1/v1 [10]),
    .ZN(\V1/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M3/M1/_1_  (.A(\V1/s1 [2]),
    .B(\V1/v1 [10]),
    .Z(\V1/A2/A1/A1/M3/s1 ));
 AND2_X1 \V1/A2/A1/A1/M3/M2/_0_  (.A1(\V1/A2/A1/A1/M3/s1 ),
    .A2(\V1/A2/A1/A1/c2 ),
    .ZN(\V1/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M3/M2/_1_  (.A(\V1/A2/A1/A1/M3/s1 ),
    .B(\V1/A2/A1/A1/c2 ),
    .Z(v1[10]));
 OR2_X1 \V1/A2/A1/A1/M3/_0_  (.A1(\V1/A2/A1/A1/M3/c1 ),
    .A2(\V1/A2/A1/A1/M3/c2 ),
    .ZN(\V1/A2/A1/A1/c3 ));
 AND2_X1 \V1/A2/A1/A1/M4/M1/_0_  (.A1(\V1/s1 [3]),
    .A2(\V1/v1 [11]),
    .ZN(\V1/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A2/A1/A1/M4/M1/_1_  (.A(\V1/s1 [3]),
    .B(\V1/v1 [11]),
    .Z(\V1/A2/A1/A1/M4/s1 ));
 AND2_X1 \V1/A2/A1/A1/M4/M2/_0_  (.A1(\V1/A2/A1/A1/M4/s1 ),
    .A2(\V1/A2/A1/A1/c3 ),
    .ZN(\V1/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A2/A1/A1/M4/M2/_1_  (.A(\V1/A2/A1/A1/M4/s1 ),
    .B(\V1/A2/A1/A1/c3 ),
    .Z(v1[11]));
 OR2_X1 \V1/A2/A1/A1/M4/_0_  (.A1(\V1/A2/A1/A1/M4/c1 ),
    .A2(\V1/A2/A1/A1/M4/c2 ),
    .ZN(\V1/A2/A1/c1 ));
 AND2_X1 \V1/A2/A1/A2/M1/M1/_0_  (.A1(\V1/s1 [4]),
    .A2(\V1/v1 [12]),
    .ZN(\V1/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M1/M1/_1_  (.A(\V1/s1 [4]),
    .B(\V1/v1 [12]),
    .Z(\V1/A2/A1/A2/M1/s1 ));
 AND2_X1 \V1/A2/A1/A2/M1/M2/_0_  (.A1(\V1/A2/A1/A2/M1/s1 ),
    .A2(\V1/A2/A1/c1 ),
    .ZN(\V1/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M1/M2/_1_  (.A(\V1/A2/A1/A2/M1/s1 ),
    .B(\V1/A2/A1/c1 ),
    .Z(v1[12]));
 OR2_X1 \V1/A2/A1/A2/M1/_0_  (.A1(\V1/A2/A1/A2/M1/c1 ),
    .A2(\V1/A2/A1/A2/M1/c2 ),
    .ZN(\V1/A2/A1/A2/c1 ));
 AND2_X1 \V1/A2/A1/A2/M2/M1/_0_  (.A1(\V1/s1 [5]),
    .A2(\V1/v1 [13]),
    .ZN(\V1/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M2/M1/_1_  (.A(\V1/s1 [5]),
    .B(\V1/v1 [13]),
    .Z(\V1/A2/A1/A2/M2/s1 ));
 AND2_X1 \V1/A2/A1/A2/M2/M2/_0_  (.A1(\V1/A2/A1/A2/M2/s1 ),
    .A2(\V1/A2/A1/A2/c1 ),
    .ZN(\V1/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M2/M2/_1_  (.A(\V1/A2/A1/A2/M2/s1 ),
    .B(\V1/A2/A1/A2/c1 ),
    .Z(v1[13]));
 OR2_X2 \V1/A2/A1/A2/M2/_0_  (.A1(\V1/A2/A1/A2/M2/c1 ),
    .A2(\V1/A2/A1/A2/M2/c2 ),
    .ZN(\V1/A2/A1/A2/c2 ));
 AND2_X1 \V1/A2/A1/A2/M3/M1/_0_  (.A1(\V1/s1 [6]),
    .A2(\V1/v1 [14]),
    .ZN(\V1/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M3/M1/_1_  (.A(\V1/s1 [6]),
    .B(\V1/v1 [14]),
    .Z(\V1/A2/A1/A2/M3/s1 ));
 AND2_X1 \V1/A2/A1/A2/M3/M2/_0_  (.A1(\V1/A2/A1/A2/M3/s1 ),
    .A2(\V1/A2/A1/A2/c2 ),
    .ZN(\V1/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M3/M2/_1_  (.A(\V1/A2/A1/A2/M3/s1 ),
    .B(\V1/A2/A1/A2/c2 ),
    .Z(v1[14]));
 OR2_X1 \V1/A2/A1/A2/M3/_0_  (.A1(\V1/A2/A1/A2/M3/c1 ),
    .A2(\V1/A2/A1/A2/M3/c2 ),
    .ZN(\V1/A2/A1/A2/c3 ));
 AND2_X1 \V1/A2/A1/A2/M4/M1/_0_  (.A1(\V1/s1 [7]),
    .A2(\V1/v1 [15]),
    .ZN(\V1/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A2/A1/A2/M4/M1/_1_  (.A(\V1/s1 [7]),
    .B(\V1/v1 [15]),
    .Z(\V1/A2/A1/A2/M4/s1 ));
 AND2_X1 \V1/A2/A1/A2/M4/M2/_0_  (.A1(\V1/A2/A1/A2/M4/s1 ),
    .A2(\V1/A2/A1/A2/c3 ),
    .ZN(\V1/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A2/A1/A2/M4/M2/_1_  (.A(\V1/A2/A1/A2/M4/s1 ),
    .B(\V1/A2/A1/A2/c3 ),
    .Z(v1[15]));
 OR2_X1 \V1/A2/A1/A2/M4/_0_  (.A1(\V1/A2/A1/A2/M4/c1 ),
    .A2(\V1/A2/A1/A2/M4/c2 ),
    .ZN(\V1/A2/c1 ));
 AND2_X1 \V1/A2/A2/A1/M1/M1/_0_  (.A1(\V1/s1 [8]),
    .A2(net3),
    .ZN(\V1/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M1/M1/_1_  (.A(\V1/s1 [8]),
    .B(net3),
    .Z(\V1/A2/A2/A1/M1/s1 ));
 AND2_X1 \V1/A2/A2/A1/M1/M2/_0_  (.A1(\V1/A2/A2/A1/M1/s1 ),
    .A2(\V1/A2/c1 ),
    .ZN(\V1/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M1/M2/_1_  (.A(\V1/A2/A2/A1/M1/s1 ),
    .B(\V1/A2/c1 ),
    .Z(\V1/s2 [8]));
 OR2_X1 \V1/A2/A2/A1/M1/_0_  (.A1(\V1/A2/A2/A1/M1/c1 ),
    .A2(\V1/A2/A2/A1/M1/c2 ),
    .ZN(\V1/A2/A2/A1/c1 ));
 AND2_X1 \V1/A2/A2/A1/M2/M1/_0_  (.A1(\V1/s1 [9]),
    .A2(net3),
    .ZN(\V1/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M2/M1/_1_  (.A(\V1/s1 [9]),
    .B(net3),
    .Z(\V1/A2/A2/A1/M2/s1 ));
 AND2_X1 \V1/A2/A2/A1/M2/M2/_0_  (.A1(\V1/A2/A2/A1/M2/s1 ),
    .A2(\V1/A2/A2/A1/c1 ),
    .ZN(\V1/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M2/M2/_1_  (.A(\V1/A2/A2/A1/M2/s1 ),
    .B(\V1/A2/A2/A1/c1 ),
    .Z(\V1/s2 [9]));
 OR2_X1 \V1/A2/A2/A1/M2/_0_  (.A1(\V1/A2/A2/A1/M2/c1 ),
    .A2(\V1/A2/A2/A1/M2/c2 ),
    .ZN(\V1/A2/A2/A1/c2 ));
 AND2_X1 \V1/A2/A2/A1/M3/M1/_0_  (.A1(\V1/s1 [10]),
    .A2(net3),
    .ZN(\V1/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M3/M1/_1_  (.A(\V1/s1 [10]),
    .B(net3),
    .Z(\V1/A2/A2/A1/M3/s1 ));
 AND2_X1 \V1/A2/A2/A1/M3/M2/_0_  (.A1(\V1/A2/A2/A1/M3/s1 ),
    .A2(\V1/A2/A2/A1/c2 ),
    .ZN(\V1/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M3/M2/_1_  (.A(\V1/A2/A2/A1/M3/s1 ),
    .B(\V1/A2/A2/A1/c2 ),
    .Z(\V1/s2 [10]));
 OR2_X1 \V1/A2/A2/A1/M3/_0_  (.A1(\V1/A2/A2/A1/M3/c1 ),
    .A2(\V1/A2/A2/A1/M3/c2 ),
    .ZN(\V1/A2/A2/A1/c3 ));
 AND2_X1 \V1/A2/A2/A1/M4/M1/_0_  (.A1(\V1/s1 [11]),
    .A2(net3),
    .ZN(\V1/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A2/A2/A1/M4/M1/_1_  (.A(\V1/s1 [11]),
    .B(net3),
    .Z(\V1/A2/A2/A1/M4/s1 ));
 AND2_X1 \V1/A2/A2/A1/M4/M2/_0_  (.A1(\V1/A2/A2/A1/M4/s1 ),
    .A2(\V1/A2/A2/A1/c3 ),
    .ZN(\V1/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A2/A2/A1/M4/M2/_1_  (.A(\V1/A2/A2/A1/M4/s1 ),
    .B(\V1/A2/A2/A1/c3 ),
    .Z(\V1/s2 [11]));
 OR2_X1 \V1/A2/A2/A1/M4/_0_  (.A1(\V1/A2/A2/A1/M4/c1 ),
    .A2(\V1/A2/A2/A1/M4/c2 ),
    .ZN(\V1/A2/A2/c1 ));
 AND2_X1 \V1/A2/A2/A2/M1/M1/_0_  (.A1(\V1/s1 [12]),
    .A2(net3),
    .ZN(\V1/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M1/M1/_1_  (.A(\V1/s1 [12]),
    .B(net3),
    .Z(\V1/A2/A2/A2/M1/s1 ));
 AND2_X1 \V1/A2/A2/A2/M1/M2/_0_  (.A1(\V1/A2/A2/A2/M1/s1 ),
    .A2(\V1/A2/A2/c1 ),
    .ZN(\V1/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M1/M2/_1_  (.A(\V1/A2/A2/A2/M1/s1 ),
    .B(\V1/A2/A2/c1 ),
    .Z(\V1/s2 [12]));
 OR2_X1 \V1/A2/A2/A2/M1/_0_  (.A1(\V1/A2/A2/A2/M1/c1 ),
    .A2(\V1/A2/A2/A2/M1/c2 ),
    .ZN(\V1/A2/A2/A2/c1 ));
 AND2_X1 \V1/A2/A2/A2/M2/M1/_0_  (.A1(\V1/s1 [13]),
    .A2(net3),
    .ZN(\V1/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M2/M1/_1_  (.A(\V1/s1 [13]),
    .B(net3),
    .Z(\V1/A2/A2/A2/M2/s1 ));
 AND2_X1 \V1/A2/A2/A2/M2/M2/_0_  (.A1(\V1/A2/A2/A2/M2/s1 ),
    .A2(\V1/A2/A2/A2/c1 ),
    .ZN(\V1/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M2/M2/_1_  (.A(\V1/A2/A2/A2/M2/s1 ),
    .B(\V1/A2/A2/A2/c1 ),
    .Z(\V1/s2 [13]));
 OR2_X1 \V1/A2/A2/A2/M2/_0_  (.A1(\V1/A2/A2/A2/M2/c1 ),
    .A2(\V1/A2/A2/A2/M2/c2 ),
    .ZN(\V1/A2/A2/A2/c2 ));
 AND2_X1 \V1/A2/A2/A2/M3/M1/_0_  (.A1(\V1/s1 [14]),
    .A2(net3),
    .ZN(\V1/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M3/M1/_1_  (.A(\V1/s1 [14]),
    .B(net3),
    .Z(\V1/A2/A2/A2/M3/s1 ));
 AND2_X1 \V1/A2/A2/A2/M3/M2/_0_  (.A1(\V1/A2/A2/A2/M3/s1 ),
    .A2(\V1/A2/A2/A2/c2 ),
    .ZN(\V1/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M3/M2/_1_  (.A(\V1/A2/A2/A2/M3/s1 ),
    .B(\V1/A2/A2/A2/c2 ),
    .Z(\V1/s2 [14]));
 OR2_X1 \V1/A2/A2/A2/M3/_0_  (.A1(\V1/A2/A2/A2/M3/c1 ),
    .A2(\V1/A2/A2/A2/M3/c2 ),
    .ZN(\V1/A2/A2/A2/c3 ));
 AND2_X1 \V1/A2/A2/A2/M4/M1/_0_  (.A1(\V1/s1 [15]),
    .A2(net3),
    .ZN(\V1/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A2/A2/A2/M4/M1/_1_  (.A(\V1/s1 [15]),
    .B(net3),
    .Z(\V1/A2/A2/A2/M4/s1 ));
 AND2_X1 \V1/A2/A2/A2/M4/M2/_0_  (.A1(\V1/A2/A2/A2/M4/s1 ),
    .A2(\V1/A2/A2/A2/c3 ),
    .ZN(\V1/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A2/A2/A2/M4/M2/_1_  (.A(\V1/A2/A2/A2/M4/s1 ),
    .B(\V1/A2/A2/A2/c3 ),
    .Z(\V1/s2 [15]));
 OR2_X1 \V1/A2/A2/A2/M4/_0_  (.A1(\V1/A2/A2/A2/M4/c1 ),
    .A2(\V1/A2/A2/A2/M4/c2 ),
    .ZN(\V1/c2 ));
 AND2_X1 \V1/A3/A1/A1/M1/M1/_0_  (.A1(\V1/v4 [0]),
    .A2(\V1/s2 [8]),
    .ZN(\V1/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M1/M1/_1_  (.A(\V1/v4 [0]),
    .B(\V1/s2 [8]),
    .Z(\V1/A3/A1/A1/M1/s1 ));
 AND2_X1 \V1/A3/A1/A1/M1/M2/_0_  (.A1(\V1/A3/A1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M1/M2/_1_  (.A(\V1/A3/A1/A1/M1/s1 ),
    .B(net3),
    .Z(v1[16]));
 OR2_X1 \V1/A3/A1/A1/M1/_0_  (.A1(\V1/A3/A1/A1/M1/c1 ),
    .A2(\V1/A3/A1/A1/M1/c2 ),
    .ZN(\V1/A3/A1/A1/c1 ));
 AND2_X1 \V1/A3/A1/A1/M2/M1/_0_  (.A1(\V1/v4 [1]),
    .A2(\V1/s2 [9]),
    .ZN(\V1/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M2/M1/_1_  (.A(\V1/v4 [1]),
    .B(\V1/s2 [9]),
    .Z(\V1/A3/A1/A1/M2/s1 ));
 AND2_X1 \V1/A3/A1/A1/M2/M2/_0_  (.A1(\V1/A3/A1/A1/M2/s1 ),
    .A2(\V1/A3/A1/A1/c1 ),
    .ZN(\V1/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M2/M2/_1_  (.A(\V1/A3/A1/A1/M2/s1 ),
    .B(\V1/A3/A1/A1/c1 ),
    .Z(v1[17]));
 OR2_X1 \V1/A3/A1/A1/M2/_0_  (.A1(\V1/A3/A1/A1/M2/c1 ),
    .A2(\V1/A3/A1/A1/M2/c2 ),
    .ZN(\V1/A3/A1/A1/c2 ));
 AND2_X1 \V1/A3/A1/A1/M3/M1/_0_  (.A1(\V1/v4 [2]),
    .A2(\V1/s2 [10]),
    .ZN(\V1/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M3/M1/_1_  (.A(\V1/v4 [2]),
    .B(\V1/s2 [10]),
    .Z(\V1/A3/A1/A1/M3/s1 ));
 AND2_X1 \V1/A3/A1/A1/M3/M2/_0_  (.A1(\V1/A3/A1/A1/M3/s1 ),
    .A2(\V1/A3/A1/A1/c2 ),
    .ZN(\V1/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M3/M2/_1_  (.A(\V1/A3/A1/A1/M3/s1 ),
    .B(\V1/A3/A1/A1/c2 ),
    .Z(v1[18]));
 OR2_X1 \V1/A3/A1/A1/M3/_0_  (.A1(\V1/A3/A1/A1/M3/c1 ),
    .A2(\V1/A3/A1/A1/M3/c2 ),
    .ZN(\V1/A3/A1/A1/c3 ));
 AND2_X1 \V1/A3/A1/A1/M4/M1/_0_  (.A1(\V1/v4 [3]),
    .A2(\V1/s2 [11]),
    .ZN(\V1/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V1/A3/A1/A1/M4/M1/_1_  (.A(\V1/v4 [3]),
    .B(\V1/s2 [11]),
    .Z(\V1/A3/A1/A1/M4/s1 ));
 AND2_X1 \V1/A3/A1/A1/M4/M2/_0_  (.A1(\V1/A3/A1/A1/M4/s1 ),
    .A2(\V1/A3/A1/A1/c3 ),
    .ZN(\V1/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V1/A3/A1/A1/M4/M2/_1_  (.A(\V1/A3/A1/A1/M4/s1 ),
    .B(\V1/A3/A1/A1/c3 ),
    .Z(v1[19]));
 OR2_X1 \V1/A3/A1/A1/M4/_0_  (.A1(\V1/A3/A1/A1/M4/c1 ),
    .A2(\V1/A3/A1/A1/M4/c2 ),
    .ZN(\V1/A3/A1/c1 ));
 AND2_X1 \V1/A3/A1/A2/M1/M1/_0_  (.A1(\V1/v4 [4]),
    .A2(\V1/s2 [12]),
    .ZN(\V1/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M1/M1/_1_  (.A(\V1/v4 [4]),
    .B(\V1/s2 [12]),
    .Z(\V1/A3/A1/A2/M1/s1 ));
 AND2_X1 \V1/A3/A1/A2/M1/M2/_0_  (.A1(\V1/A3/A1/A2/M1/s1 ),
    .A2(\V1/A3/A1/c1 ),
    .ZN(\V1/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M1/M2/_1_  (.A(\V1/A3/A1/A2/M1/s1 ),
    .B(\V1/A3/A1/c1 ),
    .Z(v1[20]));
 OR2_X1 \V1/A3/A1/A2/M1/_0_  (.A1(\V1/A3/A1/A2/M1/c1 ),
    .A2(\V1/A3/A1/A2/M1/c2 ),
    .ZN(\V1/A3/A1/A2/c1 ));
 AND2_X1 \V1/A3/A1/A2/M2/M1/_0_  (.A1(\V1/v4 [5]),
    .A2(\V1/s2 [13]),
    .ZN(\V1/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M2/M1/_1_  (.A(\V1/v4 [5]),
    .B(\V1/s2 [13]),
    .Z(\V1/A3/A1/A2/M2/s1 ));
 AND2_X1 \V1/A3/A1/A2/M2/M2/_0_  (.A1(\V1/A3/A1/A2/M2/s1 ),
    .A2(\V1/A3/A1/A2/c1 ),
    .ZN(\V1/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M2/M2/_1_  (.A(\V1/A3/A1/A2/M2/s1 ),
    .B(\V1/A3/A1/A2/c1 ),
    .Z(v1[21]));
 OR2_X1 \V1/A3/A1/A2/M2/_0_  (.A1(\V1/A3/A1/A2/M2/c1 ),
    .A2(\V1/A3/A1/A2/M2/c2 ),
    .ZN(\V1/A3/A1/A2/c2 ));
 AND2_X1 \V1/A3/A1/A2/M3/M1/_0_  (.A1(\V1/v4 [6]),
    .A2(\V1/s2 [14]),
    .ZN(\V1/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M3/M1/_1_  (.A(\V1/v4 [6]),
    .B(\V1/s2 [14]),
    .Z(\V1/A3/A1/A2/M3/s1 ));
 AND2_X1 \V1/A3/A1/A2/M3/M2/_0_  (.A1(\V1/A3/A1/A2/M3/s1 ),
    .A2(\V1/A3/A1/A2/c2 ),
    .ZN(\V1/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M3/M2/_1_  (.A(\V1/A3/A1/A2/M3/s1 ),
    .B(\V1/A3/A1/A2/c2 ),
    .Z(v1[22]));
 OR2_X1 \V1/A3/A1/A2/M3/_0_  (.A1(\V1/A3/A1/A2/M3/c1 ),
    .A2(\V1/A3/A1/A2/M3/c2 ),
    .ZN(\V1/A3/A1/A2/c3 ));
 AND2_X1 \V1/A3/A1/A2/M4/M1/_0_  (.A1(\V1/v4 [7]),
    .A2(\V1/s2 [15]),
    .ZN(\V1/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V1/A3/A1/A2/M4/M1/_1_  (.A(\V1/v4 [7]),
    .B(\V1/s2 [15]),
    .Z(\V1/A3/A1/A2/M4/s1 ));
 AND2_X1 \V1/A3/A1/A2/M4/M2/_0_  (.A1(\V1/A3/A1/A2/M4/s1 ),
    .A2(\V1/A3/A1/A2/c3 ),
    .ZN(\V1/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V1/A3/A1/A2/M4/M2/_1_  (.A(\V1/A3/A1/A2/M4/s1 ),
    .B(\V1/A3/A1/A2/c3 ),
    .Z(v1[23]));
 OR2_X2 \V1/A3/A1/A2/M4/_0_  (.A1(\V1/A3/A1/A2/M4/c1 ),
    .A2(\V1/A3/A1/A2/M4/c2 ),
    .ZN(\V1/A3/c1 ));
 AND2_X1 \V1/A3/A2/A1/M1/M1/_0_  (.A1(\V1/v4 [8]),
    .A2(\V1/c3 ),
    .ZN(\V1/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M1/M1/_1_  (.A(\V1/v4 [8]),
    .B(\V1/c3 ),
    .Z(\V1/A3/A2/A1/M1/s1 ));
 AND2_X1 \V1/A3/A2/A1/M1/M2/_0_  (.A1(\V1/A3/A2/A1/M1/s1 ),
    .A2(\V1/A3/c1 ),
    .ZN(\V1/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M1/M2/_1_  (.A(\V1/A3/A2/A1/M1/s1 ),
    .B(\V1/A3/c1 ),
    .Z(v1[24]));
 OR2_X1 \V1/A3/A2/A1/M1/_0_  (.A1(\V1/A3/A2/A1/M1/c1 ),
    .A2(\V1/A3/A2/A1/M1/c2 ),
    .ZN(\V1/A3/A2/A1/c1 ));
 AND2_X1 \V1/A3/A2/A1/M2/M1/_0_  (.A1(\V1/v4 [9]),
    .A2(net6),
    .ZN(\V1/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M2/M1/_1_  (.A(\V1/v4 [9]),
    .B(net6),
    .Z(\V1/A3/A2/A1/M2/s1 ));
 AND2_X1 \V1/A3/A2/A1/M2/M2/_0_  (.A1(\V1/A3/A2/A1/M2/s1 ),
    .A2(\V1/A3/A2/A1/c1 ),
    .ZN(\V1/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M2/M2/_1_  (.A(\V1/A3/A2/A1/M2/s1 ),
    .B(\V1/A3/A2/A1/c1 ),
    .Z(v1[25]));
 OR2_X1 \V1/A3/A2/A1/M2/_0_  (.A1(\V1/A3/A2/A1/M2/c1 ),
    .A2(\V1/A3/A2/A1/M2/c2 ),
    .ZN(\V1/A3/A2/A1/c2 ));
 AND2_X1 \V1/A3/A2/A1/M3/M1/_0_  (.A1(\V1/v4 [10]),
    .A2(net6),
    .ZN(\V1/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M3/M1/_1_  (.A(\V1/v4 [10]),
    .B(net6),
    .Z(\V1/A3/A2/A1/M3/s1 ));
 AND2_X1 \V1/A3/A2/A1/M3/M2/_0_  (.A1(\V1/A3/A2/A1/M3/s1 ),
    .A2(\V1/A3/A2/A1/c2 ),
    .ZN(\V1/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M3/M2/_1_  (.A(\V1/A3/A2/A1/M3/s1 ),
    .B(\V1/A3/A2/A1/c2 ),
    .Z(v1[26]));
 OR2_X1 \V1/A3/A2/A1/M3/_0_  (.A1(\V1/A3/A2/A1/M3/c1 ),
    .A2(\V1/A3/A2/A1/M3/c2 ),
    .ZN(\V1/A3/A2/A1/c3 ));
 AND2_X1 \V1/A3/A2/A1/M4/M1/_0_  (.A1(\V1/v4 [11]),
    .A2(net6),
    .ZN(\V1/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V1/A3/A2/A1/M4/M1/_1_  (.A(\V1/v4 [11]),
    .B(net6),
    .Z(\V1/A3/A2/A1/M4/s1 ));
 AND2_X1 \V1/A3/A2/A1/M4/M2/_0_  (.A1(\V1/A3/A2/A1/M4/s1 ),
    .A2(\V1/A3/A2/A1/c3 ),
    .ZN(\V1/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V1/A3/A2/A1/M4/M2/_1_  (.A(\V1/A3/A2/A1/M4/s1 ),
    .B(\V1/A3/A2/A1/c3 ),
    .Z(v1[27]));
 OR2_X1 \V1/A3/A2/A1/M4/_0_  (.A1(\V1/A3/A2/A1/M4/c1 ),
    .A2(\V1/A3/A2/A1/M4/c2 ),
    .ZN(\V1/A3/A2/c1 ));
 AND2_X1 \V1/A3/A2/A2/M1/M1/_0_  (.A1(\V1/v4 [12]),
    .A2(net6),
    .ZN(\V1/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M1/M1/_1_  (.A(\V1/v4 [12]),
    .B(net6),
    .Z(\V1/A3/A2/A2/M1/s1 ));
 AND2_X1 \V1/A3/A2/A2/M1/M2/_0_  (.A1(\V1/A3/A2/A2/M1/s1 ),
    .A2(\V1/A3/A2/c1 ),
    .ZN(\V1/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M1/M2/_1_  (.A(\V1/A3/A2/A2/M1/s1 ),
    .B(\V1/A3/A2/c1 ),
    .Z(v1[28]));
 OR2_X1 \V1/A3/A2/A2/M1/_0_  (.A1(\V1/A3/A2/A2/M1/c1 ),
    .A2(\V1/A3/A2/A2/M1/c2 ),
    .ZN(\V1/A3/A2/A2/c1 ));
 AND2_X1 \V1/A3/A2/A2/M2/M1/_0_  (.A1(\V1/v4 [13]),
    .A2(net6),
    .ZN(\V1/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M2/M1/_1_  (.A(\V1/v4 [13]),
    .B(net6),
    .Z(\V1/A3/A2/A2/M2/s1 ));
 AND2_X1 \V1/A3/A2/A2/M2/M2/_0_  (.A1(\V1/A3/A2/A2/M2/s1 ),
    .A2(\V1/A3/A2/A2/c1 ),
    .ZN(\V1/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M2/M2/_1_  (.A(\V1/A3/A2/A2/M2/s1 ),
    .B(\V1/A3/A2/A2/c1 ),
    .Z(v1[29]));
 OR2_X1 \V1/A3/A2/A2/M2/_0_  (.A1(\V1/A3/A2/A2/M2/c1 ),
    .A2(\V1/A3/A2/A2/M2/c2 ),
    .ZN(\V1/A3/A2/A2/c2 ));
 AND2_X1 \V1/A3/A2/A2/M3/M1/_0_  (.A1(\V1/v4 [14]),
    .A2(net6),
    .ZN(\V1/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M3/M1/_1_  (.A(\V1/v4 [14]),
    .B(net6),
    .Z(\V1/A3/A2/A2/M3/s1 ));
 AND2_X1 \V1/A3/A2/A2/M3/M2/_0_  (.A1(\V1/A3/A2/A2/M3/s1 ),
    .A2(\V1/A3/A2/A2/c2 ),
    .ZN(\V1/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M3/M2/_1_  (.A(\V1/A3/A2/A2/M3/s1 ),
    .B(\V1/A3/A2/A2/c2 ),
    .Z(v1[30]));
 OR2_X1 \V1/A3/A2/A2/M3/_0_  (.A1(\V1/A3/A2/A2/M3/c1 ),
    .A2(\V1/A3/A2/A2/M3/c2 ),
    .ZN(\V1/A3/A2/A2/c3 ));
 AND2_X1 \V1/A3/A2/A2/M4/M1/_0_  (.A1(\V1/v4 [15]),
    .A2(net6),
    .ZN(\V1/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V1/A3/A2/A2/M4/M1/_1_  (.A(\V1/v4 [15]),
    .B(net6),
    .Z(\V1/A3/A2/A2/M4/s1 ));
 AND2_X1 \V1/A3/A2/A2/M4/M2/_0_  (.A1(\V1/A3/A2/A2/M4/s1 ),
    .A2(\V1/A3/A2/A2/c3 ),
    .ZN(\V1/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V1/A3/A2/A2/M4/M2/_1_  (.A(\V1/A3/A2/A2/M4/s1 ),
    .B(\V1/A3/A2/A2/c3 ),
    .Z(v1[31]));
 OR2_X1 \V1/A3/A2/A2/M4/_0_  (.A1(\V1/A3/A2/A2/M4/c1 ),
    .A2(\V1/A3/A2/A2/M4/c2 ),
    .ZN(\V1/overflow ));
 AND2_X1 \V1/V1/A1/A1/M1/M1/_0_  (.A1(\V1/V1/v2 [0]),
    .A2(\V1/V1/v3 [0]),
    .ZN(\V1/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M1/M1/_1_  (.A(\V1/V1/v2 [0]),
    .B(\V1/V1/v3 [0]),
    .Z(\V1/V1/A1/A1/M1/s1 ));
 AND2_X1 \V1/V1/A1/A1/M1/M2/_0_  (.A1(\V1/V1/A1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M1/M2/_1_  (.A(\V1/V1/A1/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/s1 [0]));
 OR2_X1 \V1/V1/A1/A1/M1/_0_  (.A1(\V1/V1/A1/A1/M1/c1 ),
    .A2(\V1/V1/A1/A1/M1/c2 ),
    .ZN(\V1/V1/A1/A1/c1 ));
 AND2_X1 \V1/V1/A1/A1/M2/M1/_0_  (.A1(\V1/V1/v2 [1]),
    .A2(\V1/V1/v3 [1]),
    .ZN(\V1/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M2/M1/_1_  (.A(\V1/V1/v2 [1]),
    .B(\V1/V1/v3 [1]),
    .Z(\V1/V1/A1/A1/M2/s1 ));
 AND2_X1 \V1/V1/A1/A1/M2/M2/_0_  (.A1(\V1/V1/A1/A1/M2/s1 ),
    .A2(\V1/V1/A1/A1/c1 ),
    .ZN(\V1/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M2/M2/_1_  (.A(\V1/V1/A1/A1/M2/s1 ),
    .B(\V1/V1/A1/A1/c1 ),
    .Z(\V1/V1/s1 [1]));
 OR2_X1 \V1/V1/A1/A1/M2/_0_  (.A1(\V1/V1/A1/A1/M2/c1 ),
    .A2(\V1/V1/A1/A1/M2/c2 ),
    .ZN(\V1/V1/A1/A1/c2 ));
 AND2_X1 \V1/V1/A1/A1/M3/M1/_0_  (.A1(\V1/V1/v2 [2]),
    .A2(\V1/V1/v3 [2]),
    .ZN(\V1/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M3/M1/_1_  (.A(\V1/V1/v2 [2]),
    .B(\V1/V1/v3 [2]),
    .Z(\V1/V1/A1/A1/M3/s1 ));
 AND2_X1 \V1/V1/A1/A1/M3/M2/_0_  (.A1(\V1/V1/A1/A1/M3/s1 ),
    .A2(\V1/V1/A1/A1/c2 ),
    .ZN(\V1/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M3/M2/_1_  (.A(\V1/V1/A1/A1/M3/s1 ),
    .B(\V1/V1/A1/A1/c2 ),
    .Z(\V1/V1/s1 [2]));
 OR2_X1 \V1/V1/A1/A1/M3/_0_  (.A1(\V1/V1/A1/A1/M3/c1 ),
    .A2(\V1/V1/A1/A1/M3/c2 ),
    .ZN(\V1/V1/A1/A1/c3 ));
 AND2_X1 \V1/V1/A1/A1/M4/M1/_0_  (.A1(\V1/V1/v2 [3]),
    .A2(\V1/V1/v3 [3]),
    .ZN(\V1/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A1/A1/M4/M1/_1_  (.A(\V1/V1/v2 [3]),
    .B(\V1/V1/v3 [3]),
    .Z(\V1/V1/A1/A1/M4/s1 ));
 AND2_X1 \V1/V1/A1/A1/M4/M2/_0_  (.A1(\V1/V1/A1/A1/M4/s1 ),
    .A2(\V1/V1/A1/A1/c3 ),
    .ZN(\V1/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V1/A1/A1/M4/M2/_1_  (.A(\V1/V1/A1/A1/M4/s1 ),
    .B(\V1/V1/A1/A1/c3 ),
    .Z(\V1/V1/s1 [3]));
 OR2_X1 \V1/V1/A1/A1/M4/_0_  (.A1(\V1/V1/A1/A1/M4/c1 ),
    .A2(\V1/V1/A1/A1/M4/c2 ),
    .ZN(\V1/V1/A1/c1 ));
 AND2_X1 \V1/V1/A1/A2/M1/M1/_0_  (.A1(\V1/V1/v2 [4]),
    .A2(\V1/V1/v3 [4]),
    .ZN(\V1/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M1/M1/_1_  (.A(\V1/V1/v2 [4]),
    .B(\V1/V1/v3 [4]),
    .Z(\V1/V1/A1/A2/M1/s1 ));
 AND2_X1 \V1/V1/A1/A2/M1/M2/_0_  (.A1(\V1/V1/A1/A2/M1/s1 ),
    .A2(\V1/V1/A1/c1 ),
    .ZN(\V1/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M1/M2/_1_  (.A(\V1/V1/A1/A2/M1/s1 ),
    .B(\V1/V1/A1/c1 ),
    .Z(\V1/V1/s1 [4]));
 OR2_X1 \V1/V1/A1/A2/M1/_0_  (.A1(\V1/V1/A1/A2/M1/c1 ),
    .A2(\V1/V1/A1/A2/M1/c2 ),
    .ZN(\V1/V1/A1/A2/c1 ));
 AND2_X1 \V1/V1/A1/A2/M2/M1/_0_  (.A1(\V1/V1/v2 [5]),
    .A2(\V1/V1/v3 [5]),
    .ZN(\V1/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M2/M1/_1_  (.A(\V1/V1/v2 [5]),
    .B(\V1/V1/v3 [5]),
    .Z(\V1/V1/A1/A2/M2/s1 ));
 AND2_X1 \V1/V1/A1/A2/M2/M2/_0_  (.A1(\V1/V1/A1/A2/M2/s1 ),
    .A2(\V1/V1/A1/A2/c1 ),
    .ZN(\V1/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M2/M2/_1_  (.A(\V1/V1/A1/A2/M2/s1 ),
    .B(\V1/V1/A1/A2/c1 ),
    .Z(\V1/V1/s1 [5]));
 OR2_X1 \V1/V1/A1/A2/M2/_0_  (.A1(\V1/V1/A1/A2/M2/c1 ),
    .A2(\V1/V1/A1/A2/M2/c2 ),
    .ZN(\V1/V1/A1/A2/c2 ));
 AND2_X1 \V1/V1/A1/A2/M3/M1/_0_  (.A1(\V1/V1/v2 [6]),
    .A2(\V1/V1/v3 [6]),
    .ZN(\V1/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M3/M1/_1_  (.A(\V1/V1/v2 [6]),
    .B(\V1/V1/v3 [6]),
    .Z(\V1/V1/A1/A2/M3/s1 ));
 AND2_X1 \V1/V1/A1/A2/M3/M2/_0_  (.A1(\V1/V1/A1/A2/M3/s1 ),
    .A2(\V1/V1/A1/A2/c2 ),
    .ZN(\V1/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M3/M2/_1_  (.A(\V1/V1/A1/A2/M3/s1 ),
    .B(\V1/V1/A1/A2/c2 ),
    .Z(\V1/V1/s1 [6]));
 OR2_X1 \V1/V1/A1/A2/M3/_0_  (.A1(\V1/V1/A1/A2/M3/c1 ),
    .A2(\V1/V1/A1/A2/M3/c2 ),
    .ZN(\V1/V1/A1/A2/c3 ));
 AND2_X1 \V1/V1/A1/A2/M4/M1/_0_  (.A1(\V1/V1/v2 [7]),
    .A2(\V1/V1/v3 [7]),
    .ZN(\V1/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A1/A2/M4/M1/_1_  (.A(\V1/V1/v2 [7]),
    .B(\V1/V1/v3 [7]),
    .Z(\V1/V1/A1/A2/M4/s1 ));
 AND2_X1 \V1/V1/A1/A2/M4/M2/_0_  (.A1(\V1/V1/A1/A2/M4/s1 ),
    .A2(\V1/V1/A1/A2/c3 ),
    .ZN(\V1/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A1/A2/M4/M2/_1_  (.A(\V1/V1/A1/A2/M4/s1 ),
    .B(\V1/V1/A1/A2/c3 ),
    .Z(\V1/V1/s1 [7]));
 OR2_X1 \V1/V1/A1/A2/M4/_0_  (.A1(\V1/V1/A1/A2/M4/c1 ),
    .A2(\V1/V1/A1/A2/M4/c2 ),
    .ZN(\V1/V1/c1 ));
 AND2_X1 \V1/V1/A2/A1/M1/M1/_0_  (.A1(\V1/V1/s1 [0]),
    .A2(\V1/V1/v1 [4]),
    .ZN(\V1/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M1/M1/_1_  (.A(\V1/V1/s1 [0]),
    .B(\V1/V1/v1 [4]),
    .Z(\V1/V1/A2/A1/M1/s1 ));
 AND2_X1 \V1/V1/A2/A1/M1/M2/_0_  (.A1(\V1/V1/A2/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V1/A2/A1/M1/M2/_1_  (.A(\V1/V1/A2/A1/M1/s1 ),
    .B(net4),
    .Z(v1[4]));
 OR2_X1 \V1/V1/A2/A1/M1/_0_  (.A1(\V1/V1/A2/A1/M1/c1 ),
    .A2(\V1/V1/A2/A1/M1/c2 ),
    .ZN(\V1/V1/A2/A1/c1 ));
 AND2_X1 \V1/V1/A2/A1/M2/M1/_0_  (.A1(\V1/V1/s1 [1]),
    .A2(\V1/V1/v1 [5]),
    .ZN(\V1/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M2/M1/_1_  (.A(\V1/V1/s1 [1]),
    .B(\V1/V1/v1 [5]),
    .Z(\V1/V1/A2/A1/M2/s1 ));
 AND2_X1 \V1/V1/A2/A1/M2/M2/_0_  (.A1(\V1/V1/A2/A1/M2/s1 ),
    .A2(\V1/V1/A2/A1/c1 ),
    .ZN(\V1/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V1/A2/A1/M2/M2/_1_  (.A(\V1/V1/A2/A1/M2/s1 ),
    .B(\V1/V1/A2/A1/c1 ),
    .Z(v1[5]));
 OR2_X1 \V1/V1/A2/A1/M2/_0_  (.A1(\V1/V1/A2/A1/M2/c1 ),
    .A2(\V1/V1/A2/A1/M2/c2 ),
    .ZN(\V1/V1/A2/A1/c2 ));
 AND2_X1 \V1/V1/A2/A1/M3/M1/_0_  (.A1(\V1/V1/s1 [2]),
    .A2(\V1/V1/v1 [6]),
    .ZN(\V1/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M3/M1/_1_  (.A(\V1/V1/s1 [2]),
    .B(\V1/V1/v1 [6]),
    .Z(\V1/V1/A2/A1/M3/s1 ));
 AND2_X1 \V1/V1/A2/A1/M3/M2/_0_  (.A1(\V1/V1/A2/A1/M3/s1 ),
    .A2(\V1/V1/A2/A1/c2 ),
    .ZN(\V1/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V1/A2/A1/M3/M2/_1_  (.A(\V1/V1/A2/A1/M3/s1 ),
    .B(\V1/V1/A2/A1/c2 ),
    .Z(v1[6]));
 OR2_X1 \V1/V1/A2/A1/M3/_0_  (.A1(\V1/V1/A2/A1/M3/c1 ),
    .A2(\V1/V1/A2/A1/M3/c2 ),
    .ZN(\V1/V1/A2/A1/c3 ));
 AND2_X1 \V1/V1/A2/A1/M4/M1/_0_  (.A1(\V1/V1/s1 [3]),
    .A2(\V1/V1/v1 [7]),
    .ZN(\V1/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A2/A1/M4/M1/_1_  (.A(\V1/V1/s1 [3]),
    .B(\V1/V1/v1 [7]),
    .Z(\V1/V1/A2/A1/M4/s1 ));
 AND2_X1 \V1/V1/A2/A1/M4/M2/_0_  (.A1(\V1/V1/A2/A1/M4/s1 ),
    .A2(\V1/V1/A2/A1/c3 ),
    .ZN(\V1/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V1/A2/A1/M4/M2/_1_  (.A(\V1/V1/A2/A1/M4/s1 ),
    .B(\V1/V1/A2/A1/c3 ),
    .Z(v1[7]));
 OR2_X1 \V1/V1/A2/A1/M4/_0_  (.A1(\V1/V1/A2/A1/M4/c1 ),
    .A2(\V1/V1/A2/A1/M4/c2 ),
    .ZN(\V1/V1/A2/c1 ));
 AND2_X1 \V1/V1/A2/A2/M1/M1/_0_  (.A1(\V1/V1/s1 [4]),
    .A2(net4),
    .ZN(\V1/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M1/M1/_1_  (.A(\V1/V1/s1 [4]),
    .B(net4),
    .Z(\V1/V1/A2/A2/M1/s1 ));
 AND2_X1 \V1/V1/A2/A2/M1/M2/_0_  (.A1(\V1/V1/A2/A2/M1/s1 ),
    .A2(\V1/V1/A2/c1 ),
    .ZN(\V1/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M1/M2/_1_  (.A(\V1/V1/A2/A2/M1/s1 ),
    .B(\V1/V1/A2/c1 ),
    .Z(\V1/V1/s2 [4]));
 OR2_X1 \V1/V1/A2/A2/M1/_0_  (.A1(\V1/V1/A2/A2/M1/c1 ),
    .A2(\V1/V1/A2/A2/M1/c2 ),
    .ZN(\V1/V1/A2/A2/c1 ));
 AND2_X1 \V1/V1/A2/A2/M2/M1/_0_  (.A1(\V1/V1/s1 [5]),
    .A2(net4),
    .ZN(\V1/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M2/M1/_1_  (.A(\V1/V1/s1 [5]),
    .B(net4),
    .Z(\V1/V1/A2/A2/M2/s1 ));
 AND2_X1 \V1/V1/A2/A2/M2/M2/_0_  (.A1(\V1/V1/A2/A2/M2/s1 ),
    .A2(\V1/V1/A2/A2/c1 ),
    .ZN(\V1/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M2/M2/_1_  (.A(\V1/V1/A2/A2/M2/s1 ),
    .B(\V1/V1/A2/A2/c1 ),
    .Z(\V1/V1/s2 [5]));
 OR2_X1 \V1/V1/A2/A2/M2/_0_  (.A1(\V1/V1/A2/A2/M2/c1 ),
    .A2(\V1/V1/A2/A2/M2/c2 ),
    .ZN(\V1/V1/A2/A2/c2 ));
 AND2_X1 \V1/V1/A2/A2/M3/M1/_0_  (.A1(\V1/V1/s1 [6]),
    .A2(net4),
    .ZN(\V1/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M3/M1/_1_  (.A(\V1/V1/s1 [6]),
    .B(net4),
    .Z(\V1/V1/A2/A2/M3/s1 ));
 AND2_X1 \V1/V1/A2/A2/M3/M2/_0_  (.A1(\V1/V1/A2/A2/M3/s1 ),
    .A2(\V1/V1/A2/A2/c2 ),
    .ZN(\V1/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M3/M2/_1_  (.A(\V1/V1/A2/A2/M3/s1 ),
    .B(\V1/V1/A2/A2/c2 ),
    .Z(\V1/V1/s2 [6]));
 OR2_X1 \V1/V1/A2/A2/M3/_0_  (.A1(\V1/V1/A2/A2/M3/c1 ),
    .A2(\V1/V1/A2/A2/M3/c2 ),
    .ZN(\V1/V1/A2/A2/c3 ));
 AND2_X1 \V1/V1/A2/A2/M4/M1/_0_  (.A1(\V1/V1/s1 [7]),
    .A2(net4),
    .ZN(\V1/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A2/A2/M4/M1/_1_  (.A(\V1/V1/s1 [7]),
    .B(net4),
    .Z(\V1/V1/A2/A2/M4/s1 ));
 AND2_X1 \V1/V1/A2/A2/M4/M2/_0_  (.A1(\V1/V1/A2/A2/M4/s1 ),
    .A2(\V1/V1/A2/A2/c3 ),
    .ZN(\V1/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A2/A2/M4/M2/_1_  (.A(\V1/V1/A2/A2/M4/s1 ),
    .B(\V1/V1/A2/A2/c3 ),
    .Z(\V1/V1/s2 [7]));
 OR2_X1 \V1/V1/A2/A2/M4/_0_  (.A1(\V1/V1/A2/A2/M4/c1 ),
    .A2(\V1/V1/A2/A2/M4/c2 ),
    .ZN(\V1/V1/c2 ));
 AND2_X1 \V1/V1/A3/A1/M1/M1/_0_  (.A1(\V1/V1/v4 [0]),
    .A2(\V1/V1/s2 [4]),
    .ZN(\V1/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M1/M1/_1_  (.A(\V1/V1/v4 [0]),
    .B(\V1/V1/s2 [4]),
    .Z(\V1/V1/A3/A1/M1/s1 ));
 AND2_X1 \V1/V1/A3/A1/M1/M2/_0_  (.A1(\V1/V1/A3/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M1/M2/_1_  (.A(\V1/V1/A3/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/v1 [8]));
 OR2_X1 \V1/V1/A3/A1/M1/_0_  (.A1(\V1/V1/A3/A1/M1/c1 ),
    .A2(\V1/V1/A3/A1/M1/c2 ),
    .ZN(\V1/V1/A3/A1/c1 ));
 AND2_X1 \V1/V1/A3/A1/M2/M1/_0_  (.A1(\V1/V1/v4 [1]),
    .A2(\V1/V1/s2 [5]),
    .ZN(\V1/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M2/M1/_1_  (.A(\V1/V1/v4 [1]),
    .B(\V1/V1/s2 [5]),
    .Z(\V1/V1/A3/A1/M2/s1 ));
 AND2_X1 \V1/V1/A3/A1/M2/M2/_0_  (.A1(\V1/V1/A3/A1/M2/s1 ),
    .A2(\V1/V1/A3/A1/c1 ),
    .ZN(\V1/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M2/M2/_1_  (.A(\V1/V1/A3/A1/M2/s1 ),
    .B(\V1/V1/A3/A1/c1 ),
    .Z(\V1/v1 [9]));
 OR2_X1 \V1/V1/A3/A1/M2/_0_  (.A1(\V1/V1/A3/A1/M2/c1 ),
    .A2(\V1/V1/A3/A1/M2/c2 ),
    .ZN(\V1/V1/A3/A1/c2 ));
 AND2_X1 \V1/V1/A3/A1/M3/M1/_0_  (.A1(\V1/V1/v4 [2]),
    .A2(\V1/V1/s2 [6]),
    .ZN(\V1/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M3/M1/_1_  (.A(\V1/V1/v4 [2]),
    .B(\V1/V1/s2 [6]),
    .Z(\V1/V1/A3/A1/M3/s1 ));
 AND2_X1 \V1/V1/A3/A1/M3/M2/_0_  (.A1(\V1/V1/A3/A1/M3/s1 ),
    .A2(\V1/V1/A3/A1/c2 ),
    .ZN(\V1/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M3/M2/_1_  (.A(\V1/V1/A3/A1/M3/s1 ),
    .B(\V1/V1/A3/A1/c2 ),
    .Z(\V1/v1 [10]));
 OR2_X1 \V1/V1/A3/A1/M3/_0_  (.A1(\V1/V1/A3/A1/M3/c1 ),
    .A2(\V1/V1/A3/A1/M3/c2 ),
    .ZN(\V1/V1/A3/A1/c3 ));
 AND2_X1 \V1/V1/A3/A1/M4/M1/_0_  (.A1(\V1/V1/v4 [3]),
    .A2(\V1/V1/s2 [7]),
    .ZN(\V1/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V1/A3/A1/M4/M1/_1_  (.A(\V1/V1/v4 [3]),
    .B(\V1/V1/s2 [7]),
    .Z(\V1/V1/A3/A1/M4/s1 ));
 AND2_X1 \V1/V1/A3/A1/M4/M2/_0_  (.A1(\V1/V1/A3/A1/M4/s1 ),
    .A2(\V1/V1/A3/A1/c3 ),
    .ZN(\V1/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V1/A3/A1/M4/M2/_1_  (.A(\V1/V1/A3/A1/M4/s1 ),
    .B(\V1/V1/A3/A1/c3 ),
    .Z(\V1/v1 [11]));
 OR2_X1 \V1/V1/A3/A1/M4/_0_  (.A1(\V1/V1/A3/A1/M4/c1 ),
    .A2(\V1/V1/A3/A1/M4/c2 ),
    .ZN(\V1/V1/A3/c1 ));
 AND2_X1 \V1/V1/A3/A2/M1/M1/_0_  (.A1(\V1/V1/v4 [4]),
    .A2(\V1/V1/c3 ),
    .ZN(\V1/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M1/M1/_1_  (.A(\V1/V1/v4 [4]),
    .B(\V1/V1/c3 ),
    .Z(\V1/V1/A3/A2/M1/s1 ));
 AND2_X1 \V1/V1/A3/A2/M1/M2/_0_  (.A1(\V1/V1/A3/A2/M1/s1 ),
    .A2(\V1/V1/A3/c1 ),
    .ZN(\V1/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M1/M2/_1_  (.A(\V1/V1/A3/A2/M1/s1 ),
    .B(\V1/V1/A3/c1 ),
    .Z(\V1/v1 [12]));
 OR2_X1 \V1/V1/A3/A2/M1/_0_  (.A1(\V1/V1/A3/A2/M1/c1 ),
    .A2(\V1/V1/A3/A2/M1/c2 ),
    .ZN(\V1/V1/A3/A2/c1 ));
 AND2_X1 \V1/V1/A3/A2/M2/M1/_0_  (.A1(\V1/V1/v4 [5]),
    .A2(net4),
    .ZN(\V1/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M2/M1/_1_  (.A(\V1/V1/v4 [5]),
    .B(net4),
    .Z(\V1/V1/A3/A2/M2/s1 ));
 AND2_X1 \V1/V1/A3/A2/M2/M2/_0_  (.A1(\V1/V1/A3/A2/M2/s1 ),
    .A2(\V1/V1/A3/A2/c1 ),
    .ZN(\V1/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M2/M2/_1_  (.A(\V1/V1/A3/A2/M2/s1 ),
    .B(\V1/V1/A3/A2/c1 ),
    .Z(\V1/v1 [13]));
 OR2_X1 \V1/V1/A3/A2/M2/_0_  (.A1(\V1/V1/A3/A2/M2/c1 ),
    .A2(\V1/V1/A3/A2/M2/c2 ),
    .ZN(\V1/V1/A3/A2/c2 ));
 AND2_X1 \V1/V1/A3/A2/M3/M1/_0_  (.A1(\V1/V1/v4 [6]),
    .A2(net4),
    .ZN(\V1/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M3/M1/_1_  (.A(\V1/V1/v4 [6]),
    .B(net4),
    .Z(\V1/V1/A3/A2/M3/s1 ));
 AND2_X1 \V1/V1/A3/A2/M3/M2/_0_  (.A1(\V1/V1/A3/A2/M3/s1 ),
    .A2(\V1/V1/A3/A2/c2 ),
    .ZN(\V1/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M3/M2/_1_  (.A(\V1/V1/A3/A2/M3/s1 ),
    .B(\V1/V1/A3/A2/c2 ),
    .Z(\V1/v1 [14]));
 OR2_X1 \V1/V1/A3/A2/M3/_0_  (.A1(\V1/V1/A3/A2/M3/c1 ),
    .A2(\V1/V1/A3/A2/M3/c2 ),
    .ZN(\V1/V1/A3/A2/c3 ));
 AND2_X1 \V1/V1/A3/A2/M4/M1/_0_  (.A1(\V1/V1/v4 [7]),
    .A2(net4),
    .ZN(\V1/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V1/A3/A2/M4/M1/_1_  (.A(\V1/V1/v4 [7]),
    .B(net4),
    .Z(\V1/V1/A3/A2/M4/s1 ));
 AND2_X1 \V1/V1/A3/A2/M4/M2/_0_  (.A1(\V1/V1/A3/A2/M4/s1 ),
    .A2(\V1/V1/A3/A2/c3 ),
    .ZN(\V1/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V1/A3/A2/M4/M2/_1_  (.A(\V1/V1/A3/A2/M4/s1 ),
    .B(\V1/V1/A3/A2/c3 ),
    .Z(\V1/v1 [15]));
 OR2_X1 \V1/V1/A3/A2/M4/_0_  (.A1(\V1/V1/A3/A2/M4/c1 ),
    .A2(\V1/V1/A3/A2/M4/c2 ),
    .ZN(\V1/V1/overflow ));
 AND2_X1 \V1/V1/V1/A1/M1/M1/_0_  (.A1(\V1/V1/V1/v2 [0]),
    .A2(\V1/V1/V1/v3 [0]),
    .ZN(\V1/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M1/M1/_1_  (.A(\V1/V1/V1/v2 [0]),
    .B(\V1/V1/V1/v3 [0]),
    .Z(\V1/V1/V1/A1/M1/s1 ));
 AND2_X1 \V1/V1/V1/A1/M1/M2/_0_  (.A1(\V1/V1/V1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M1/M2/_1_  (.A(\V1/V1/V1/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/V1/s1 [0]));
 OR2_X1 \V1/V1/V1/A1/M1/_0_  (.A1(\V1/V1/V1/A1/M1/c1 ),
    .A2(\V1/V1/V1/A1/M1/c2 ),
    .ZN(\V1/V1/V1/A1/c1 ));
 AND2_X1 \V1/V1/V1/A1/M2/M1/_0_  (.A1(\V1/V1/V1/v2 [1]),
    .A2(\V1/V1/V1/v3 [1]),
    .ZN(\V1/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M2/M1/_1_  (.A(\V1/V1/V1/v2 [1]),
    .B(\V1/V1/V1/v3 [1]),
    .Z(\V1/V1/V1/A1/M2/s1 ));
 AND2_X1 \V1/V1/V1/A1/M2/M2/_0_  (.A1(\V1/V1/V1/A1/M2/s1 ),
    .A2(\V1/V1/V1/A1/c1 ),
    .ZN(\V1/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M2/M2/_1_  (.A(\V1/V1/V1/A1/M2/s1 ),
    .B(\V1/V1/V1/A1/c1 ),
    .Z(\V1/V1/V1/s1 [1]));
 OR2_X1 \V1/V1/V1/A1/M2/_0_  (.A1(\V1/V1/V1/A1/M2/c1 ),
    .A2(\V1/V1/V1/A1/M2/c2 ),
    .ZN(\V1/V1/V1/A1/c2 ));
 AND2_X1 \V1/V1/V1/A1/M3/M1/_0_  (.A1(\V1/V1/V1/v2 [2]),
    .A2(\V1/V1/V1/v3 [2]),
    .ZN(\V1/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M3/M1/_1_  (.A(\V1/V1/V1/v2 [2]),
    .B(\V1/V1/V1/v3 [2]),
    .Z(\V1/V1/V1/A1/M3/s1 ));
 AND2_X1 \V1/V1/V1/A1/M3/M2/_0_  (.A1(\V1/V1/V1/A1/M3/s1 ),
    .A2(\V1/V1/V1/A1/c2 ),
    .ZN(\V1/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M3/M2/_1_  (.A(\V1/V1/V1/A1/M3/s1 ),
    .B(\V1/V1/V1/A1/c2 ),
    .Z(\V1/V1/V1/s1 [2]));
 OR2_X1 \V1/V1/V1/A1/M3/_0_  (.A1(\V1/V1/V1/A1/M3/c1 ),
    .A2(\V1/V1/V1/A1/M3/c2 ),
    .ZN(\V1/V1/V1/A1/c3 ));
 AND2_X1 \V1/V1/V1/A1/M4/M1/_0_  (.A1(\V1/V1/V1/v2 [3]),
    .A2(\V1/V1/V1/v3 [3]),
    .ZN(\V1/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A1/M4/M1/_1_  (.A(\V1/V1/V1/v2 [3]),
    .B(\V1/V1/V1/v3 [3]),
    .Z(\V1/V1/V1/A1/M4/s1 ));
 AND2_X1 \V1/V1/V1/A1/M4/M2/_0_  (.A1(\V1/V1/V1/A1/M4/s1 ),
    .A2(\V1/V1/V1/A1/c3 ),
    .ZN(\V1/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A1/M4/M2/_1_  (.A(\V1/V1/V1/A1/M4/s1 ),
    .B(\V1/V1/V1/A1/c3 ),
    .Z(\V1/V1/V1/s1 [3]));
 OR2_X1 \V1/V1/V1/A1/M4/_0_  (.A1(\V1/V1/V1/A1/M4/c1 ),
    .A2(\V1/V1/V1/A1/M4/c2 ),
    .ZN(\V1/V1/V1/c1 ));
 AND2_X1 \V1/V1/V1/A2/M1/M1/_0_  (.A1(\V1/V1/V1/s1 [0]),
    .A2(\V1/V1/V1/v1 [2]),
    .ZN(\V1/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M1/M1/_1_  (.A(\V1/V1/V1/s1 [0]),
    .B(\V1/V1/V1/v1 [2]),
    .Z(\V1/V1/V1/A2/M1/s1 ));
 AND2_X1 \V1/V1/V1/A2/M1/M2/_0_  (.A1(\V1/V1/V1/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M1/M2/_1_  (.A(\V1/V1/V1/A2/M1/s1 ),
    .B(net4),
    .Z(v1[2]));
 OR2_X1 \V1/V1/V1/A2/M1/_0_  (.A1(\V1/V1/V1/A2/M1/c1 ),
    .A2(\V1/V1/V1/A2/M1/c2 ),
    .ZN(\V1/V1/V1/A2/c1 ));
 AND2_X1 \V1/V1/V1/A2/M2/M1/_0_  (.A1(\V1/V1/V1/s1 [1]),
    .A2(\V1/V1/V1/v1 [3]),
    .ZN(\V1/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M2/M1/_1_  (.A(\V1/V1/V1/s1 [1]),
    .B(\V1/V1/V1/v1 [3]),
    .Z(\V1/V1/V1/A2/M2/s1 ));
 AND2_X1 \V1/V1/V1/A2/M2/M2/_0_  (.A1(\V1/V1/V1/A2/M2/s1 ),
    .A2(\V1/V1/V1/A2/c1 ),
    .ZN(\V1/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M2/M2/_1_  (.A(\V1/V1/V1/A2/M2/s1 ),
    .B(\V1/V1/V1/A2/c1 ),
    .Z(v1[3]));
 OR2_X1 \V1/V1/V1/A2/M2/_0_  (.A1(\V1/V1/V1/A2/M2/c1 ),
    .A2(\V1/V1/V1/A2/M2/c2 ),
    .ZN(\V1/V1/V1/A2/c2 ));
 AND2_X1 \V1/V1/V1/A2/M3/M1/_0_  (.A1(\V1/V1/V1/s1 [2]),
    .A2(net4),
    .ZN(\V1/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M3/M1/_1_  (.A(\V1/V1/V1/s1 [2]),
    .B(net4),
    .Z(\V1/V1/V1/A2/M3/s1 ));
 AND2_X1 \V1/V1/V1/A2/M3/M2/_0_  (.A1(\V1/V1/V1/A2/M3/s1 ),
    .A2(\V1/V1/V1/A2/c2 ),
    .ZN(\V1/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M3/M2/_1_  (.A(\V1/V1/V1/A2/M3/s1 ),
    .B(\V1/V1/V1/A2/c2 ),
    .Z(\V1/V1/V1/s2 [2]));
 OR2_X1 \V1/V1/V1/A2/M3/_0_  (.A1(\V1/V1/V1/A2/M3/c1 ),
    .A2(\V1/V1/V1/A2/M3/c2 ),
    .ZN(\V1/V1/V1/A2/c3 ));
 AND2_X1 \V1/V1/V1/A2/M4/M1/_0_  (.A1(\V1/V1/V1/s1 [3]),
    .A2(net4),
    .ZN(\V1/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A2/M4/M1/_1_  (.A(\V1/V1/V1/s1 [3]),
    .B(net4),
    .Z(\V1/V1/V1/A2/M4/s1 ));
 AND2_X1 \V1/V1/V1/A2/M4/M2/_0_  (.A1(\V1/V1/V1/A2/M4/s1 ),
    .A2(\V1/V1/V1/A2/c3 ),
    .ZN(\V1/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A2/M4/M2/_1_  (.A(\V1/V1/V1/A2/M4/s1 ),
    .B(\V1/V1/V1/A2/c3 ),
    .Z(\V1/V1/V1/s2 [3]));
 OR2_X1 \V1/V1/V1/A2/M4/_0_  (.A1(\V1/V1/V1/A2/M4/c1 ),
    .A2(\V1/V1/V1/A2/M4/c2 ),
    .ZN(\V1/V1/V1/c2 ));
 AND2_X1 \V1/V1/V1/A3/M1/M1/_0_  (.A1(\V1/V1/V1/v4 [0]),
    .A2(\V1/V1/V1/s2 [2]),
    .ZN(\V1/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M1/M1/_1_  (.A(\V1/V1/V1/v4 [0]),
    .B(\V1/V1/V1/s2 [2]),
    .Z(\V1/V1/V1/A3/M1/s1 ));
 AND2_X1 \V1/V1/V1/A3/M1/M2/_0_  (.A1(\V1/V1/V1/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M1/M2/_1_  (.A(\V1/V1/V1/A3/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/v1 [4]));
 OR2_X1 \V1/V1/V1/A3/M1/_0_  (.A1(\V1/V1/V1/A3/M1/c1 ),
    .A2(\V1/V1/V1/A3/M1/c2 ),
    .ZN(\V1/V1/V1/A3/c1 ));
 AND2_X1 \V1/V1/V1/A3/M2/M1/_0_  (.A1(\V1/V1/V1/v4 [1]),
    .A2(\V1/V1/V1/s2 [3]),
    .ZN(\V1/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M2/M1/_1_  (.A(\V1/V1/V1/v4 [1]),
    .B(\V1/V1/V1/s2 [3]),
    .Z(\V1/V1/V1/A3/M2/s1 ));
 AND2_X1 \V1/V1/V1/A3/M2/M2/_0_  (.A1(\V1/V1/V1/A3/M2/s1 ),
    .A2(\V1/V1/V1/A3/c1 ),
    .ZN(\V1/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M2/M2/_1_  (.A(\V1/V1/V1/A3/M2/s1 ),
    .B(\V1/V1/V1/A3/c1 ),
    .Z(\V1/V1/v1 [5]));
 OR2_X1 \V1/V1/V1/A3/M2/_0_  (.A1(\V1/V1/V1/A3/M2/c1 ),
    .A2(\V1/V1/V1/A3/M2/c2 ),
    .ZN(\V1/V1/V1/A3/c2 ));
 AND2_X1 \V1/V1/V1/A3/M3/M1/_0_  (.A1(\V1/V1/V1/v4 [2]),
    .A2(\V1/V1/V1/c3 ),
    .ZN(\V1/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M3/M1/_1_  (.A(\V1/V1/V1/v4 [2]),
    .B(\V1/V1/V1/c3 ),
    .Z(\V1/V1/V1/A3/M3/s1 ));
 AND2_X1 \V1/V1/V1/A3/M3/M2/_0_  (.A1(\V1/V1/V1/A3/M3/s1 ),
    .A2(\V1/V1/V1/A3/c2 ),
    .ZN(\V1/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M3/M2/_1_  (.A(\V1/V1/V1/A3/M3/s1 ),
    .B(\V1/V1/V1/A3/c2 ),
    .Z(\V1/V1/v1 [6]));
 OR2_X1 \V1/V1/V1/A3/M3/_0_  (.A1(\V1/V1/V1/A3/M3/c1 ),
    .A2(\V1/V1/V1/A3/M3/c2 ),
    .ZN(\V1/V1/V1/A3/c3 ));
 AND2_X1 \V1/V1/V1/A3/M4/M1/_0_  (.A1(\V1/V1/V1/v4 [3]),
    .A2(net4),
    .ZN(\V1/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V1/A3/M4/M1/_1_  (.A(\V1/V1/V1/v4 [3]),
    .B(net4),
    .Z(\V1/V1/V1/A3/M4/s1 ));
 AND2_X1 \V1/V1/V1/A3/M4/M2/_0_  (.A1(\V1/V1/V1/A3/M4/s1 ),
    .A2(\V1/V1/V1/A3/c3 ),
    .ZN(\V1/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V1/A3/M4/M2/_1_  (.A(\V1/V1/V1/A3/M4/s1 ),
    .B(\V1/V1/V1/A3/c3 ),
    .Z(\V1/V1/v1 [7]));
 OR2_X1 \V1/V1/V1/A3/M4/_0_  (.A1(\V1/V1/V1/A3/M4/c1 ),
    .A2(\V1/V1/V1/A3/M4/c2 ),
    .ZN(\V1/V1/V1/overflow ));
 AND2_X1 \V1/V1/V1/V1/HA1/_0_  (.A1(\V1/V1/V1/V1/w2 ),
    .A2(\V1/V1/V1/V1/w1 ),
    .ZN(\V1/V1/V1/V1/w4 ));
 XOR2_X2 \V1/V1/V1/V1/HA1/_1_  (.A(\V1/V1/V1/V1/w2 ),
    .B(\V1/V1/V1/V1/w1 ),
    .Z(v1[1]));
 AND2_X1 \V1/V1/V1/V1/HA2/_0_  (.A1(\V1/V1/V1/V1/w4 ),
    .A2(\V1/V1/V1/V1/w3 ),
    .ZN(\V1/V1/V1/v1 [3]));
 XOR2_X2 \V1/V1/V1/V1/HA2/_1_  (.A(\V1/V1/V1/V1/w4 ),
    .B(\V1/V1/V1/V1/w3 ),
    .Z(\V1/V1/V1/v1 [2]));
 AND2_X2 \V1/V1/V1/V1/_0_  (.A1(A[0]),
    .A2(net23),
    .ZN(v1[0]));
 AND2_X1 \V1/V1/V1/V1/_1_  (.A1(net48),
    .A2(B[1]),
    .ZN(\V1/V1/V1/V1/w1 ));
 AND2_X1 \V1/V1/V1/V1/_2_  (.A1(net23),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V1/w2 ));
 AND2_X1 \V1/V1/V1/V1/_3_  (.A1(B[1]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V1/w3 ));
 AND2_X1 \V1/V1/V1/V2/HA1/_0_  (.A1(\V1/V1/V1/V2/w2 ),
    .A2(\V1/V1/V1/V2/w1 ),
    .ZN(\V1/V1/V1/V2/w4 ));
 XOR2_X2 \V1/V1/V1/V2/HA1/_1_  (.A(\V1/V1/V1/V2/w2 ),
    .B(\V1/V1/V1/V2/w1 ),
    .Z(\V1/V1/V1/v2 [1]));
 AND2_X1 \V1/V1/V1/V2/HA2/_0_  (.A1(\V1/V1/V1/V2/w4 ),
    .A2(\V1/V1/V1/V2/w3 ),
    .ZN(\V1/V1/V1/v2 [3]));
 XOR2_X2 \V1/V1/V1/V2/HA2/_1_  (.A(\V1/V1/V1/V2/w4 ),
    .B(\V1/V1/V1/V2/w3 ),
    .Z(\V1/V1/V1/v2 [2]));
 AND2_X1 \V1/V1/V1/V2/_0_  (.A1(A[2]),
    .A2(net23),
    .ZN(\V1/V1/V1/v2 [0]));
 AND2_X1 \V1/V1/V1/V2/_1_  (.A1(A[2]),
    .A2(B[1]),
    .ZN(\V1/V1/V1/V2/w1 ));
 AND2_X1 \V1/V1/V1/V2/_2_  (.A1(net23),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V2/w2 ));
 AND2_X1 \V1/V1/V1/V2/_3_  (.A1(B[1]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V2/w3 ));
 AND2_X1 \V1/V1/V1/V3/HA1/_0_  (.A1(\V1/V1/V1/V3/w2 ),
    .A2(\V1/V1/V1/V3/w1 ),
    .ZN(\V1/V1/V1/V3/w4 ));
 XOR2_X2 \V1/V1/V1/V3/HA1/_1_  (.A(\V1/V1/V1/V3/w2 ),
    .B(\V1/V1/V1/V3/w1 ),
    .Z(\V1/V1/V1/v3 [1]));
 AND2_X1 \V1/V1/V1/V3/HA2/_0_  (.A1(\V1/V1/V1/V3/w4 ),
    .A2(\V1/V1/V1/V3/w3 ),
    .ZN(\V1/V1/V1/v3 [3]));
 XOR2_X2 \V1/V1/V1/V3/HA2/_1_  (.A(\V1/V1/V1/V3/w4 ),
    .B(\V1/V1/V1/V3/w3 ),
    .Z(\V1/V1/V1/v3 [2]));
 AND2_X1 \V1/V1/V1/V3/_0_  (.A1(net48),
    .A2(B[2]),
    .ZN(\V1/V1/V1/v3 [0]));
 AND2_X1 \V1/V1/V1/V3/_1_  (.A1(net48),
    .A2(B[3]),
    .ZN(\V1/V1/V1/V3/w1 ));
 AND2_X1 \V1/V1/V1/V3/_2_  (.A1(B[2]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V3/w2 ));
 AND2_X1 \V1/V1/V1/V3/_3_  (.A1(B[3]),
    .A2(A[1]),
    .ZN(\V1/V1/V1/V3/w3 ));
 AND2_X1 \V1/V1/V1/V4/HA1/_0_  (.A1(\V1/V1/V1/V4/w2 ),
    .A2(\V1/V1/V1/V4/w1 ),
    .ZN(\V1/V1/V1/V4/w4 ));
 XOR2_X2 \V1/V1/V1/V4/HA1/_1_  (.A(\V1/V1/V1/V4/w2 ),
    .B(\V1/V1/V1/V4/w1 ),
    .Z(\V1/V1/V1/v4 [1]));
 AND2_X1 \V1/V1/V1/V4/HA2/_0_  (.A1(\V1/V1/V1/V4/w4 ),
    .A2(\V1/V1/V1/V4/w3 ),
    .ZN(\V1/V1/V1/v4 [3]));
 XOR2_X2 \V1/V1/V1/V4/HA2/_1_  (.A(\V1/V1/V1/V4/w4 ),
    .B(\V1/V1/V1/V4/w3 ),
    .Z(\V1/V1/V1/v4 [2]));
 AND2_X1 \V1/V1/V1/V4/_0_  (.A1(A[2]),
    .A2(B[2]),
    .ZN(\V1/V1/V1/v4 [0]));
 AND2_X1 \V1/V1/V1/V4/_1_  (.A1(A[2]),
    .A2(B[3]),
    .ZN(\V1/V1/V1/V4/w1 ));
 AND2_X1 \V1/V1/V1/V4/_2_  (.A1(B[2]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V4/w2 ));
 AND2_X1 \V1/V1/V1/V4/_3_  (.A1(B[3]),
    .A2(A[3]),
    .ZN(\V1/V1/V1/V4/w3 ));
 OR2_X1 \V1/V1/V1/_0_  (.A1(\V1/V1/V1/c1 ),
    .A2(\V1/V1/V1/c2 ),
    .ZN(\V1/V1/V1/c3 ));
 AND2_X1 \V1/V1/V2/A1/M1/M1/_0_  (.A1(\V1/V1/V2/v2 [0]),
    .A2(\V1/V1/V2/v3 [0]),
    .ZN(\V1/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M1/M1/_1_  (.A(\V1/V1/V2/v2 [0]),
    .B(\V1/V1/V2/v3 [0]),
    .Z(\V1/V1/V2/A1/M1/s1 ));
 AND2_X1 \V1/V1/V2/A1/M1/M2/_0_  (.A1(\V1/V1/V2/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M1/M2/_1_  (.A(\V1/V1/V2/A1/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/V2/s1 [0]));
 OR2_X1 \V1/V1/V2/A1/M1/_0_  (.A1(\V1/V1/V2/A1/M1/c1 ),
    .A2(\V1/V1/V2/A1/M1/c2 ),
    .ZN(\V1/V1/V2/A1/c1 ));
 AND2_X1 \V1/V1/V2/A1/M2/M1/_0_  (.A1(\V1/V1/V2/v2 [1]),
    .A2(\V1/V1/V2/v3 [1]),
    .ZN(\V1/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M2/M1/_1_  (.A(\V1/V1/V2/v2 [1]),
    .B(\V1/V1/V2/v3 [1]),
    .Z(\V1/V1/V2/A1/M2/s1 ));
 AND2_X1 \V1/V1/V2/A1/M2/M2/_0_  (.A1(\V1/V1/V2/A1/M2/s1 ),
    .A2(\V1/V1/V2/A1/c1 ),
    .ZN(\V1/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M2/M2/_1_  (.A(\V1/V1/V2/A1/M2/s1 ),
    .B(\V1/V1/V2/A1/c1 ),
    .Z(\V1/V1/V2/s1 [1]));
 OR2_X1 \V1/V1/V2/A1/M2/_0_  (.A1(\V1/V1/V2/A1/M2/c1 ),
    .A2(\V1/V1/V2/A1/M2/c2 ),
    .ZN(\V1/V1/V2/A1/c2 ));
 AND2_X1 \V1/V1/V2/A1/M3/M1/_0_  (.A1(\V1/V1/V2/v2 [2]),
    .A2(\V1/V1/V2/v3 [2]),
    .ZN(\V1/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M3/M1/_1_  (.A(\V1/V1/V2/v2 [2]),
    .B(\V1/V1/V2/v3 [2]),
    .Z(\V1/V1/V2/A1/M3/s1 ));
 AND2_X1 \V1/V1/V2/A1/M3/M2/_0_  (.A1(\V1/V1/V2/A1/M3/s1 ),
    .A2(\V1/V1/V2/A1/c2 ),
    .ZN(\V1/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M3/M2/_1_  (.A(\V1/V1/V2/A1/M3/s1 ),
    .B(\V1/V1/V2/A1/c2 ),
    .Z(\V1/V1/V2/s1 [2]));
 OR2_X1 \V1/V1/V2/A1/M3/_0_  (.A1(\V1/V1/V2/A1/M3/c1 ),
    .A2(\V1/V1/V2/A1/M3/c2 ),
    .ZN(\V1/V1/V2/A1/c3 ));
 AND2_X1 \V1/V1/V2/A1/M4/M1/_0_  (.A1(\V1/V1/V2/v2 [3]),
    .A2(\V1/V1/V2/v3 [3]),
    .ZN(\V1/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A1/M4/M1/_1_  (.A(\V1/V1/V2/v2 [3]),
    .B(\V1/V1/V2/v3 [3]),
    .Z(\V1/V1/V2/A1/M4/s1 ));
 AND2_X1 \V1/V1/V2/A1/M4/M2/_0_  (.A1(\V1/V1/V2/A1/M4/s1 ),
    .A2(\V1/V1/V2/A1/c3 ),
    .ZN(\V1/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A1/M4/M2/_1_  (.A(\V1/V1/V2/A1/M4/s1 ),
    .B(\V1/V1/V2/A1/c3 ),
    .Z(\V1/V1/V2/s1 [3]));
 OR2_X1 \V1/V1/V2/A1/M4/_0_  (.A1(\V1/V1/V2/A1/M4/c1 ),
    .A2(\V1/V1/V2/A1/M4/c2 ),
    .ZN(\V1/V1/V2/c1 ));
 AND2_X1 \V1/V1/V2/A2/M1/M1/_0_  (.A1(\V1/V1/V2/s1 [0]),
    .A2(\V1/V1/V2/v1 [2]),
    .ZN(\V1/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M1/M1/_1_  (.A(\V1/V1/V2/s1 [0]),
    .B(\V1/V1/V2/v1 [2]),
    .Z(\V1/V1/V2/A2/M1/s1 ));
 AND2_X1 \V1/V1/V2/A2/M1/M2/_0_  (.A1(\V1/V1/V2/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M1/M2/_1_  (.A(\V1/V1/V2/A2/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/v2 [2]));
 OR2_X1 \V1/V1/V2/A2/M1/_0_  (.A1(\V1/V1/V2/A2/M1/c1 ),
    .A2(\V1/V1/V2/A2/M1/c2 ),
    .ZN(\V1/V1/V2/A2/c1 ));
 AND2_X1 \V1/V1/V2/A2/M2/M1/_0_  (.A1(\V1/V1/V2/s1 [1]),
    .A2(\V1/V1/V2/v1 [3]),
    .ZN(\V1/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M2/M1/_1_  (.A(\V1/V1/V2/s1 [1]),
    .B(\V1/V1/V2/v1 [3]),
    .Z(\V1/V1/V2/A2/M2/s1 ));
 AND2_X1 \V1/V1/V2/A2/M2/M2/_0_  (.A1(\V1/V1/V2/A2/M2/s1 ),
    .A2(\V1/V1/V2/A2/c1 ),
    .ZN(\V1/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M2/M2/_1_  (.A(\V1/V1/V2/A2/M2/s1 ),
    .B(\V1/V1/V2/A2/c1 ),
    .Z(\V1/V1/v2 [3]));
 OR2_X1 \V1/V1/V2/A2/M2/_0_  (.A1(\V1/V1/V2/A2/M2/c1 ),
    .A2(\V1/V1/V2/A2/M2/c2 ),
    .ZN(\V1/V1/V2/A2/c2 ));
 AND2_X1 \V1/V1/V2/A2/M3/M1/_0_  (.A1(\V1/V1/V2/s1 [2]),
    .A2(net2),
    .ZN(\V1/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M3/M1/_1_  (.A(\V1/V1/V2/s1 [2]),
    .B(net2),
    .Z(\V1/V1/V2/A2/M3/s1 ));
 AND2_X1 \V1/V1/V2/A2/M3/M2/_0_  (.A1(\V1/V1/V2/A2/M3/s1 ),
    .A2(\V1/V1/V2/A2/c2 ),
    .ZN(\V1/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M3/M2/_1_  (.A(\V1/V1/V2/A2/M3/s1 ),
    .B(\V1/V1/V2/A2/c2 ),
    .Z(\V1/V1/V2/s2 [2]));
 OR2_X1 \V1/V1/V2/A2/M3/_0_  (.A1(\V1/V1/V2/A2/M3/c1 ),
    .A2(\V1/V1/V2/A2/M3/c2 ),
    .ZN(\V1/V1/V2/A2/c3 ));
 AND2_X1 \V1/V1/V2/A2/M4/M1/_0_  (.A1(\V1/V1/V2/s1 [3]),
    .A2(net2),
    .ZN(\V1/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A2/M4/M1/_1_  (.A(\V1/V1/V2/s1 [3]),
    .B(net2),
    .Z(\V1/V1/V2/A2/M4/s1 ));
 AND2_X1 \V1/V1/V2/A2/M4/M2/_0_  (.A1(\V1/V1/V2/A2/M4/s1 ),
    .A2(\V1/V1/V2/A2/c3 ),
    .ZN(\V1/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A2/M4/M2/_1_  (.A(\V1/V1/V2/A2/M4/s1 ),
    .B(\V1/V1/V2/A2/c3 ),
    .Z(\V1/V1/V2/s2 [3]));
 OR2_X1 \V1/V1/V2/A2/M4/_0_  (.A1(\V1/V1/V2/A2/M4/c1 ),
    .A2(\V1/V1/V2/A2/M4/c2 ),
    .ZN(\V1/V1/V2/c2 ));
 AND2_X1 \V1/V1/V2/A3/M1/M1/_0_  (.A1(\V1/V1/V2/v4 [0]),
    .A2(\V1/V1/V2/s2 [2]),
    .ZN(\V1/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M1/M1/_1_  (.A(\V1/V1/V2/v4 [0]),
    .B(\V1/V1/V2/s2 [2]),
    .Z(\V1/V1/V2/A3/M1/s1 ));
 AND2_X1 \V1/V1/V2/A3/M1/M2/_0_  (.A1(\V1/V1/V2/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M1/M2/_1_  (.A(\V1/V1/V2/A3/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/v2 [4]));
 OR2_X1 \V1/V1/V2/A3/M1/_0_  (.A1(\V1/V1/V2/A3/M1/c1 ),
    .A2(\V1/V1/V2/A3/M1/c2 ),
    .ZN(\V1/V1/V2/A3/c1 ));
 AND2_X1 \V1/V1/V2/A3/M2/M1/_0_  (.A1(\V1/V1/V2/v4 [1]),
    .A2(\V1/V1/V2/s2 [3]),
    .ZN(\V1/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M2/M1/_1_  (.A(\V1/V1/V2/v4 [1]),
    .B(\V1/V1/V2/s2 [3]),
    .Z(\V1/V1/V2/A3/M2/s1 ));
 AND2_X1 \V1/V1/V2/A3/M2/M2/_0_  (.A1(\V1/V1/V2/A3/M2/s1 ),
    .A2(\V1/V1/V2/A3/c1 ),
    .ZN(\V1/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M2/M2/_1_  (.A(\V1/V1/V2/A3/M2/s1 ),
    .B(\V1/V1/V2/A3/c1 ),
    .Z(\V1/V1/v2 [5]));
 OR2_X1 \V1/V1/V2/A3/M2/_0_  (.A1(\V1/V1/V2/A3/M2/c1 ),
    .A2(\V1/V1/V2/A3/M2/c2 ),
    .ZN(\V1/V1/V2/A3/c2 ));
 AND2_X1 \V1/V1/V2/A3/M3/M1/_0_  (.A1(\V1/V1/V2/v4 [2]),
    .A2(\V1/V1/V2/c3 ),
    .ZN(\V1/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M3/M1/_1_  (.A(\V1/V1/V2/v4 [2]),
    .B(\V1/V1/V2/c3 ),
    .Z(\V1/V1/V2/A3/M3/s1 ));
 AND2_X1 \V1/V1/V2/A3/M3/M2/_0_  (.A1(\V1/V1/V2/A3/M3/s1 ),
    .A2(\V1/V1/V2/A3/c2 ),
    .ZN(\V1/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M3/M2/_1_  (.A(\V1/V1/V2/A3/M3/s1 ),
    .B(\V1/V1/V2/A3/c2 ),
    .Z(\V1/V1/v2 [6]));
 OR2_X1 \V1/V1/V2/A3/M3/_0_  (.A1(\V1/V1/V2/A3/M3/c1 ),
    .A2(\V1/V1/V2/A3/M3/c2 ),
    .ZN(\V1/V1/V2/A3/c3 ));
 AND2_X1 \V1/V1/V2/A3/M4/M1/_0_  (.A1(\V1/V1/V2/v4 [3]),
    .A2(net2),
    .ZN(\V1/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V2/A3/M4/M1/_1_  (.A(\V1/V1/V2/v4 [3]),
    .B(net2),
    .Z(\V1/V1/V2/A3/M4/s1 ));
 AND2_X1 \V1/V1/V2/A3/M4/M2/_0_  (.A1(\V1/V1/V2/A3/M4/s1 ),
    .A2(\V1/V1/V2/A3/c3 ),
    .ZN(\V1/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V2/A3/M4/M2/_1_  (.A(\V1/V1/V2/A3/M4/s1 ),
    .B(\V1/V1/V2/A3/c3 ),
    .Z(\V1/V1/v2 [7]));
 OR2_X1 \V1/V1/V2/A3/M4/_0_  (.A1(\V1/V1/V2/A3/M4/c1 ),
    .A2(\V1/V1/V2/A3/M4/c2 ),
    .ZN(\V1/V1/V2/overflow ));
 AND2_X1 \V1/V1/V2/V1/HA1/_0_  (.A1(\V1/V1/V2/V1/w2 ),
    .A2(\V1/V1/V2/V1/w1 ),
    .ZN(\V1/V1/V2/V1/w4 ));
 XOR2_X2 \V1/V1/V2/V1/HA1/_1_  (.A(\V1/V1/V2/V1/w2 ),
    .B(\V1/V1/V2/V1/w1 ),
    .Z(\V1/V1/v2 [1]));
 AND2_X1 \V1/V1/V2/V1/HA2/_0_  (.A1(\V1/V1/V2/V1/w4 ),
    .A2(\V1/V1/V2/V1/w3 ),
    .ZN(\V1/V1/V2/v1 [3]));
 XOR2_X2 \V1/V1/V2/V1/HA2/_1_  (.A(\V1/V1/V2/V1/w4 ),
    .B(\V1/V1/V2/V1/w3 ),
    .Z(\V1/V1/V2/v1 [2]));
 AND2_X1 \V1/V1/V2/V1/_0_  (.A1(A[4]),
    .A2(B[0]),
    .ZN(\V1/V1/v2 [0]));
 AND2_X1 \V1/V1/V2/V1/_1_  (.A1(A[4]),
    .A2(B[1]),
    .ZN(\V1/V1/V2/V1/w1 ));
 AND2_X1 \V1/V1/V2/V1/_2_  (.A1(B[0]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V1/w2 ));
 AND2_X1 \V1/V1/V2/V1/_3_  (.A1(B[1]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V1/w3 ));
 AND2_X1 \V1/V1/V2/V2/HA1/_0_  (.A1(\V1/V1/V2/V2/w2 ),
    .A2(\V1/V1/V2/V2/w1 ),
    .ZN(\V1/V1/V2/V2/w4 ));
 XOR2_X2 \V1/V1/V2/V2/HA1/_1_  (.A(\V1/V1/V2/V2/w2 ),
    .B(\V1/V1/V2/V2/w1 ),
    .Z(\V1/V1/V2/v2 [1]));
 AND2_X1 \V1/V1/V2/V2/HA2/_0_  (.A1(\V1/V1/V2/V2/w4 ),
    .A2(\V1/V1/V2/V2/w3 ),
    .ZN(\V1/V1/V2/v2 [3]));
 XOR2_X2 \V1/V1/V2/V2/HA2/_1_  (.A(\V1/V1/V2/V2/w4 ),
    .B(\V1/V1/V2/V2/w3 ),
    .Z(\V1/V1/V2/v2 [2]));
 AND2_X1 \V1/V1/V2/V2/_0_  (.A1(A[6]),
    .A2(B[0]),
    .ZN(\V1/V1/V2/v2 [0]));
 AND2_X1 \V1/V1/V2/V2/_1_  (.A1(A[6]),
    .A2(B[1]),
    .ZN(\V1/V1/V2/V2/w1 ));
 AND2_X1 \V1/V1/V2/V2/_2_  (.A1(B[0]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V2/w2 ));
 AND2_X1 \V1/V1/V2/V2/_3_  (.A1(B[1]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V2/w3 ));
 AND2_X1 \V1/V1/V2/V3/HA1/_0_  (.A1(\V1/V1/V2/V3/w2 ),
    .A2(\V1/V1/V2/V3/w1 ),
    .ZN(\V1/V1/V2/V3/w4 ));
 XOR2_X2 \V1/V1/V2/V3/HA1/_1_  (.A(\V1/V1/V2/V3/w2 ),
    .B(\V1/V1/V2/V3/w1 ),
    .Z(\V1/V1/V2/v3 [1]));
 AND2_X1 \V1/V1/V2/V3/HA2/_0_  (.A1(\V1/V1/V2/V3/w4 ),
    .A2(\V1/V1/V2/V3/w3 ),
    .ZN(\V1/V1/V2/v3 [3]));
 XOR2_X2 \V1/V1/V2/V3/HA2/_1_  (.A(\V1/V1/V2/V3/w4 ),
    .B(\V1/V1/V2/V3/w3 ),
    .Z(\V1/V1/V2/v3 [2]));
 AND2_X1 \V1/V1/V2/V3/_0_  (.A1(A[4]),
    .A2(B[2]),
    .ZN(\V1/V1/V2/v3 [0]));
 AND2_X1 \V1/V1/V2/V3/_1_  (.A1(A[4]),
    .A2(B[3]),
    .ZN(\V1/V1/V2/V3/w1 ));
 AND2_X1 \V1/V1/V2/V3/_2_  (.A1(B[2]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V3/w2 ));
 AND2_X1 \V1/V1/V2/V3/_3_  (.A1(B[3]),
    .A2(A[5]),
    .ZN(\V1/V1/V2/V3/w3 ));
 AND2_X1 \V1/V1/V2/V4/HA1/_0_  (.A1(\V1/V1/V2/V4/w2 ),
    .A2(\V1/V1/V2/V4/w1 ),
    .ZN(\V1/V1/V2/V4/w4 ));
 XOR2_X2 \V1/V1/V2/V4/HA1/_1_  (.A(\V1/V1/V2/V4/w2 ),
    .B(\V1/V1/V2/V4/w1 ),
    .Z(\V1/V1/V2/v4 [1]));
 AND2_X1 \V1/V1/V2/V4/HA2/_0_  (.A1(\V1/V1/V2/V4/w4 ),
    .A2(\V1/V1/V2/V4/w3 ),
    .ZN(\V1/V1/V2/v4 [3]));
 XOR2_X2 \V1/V1/V2/V4/HA2/_1_  (.A(\V1/V1/V2/V4/w4 ),
    .B(\V1/V1/V2/V4/w3 ),
    .Z(\V1/V1/V2/v4 [2]));
 AND2_X1 \V1/V1/V2/V4/_0_  (.A1(A[6]),
    .A2(B[2]),
    .ZN(\V1/V1/V2/v4 [0]));
 AND2_X1 \V1/V1/V2/V4/_1_  (.A1(A[6]),
    .A2(B[3]),
    .ZN(\V1/V1/V2/V4/w1 ));
 AND2_X1 \V1/V1/V2/V4/_2_  (.A1(B[2]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V4/w2 ));
 AND2_X1 \V1/V1/V2/V4/_3_  (.A1(B[3]),
    .A2(A[7]),
    .ZN(\V1/V1/V2/V4/w3 ));
 OR2_X1 \V1/V1/V2/_0_  (.A1(\V1/V1/V2/c1 ),
    .A2(\V1/V1/V2/c2 ),
    .ZN(\V1/V1/V2/c3 ));
 AND2_X1 \V1/V1/V3/A1/M1/M1/_0_  (.A1(\V1/V1/V3/v2 [0]),
    .A2(\V1/V1/V3/v3 [0]),
    .ZN(\V1/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M1/M1/_1_  (.A(\V1/V1/V3/v2 [0]),
    .B(\V1/V1/V3/v3 [0]),
    .Z(\V1/V1/V3/A1/M1/s1 ));
 AND2_X1 \V1/V1/V3/A1/M1/M2/_0_  (.A1(\V1/V1/V3/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M1/M2/_1_  (.A(\V1/V1/V3/A1/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/V3/s1 [0]));
 OR2_X1 \V1/V1/V3/A1/M1/_0_  (.A1(\V1/V1/V3/A1/M1/c1 ),
    .A2(\V1/V1/V3/A1/M1/c2 ),
    .ZN(\V1/V1/V3/A1/c1 ));
 AND2_X1 \V1/V1/V3/A1/M2/M1/_0_  (.A1(\V1/V1/V3/v2 [1]),
    .A2(\V1/V1/V3/v3 [1]),
    .ZN(\V1/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M2/M1/_1_  (.A(\V1/V1/V3/v2 [1]),
    .B(\V1/V1/V3/v3 [1]),
    .Z(\V1/V1/V3/A1/M2/s1 ));
 AND2_X1 \V1/V1/V3/A1/M2/M2/_0_  (.A1(\V1/V1/V3/A1/M2/s1 ),
    .A2(\V1/V1/V3/A1/c1 ),
    .ZN(\V1/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M2/M2/_1_  (.A(\V1/V1/V3/A1/M2/s1 ),
    .B(\V1/V1/V3/A1/c1 ),
    .Z(\V1/V1/V3/s1 [1]));
 OR2_X1 \V1/V1/V3/A1/M2/_0_  (.A1(\V1/V1/V3/A1/M2/c1 ),
    .A2(\V1/V1/V3/A1/M2/c2 ),
    .ZN(\V1/V1/V3/A1/c2 ));
 AND2_X1 \V1/V1/V3/A1/M3/M1/_0_  (.A1(\V1/V1/V3/v2 [2]),
    .A2(\V1/V1/V3/v3 [2]),
    .ZN(\V1/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M3/M1/_1_  (.A(\V1/V1/V3/v2 [2]),
    .B(\V1/V1/V3/v3 [2]),
    .Z(\V1/V1/V3/A1/M3/s1 ));
 AND2_X1 \V1/V1/V3/A1/M3/M2/_0_  (.A1(\V1/V1/V3/A1/M3/s1 ),
    .A2(\V1/V1/V3/A1/c2 ),
    .ZN(\V1/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M3/M2/_1_  (.A(\V1/V1/V3/A1/M3/s1 ),
    .B(\V1/V1/V3/A1/c2 ),
    .Z(\V1/V1/V3/s1 [2]));
 OR2_X1 \V1/V1/V3/A1/M3/_0_  (.A1(\V1/V1/V3/A1/M3/c1 ),
    .A2(\V1/V1/V3/A1/M3/c2 ),
    .ZN(\V1/V1/V3/A1/c3 ));
 AND2_X1 \V1/V1/V3/A1/M4/M1/_0_  (.A1(\V1/V1/V3/v2 [3]),
    .A2(\V1/V1/V3/v3 [3]),
    .ZN(\V1/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A1/M4/M1/_1_  (.A(\V1/V1/V3/v2 [3]),
    .B(\V1/V1/V3/v3 [3]),
    .Z(\V1/V1/V3/A1/M4/s1 ));
 AND2_X1 \V1/V1/V3/A1/M4/M2/_0_  (.A1(\V1/V1/V3/A1/M4/s1 ),
    .A2(\V1/V1/V3/A1/c3 ),
    .ZN(\V1/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A1/M4/M2/_1_  (.A(\V1/V1/V3/A1/M4/s1 ),
    .B(\V1/V1/V3/A1/c3 ),
    .Z(\V1/V1/V3/s1 [3]));
 OR2_X1 \V1/V1/V3/A1/M4/_0_  (.A1(\V1/V1/V3/A1/M4/c1 ),
    .A2(\V1/V1/V3/A1/M4/c2 ),
    .ZN(\V1/V1/V3/c1 ));
 AND2_X1 \V1/V1/V3/A2/M1/M1/_0_  (.A1(\V1/V1/V3/s1 [0]),
    .A2(\V1/V1/V3/v1 [2]),
    .ZN(\V1/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M1/M1/_1_  (.A(\V1/V1/V3/s1 [0]),
    .B(\V1/V1/V3/v1 [2]),
    .Z(\V1/V1/V3/A2/M1/s1 ));
 AND2_X1 \V1/V1/V3/A2/M1/M2/_0_  (.A1(\V1/V1/V3/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M1/M2/_1_  (.A(\V1/V1/V3/A2/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/v3 [2]));
 OR2_X1 \V1/V1/V3/A2/M1/_0_  (.A1(\V1/V1/V3/A2/M1/c1 ),
    .A2(\V1/V1/V3/A2/M1/c2 ),
    .ZN(\V1/V1/V3/A2/c1 ));
 AND2_X1 \V1/V1/V3/A2/M2/M1/_0_  (.A1(\V1/V1/V3/s1 [1]),
    .A2(\V1/V1/V3/v1 [3]),
    .ZN(\V1/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M2/M1/_1_  (.A(\V1/V1/V3/s1 [1]),
    .B(\V1/V1/V3/v1 [3]),
    .Z(\V1/V1/V3/A2/M2/s1 ));
 AND2_X1 \V1/V1/V3/A2/M2/M2/_0_  (.A1(\V1/V1/V3/A2/M2/s1 ),
    .A2(\V1/V1/V3/A2/c1 ),
    .ZN(\V1/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M2/M2/_1_  (.A(\V1/V1/V3/A2/M2/s1 ),
    .B(\V1/V1/V3/A2/c1 ),
    .Z(\V1/V1/v3 [3]));
 OR2_X1 \V1/V1/V3/A2/M2/_0_  (.A1(\V1/V1/V3/A2/M2/c1 ),
    .A2(\V1/V1/V3/A2/M2/c2 ),
    .ZN(\V1/V1/V3/A2/c2 ));
 AND2_X1 \V1/V1/V3/A2/M3/M1/_0_  (.A1(\V1/V1/V3/s1 [2]),
    .A2(net2),
    .ZN(\V1/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M3/M1/_1_  (.A(\V1/V1/V3/s1 [2]),
    .B(net2),
    .Z(\V1/V1/V3/A2/M3/s1 ));
 AND2_X1 \V1/V1/V3/A2/M3/M2/_0_  (.A1(\V1/V1/V3/A2/M3/s1 ),
    .A2(\V1/V1/V3/A2/c2 ),
    .ZN(\V1/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M3/M2/_1_  (.A(\V1/V1/V3/A2/M3/s1 ),
    .B(\V1/V1/V3/A2/c2 ),
    .Z(\V1/V1/V3/s2 [2]));
 OR2_X1 \V1/V1/V3/A2/M3/_0_  (.A1(\V1/V1/V3/A2/M3/c1 ),
    .A2(\V1/V1/V3/A2/M3/c2 ),
    .ZN(\V1/V1/V3/A2/c3 ));
 AND2_X1 \V1/V1/V3/A2/M4/M1/_0_  (.A1(\V1/V1/V3/s1 [3]),
    .A2(net2),
    .ZN(\V1/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A2/M4/M1/_1_  (.A(\V1/V1/V3/s1 [3]),
    .B(net2),
    .Z(\V1/V1/V3/A2/M4/s1 ));
 AND2_X1 \V1/V1/V3/A2/M4/M2/_0_  (.A1(\V1/V1/V3/A2/M4/s1 ),
    .A2(\V1/V1/V3/A2/c3 ),
    .ZN(\V1/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A2/M4/M2/_1_  (.A(\V1/V1/V3/A2/M4/s1 ),
    .B(\V1/V1/V3/A2/c3 ),
    .Z(\V1/V1/V3/s2 [3]));
 OR2_X1 \V1/V1/V3/A2/M4/_0_  (.A1(\V1/V1/V3/A2/M4/c1 ),
    .A2(\V1/V1/V3/A2/M4/c2 ),
    .ZN(\V1/V1/V3/c2 ));
 AND2_X1 \V1/V1/V3/A3/M1/M1/_0_  (.A1(\V1/V1/V3/v4 [0]),
    .A2(\V1/V1/V3/s2 [2]),
    .ZN(\V1/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M1/M1/_1_  (.A(\V1/V1/V3/v4 [0]),
    .B(\V1/V1/V3/s2 [2]),
    .Z(\V1/V1/V3/A3/M1/s1 ));
 AND2_X1 \V1/V1/V3/A3/M1/M2/_0_  (.A1(\V1/V1/V3/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V1/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M1/M2/_1_  (.A(\V1/V1/V3/A3/M1/s1 ),
    .B(net2),
    .Z(\V1/V1/v3 [4]));
 OR2_X1 \V1/V1/V3/A3/M1/_0_  (.A1(\V1/V1/V3/A3/M1/c1 ),
    .A2(\V1/V1/V3/A3/M1/c2 ),
    .ZN(\V1/V1/V3/A3/c1 ));
 AND2_X1 \V1/V1/V3/A3/M2/M1/_0_  (.A1(\V1/V1/V3/v4 [1]),
    .A2(\V1/V1/V3/s2 [3]),
    .ZN(\V1/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M2/M1/_1_  (.A(\V1/V1/V3/v4 [1]),
    .B(\V1/V1/V3/s2 [3]),
    .Z(\V1/V1/V3/A3/M2/s1 ));
 AND2_X1 \V1/V1/V3/A3/M2/M2/_0_  (.A1(\V1/V1/V3/A3/M2/s1 ),
    .A2(\V1/V1/V3/A3/c1 ),
    .ZN(\V1/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M2/M2/_1_  (.A(\V1/V1/V3/A3/M2/s1 ),
    .B(\V1/V1/V3/A3/c1 ),
    .Z(\V1/V1/v3 [5]));
 OR2_X1 \V1/V1/V3/A3/M2/_0_  (.A1(\V1/V1/V3/A3/M2/c1 ),
    .A2(\V1/V1/V3/A3/M2/c2 ),
    .ZN(\V1/V1/V3/A3/c2 ));
 AND2_X1 \V1/V1/V3/A3/M3/M1/_0_  (.A1(\V1/V1/V3/v4 [2]),
    .A2(\V1/V1/V3/c3 ),
    .ZN(\V1/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M3/M1/_1_  (.A(\V1/V1/V3/v4 [2]),
    .B(\V1/V1/V3/c3 ),
    .Z(\V1/V1/V3/A3/M3/s1 ));
 AND2_X1 \V1/V1/V3/A3/M3/M2/_0_  (.A1(\V1/V1/V3/A3/M3/s1 ),
    .A2(\V1/V1/V3/A3/c2 ),
    .ZN(\V1/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M3/M2/_1_  (.A(\V1/V1/V3/A3/M3/s1 ),
    .B(\V1/V1/V3/A3/c2 ),
    .Z(\V1/V1/v3 [6]));
 OR2_X1 \V1/V1/V3/A3/M3/_0_  (.A1(\V1/V1/V3/A3/M3/c1 ),
    .A2(\V1/V1/V3/A3/M3/c2 ),
    .ZN(\V1/V1/V3/A3/c3 ));
 AND2_X1 \V1/V1/V3/A3/M4/M1/_0_  (.A1(\V1/V1/V3/v4 [3]),
    .A2(net2),
    .ZN(\V1/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V3/A3/M4/M1/_1_  (.A(\V1/V1/V3/v4 [3]),
    .B(net2),
    .Z(\V1/V1/V3/A3/M4/s1 ));
 AND2_X1 \V1/V1/V3/A3/M4/M2/_0_  (.A1(\V1/V1/V3/A3/M4/s1 ),
    .A2(\V1/V1/V3/A3/c3 ),
    .ZN(\V1/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V3/A3/M4/M2/_1_  (.A(\V1/V1/V3/A3/M4/s1 ),
    .B(\V1/V1/V3/A3/c3 ),
    .Z(\V1/V1/v3 [7]));
 OR2_X1 \V1/V1/V3/A3/M4/_0_  (.A1(\V1/V1/V3/A3/M4/c1 ),
    .A2(\V1/V1/V3/A3/M4/c2 ),
    .ZN(\V1/V1/V3/overflow ));
 AND2_X1 \V1/V1/V3/V1/HA1/_0_  (.A1(\V1/V1/V3/V1/w2 ),
    .A2(\V1/V1/V3/V1/w1 ),
    .ZN(\V1/V1/V3/V1/w4 ));
 XOR2_X2 \V1/V1/V3/V1/HA1/_1_  (.A(\V1/V1/V3/V1/w2 ),
    .B(\V1/V1/V3/V1/w1 ),
    .Z(\V1/V1/v3 [1]));
 AND2_X1 \V1/V1/V3/V1/HA2/_0_  (.A1(\V1/V1/V3/V1/w4 ),
    .A2(\V1/V1/V3/V1/w3 ),
    .ZN(\V1/V1/V3/v1 [3]));
 XOR2_X2 \V1/V1/V3/V1/HA2/_1_  (.A(\V1/V1/V3/V1/w4 ),
    .B(\V1/V1/V3/V1/w3 ),
    .Z(\V1/V1/V3/v1 [2]));
 AND2_X1 \V1/V1/V3/V1/_0_  (.A1(net48),
    .A2(B[4]),
    .ZN(\V1/V1/v3 [0]));
 AND2_X1 \V1/V1/V3/V1/_1_  (.A1(net48),
    .A2(B[5]),
    .ZN(\V1/V1/V3/V1/w1 ));
 AND2_X1 \V1/V1/V3/V1/_2_  (.A1(B[4]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V1/w2 ));
 AND2_X1 \V1/V1/V3/V1/_3_  (.A1(B[5]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V1/w3 ));
 AND2_X1 \V1/V1/V3/V2/HA1/_0_  (.A1(\V1/V1/V3/V2/w2 ),
    .A2(\V1/V1/V3/V2/w1 ),
    .ZN(\V1/V1/V3/V2/w4 ));
 XOR2_X2 \V1/V1/V3/V2/HA1/_1_  (.A(\V1/V1/V3/V2/w2 ),
    .B(\V1/V1/V3/V2/w1 ),
    .Z(\V1/V1/V3/v2 [1]));
 AND2_X1 \V1/V1/V3/V2/HA2/_0_  (.A1(\V1/V1/V3/V2/w4 ),
    .A2(\V1/V1/V3/V2/w3 ),
    .ZN(\V1/V1/V3/v2 [3]));
 XOR2_X2 \V1/V1/V3/V2/HA2/_1_  (.A(\V1/V1/V3/V2/w4 ),
    .B(\V1/V1/V3/V2/w3 ),
    .Z(\V1/V1/V3/v2 [2]));
 AND2_X1 \V1/V1/V3/V2/_0_  (.A1(A[2]),
    .A2(B[4]),
    .ZN(\V1/V1/V3/v2 [0]));
 AND2_X1 \V1/V1/V3/V2/_1_  (.A1(A[2]),
    .A2(B[5]),
    .ZN(\V1/V1/V3/V2/w1 ));
 AND2_X1 \V1/V1/V3/V2/_2_  (.A1(B[4]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V2/w2 ));
 AND2_X1 \V1/V1/V3/V2/_3_  (.A1(B[5]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V2/w3 ));
 AND2_X1 \V1/V1/V3/V3/HA1/_0_  (.A1(\V1/V1/V3/V3/w2 ),
    .A2(\V1/V1/V3/V3/w1 ),
    .ZN(\V1/V1/V3/V3/w4 ));
 XOR2_X2 \V1/V1/V3/V3/HA1/_1_  (.A(\V1/V1/V3/V3/w2 ),
    .B(\V1/V1/V3/V3/w1 ),
    .Z(\V1/V1/V3/v3 [1]));
 AND2_X1 \V1/V1/V3/V3/HA2/_0_  (.A1(\V1/V1/V3/V3/w4 ),
    .A2(\V1/V1/V3/V3/w3 ),
    .ZN(\V1/V1/V3/v3 [3]));
 XOR2_X2 \V1/V1/V3/V3/HA2/_1_  (.A(\V1/V1/V3/V3/w4 ),
    .B(\V1/V1/V3/V3/w3 ),
    .Z(\V1/V1/V3/v3 [2]));
 AND2_X1 \V1/V1/V3/V3/_0_  (.A1(net48),
    .A2(B[6]),
    .ZN(\V1/V1/V3/v3 [0]));
 AND2_X1 \V1/V1/V3/V3/_1_  (.A1(net48),
    .A2(B[7]),
    .ZN(\V1/V1/V3/V3/w1 ));
 AND2_X1 \V1/V1/V3/V3/_2_  (.A1(B[6]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V3/w2 ));
 AND2_X1 \V1/V1/V3/V3/_3_  (.A1(B[7]),
    .A2(A[1]),
    .ZN(\V1/V1/V3/V3/w3 ));
 AND2_X1 \V1/V1/V3/V4/HA1/_0_  (.A1(\V1/V1/V3/V4/w2 ),
    .A2(\V1/V1/V3/V4/w1 ),
    .ZN(\V1/V1/V3/V4/w4 ));
 XOR2_X2 \V1/V1/V3/V4/HA1/_1_  (.A(\V1/V1/V3/V4/w2 ),
    .B(\V1/V1/V3/V4/w1 ),
    .Z(\V1/V1/V3/v4 [1]));
 AND2_X1 \V1/V1/V3/V4/HA2/_0_  (.A1(\V1/V1/V3/V4/w4 ),
    .A2(\V1/V1/V3/V4/w3 ),
    .ZN(\V1/V1/V3/v4 [3]));
 XOR2_X2 \V1/V1/V3/V4/HA2/_1_  (.A(\V1/V1/V3/V4/w4 ),
    .B(\V1/V1/V3/V4/w3 ),
    .Z(\V1/V1/V3/v4 [2]));
 AND2_X1 \V1/V1/V3/V4/_0_  (.A1(A[2]),
    .A2(B[6]),
    .ZN(\V1/V1/V3/v4 [0]));
 AND2_X1 \V1/V1/V3/V4/_1_  (.A1(A[2]),
    .A2(B[7]),
    .ZN(\V1/V1/V3/V4/w1 ));
 AND2_X1 \V1/V1/V3/V4/_2_  (.A1(B[6]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V4/w2 ));
 AND2_X1 \V1/V1/V3/V4/_3_  (.A1(B[7]),
    .A2(A[3]),
    .ZN(\V1/V1/V3/V4/w3 ));
 OR2_X1 \V1/V1/V3/_0_  (.A1(\V1/V1/V3/c1 ),
    .A2(\V1/V1/V3/c2 ),
    .ZN(\V1/V1/V3/c3 ));
 AND2_X1 \V1/V1/V4/A1/M1/M1/_0_  (.A1(\V1/V1/V4/v2 [0]),
    .A2(\V1/V1/V4/v3 [0]),
    .ZN(\V1/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M1/M1/_1_  (.A(\V1/V1/V4/v2 [0]),
    .B(\V1/V1/V4/v3 [0]),
    .Z(\V1/V1/V4/A1/M1/s1 ));
 AND2_X1 \V1/V1/V4/A1/M1/M2/_0_  (.A1(\V1/V1/V4/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M1/M2/_1_  (.A(\V1/V1/V4/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/V4/s1 [0]));
 OR2_X1 \V1/V1/V4/A1/M1/_0_  (.A1(\V1/V1/V4/A1/M1/c1 ),
    .A2(\V1/V1/V4/A1/M1/c2 ),
    .ZN(\V1/V1/V4/A1/c1 ));
 AND2_X1 \V1/V1/V4/A1/M2/M1/_0_  (.A1(\V1/V1/V4/v2 [1]),
    .A2(\V1/V1/V4/v3 [1]),
    .ZN(\V1/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M2/M1/_1_  (.A(\V1/V1/V4/v2 [1]),
    .B(\V1/V1/V4/v3 [1]),
    .Z(\V1/V1/V4/A1/M2/s1 ));
 AND2_X1 \V1/V1/V4/A1/M2/M2/_0_  (.A1(\V1/V1/V4/A1/M2/s1 ),
    .A2(\V1/V1/V4/A1/c1 ),
    .ZN(\V1/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M2/M2/_1_  (.A(\V1/V1/V4/A1/M2/s1 ),
    .B(\V1/V1/V4/A1/c1 ),
    .Z(\V1/V1/V4/s1 [1]));
 OR2_X1 \V1/V1/V4/A1/M2/_0_  (.A1(\V1/V1/V4/A1/M2/c1 ),
    .A2(\V1/V1/V4/A1/M2/c2 ),
    .ZN(\V1/V1/V4/A1/c2 ));
 AND2_X1 \V1/V1/V4/A1/M3/M1/_0_  (.A1(\V1/V1/V4/v2 [2]),
    .A2(\V1/V1/V4/v3 [2]),
    .ZN(\V1/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M3/M1/_1_  (.A(\V1/V1/V4/v2 [2]),
    .B(\V1/V1/V4/v3 [2]),
    .Z(\V1/V1/V4/A1/M3/s1 ));
 AND2_X1 \V1/V1/V4/A1/M3/M2/_0_  (.A1(\V1/V1/V4/A1/M3/s1 ),
    .A2(\V1/V1/V4/A1/c2 ),
    .ZN(\V1/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M3/M2/_1_  (.A(\V1/V1/V4/A1/M3/s1 ),
    .B(\V1/V1/V4/A1/c2 ),
    .Z(\V1/V1/V4/s1 [2]));
 OR2_X1 \V1/V1/V4/A1/M3/_0_  (.A1(\V1/V1/V4/A1/M3/c1 ),
    .A2(\V1/V1/V4/A1/M3/c2 ),
    .ZN(\V1/V1/V4/A1/c3 ));
 AND2_X1 \V1/V1/V4/A1/M4/M1/_0_  (.A1(\V1/V1/V4/v2 [3]),
    .A2(\V1/V1/V4/v3 [3]),
    .ZN(\V1/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A1/M4/M1/_1_  (.A(\V1/V1/V4/v2 [3]),
    .B(\V1/V1/V4/v3 [3]),
    .Z(\V1/V1/V4/A1/M4/s1 ));
 AND2_X1 \V1/V1/V4/A1/M4/M2/_0_  (.A1(\V1/V1/V4/A1/M4/s1 ),
    .A2(\V1/V1/V4/A1/c3 ),
    .ZN(\V1/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A1/M4/M2/_1_  (.A(\V1/V1/V4/A1/M4/s1 ),
    .B(\V1/V1/V4/A1/c3 ),
    .Z(\V1/V1/V4/s1 [3]));
 OR2_X1 \V1/V1/V4/A1/M4/_0_  (.A1(\V1/V1/V4/A1/M4/c1 ),
    .A2(\V1/V1/V4/A1/M4/c2 ),
    .ZN(\V1/V1/V4/c1 ));
 AND2_X1 \V1/V1/V4/A2/M1/M1/_0_  (.A1(\V1/V1/V4/s1 [0]),
    .A2(\V1/V1/V4/v1 [2]),
    .ZN(\V1/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M1/M1/_1_  (.A(\V1/V1/V4/s1 [0]),
    .B(\V1/V1/V4/v1 [2]),
    .Z(\V1/V1/V4/A2/M1/s1 ));
 AND2_X1 \V1/V1/V4/A2/M1/M2/_0_  (.A1(\V1/V1/V4/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M1/M2/_1_  (.A(\V1/V1/V4/A2/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/v4 [2]));
 OR2_X1 \V1/V1/V4/A2/M1/_0_  (.A1(\V1/V1/V4/A2/M1/c1 ),
    .A2(\V1/V1/V4/A2/M1/c2 ),
    .ZN(\V1/V1/V4/A2/c1 ));
 AND2_X1 \V1/V1/V4/A2/M2/M1/_0_  (.A1(\V1/V1/V4/s1 [1]),
    .A2(\V1/V1/V4/v1 [3]),
    .ZN(\V1/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M2/M1/_1_  (.A(\V1/V1/V4/s1 [1]),
    .B(\V1/V1/V4/v1 [3]),
    .Z(\V1/V1/V4/A2/M2/s1 ));
 AND2_X1 \V1/V1/V4/A2/M2/M2/_0_  (.A1(\V1/V1/V4/A2/M2/s1 ),
    .A2(\V1/V1/V4/A2/c1 ),
    .ZN(\V1/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M2/M2/_1_  (.A(\V1/V1/V4/A2/M2/s1 ),
    .B(\V1/V1/V4/A2/c1 ),
    .Z(\V1/V1/v4 [3]));
 OR2_X1 \V1/V1/V4/A2/M2/_0_  (.A1(\V1/V1/V4/A2/M2/c1 ),
    .A2(\V1/V1/V4/A2/M2/c2 ),
    .ZN(\V1/V1/V4/A2/c2 ));
 AND2_X1 \V1/V1/V4/A2/M3/M1/_0_  (.A1(\V1/V1/V4/s1 [2]),
    .A2(net4),
    .ZN(\V1/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M3/M1/_1_  (.A(\V1/V1/V4/s1 [2]),
    .B(net4),
    .Z(\V1/V1/V4/A2/M3/s1 ));
 AND2_X1 \V1/V1/V4/A2/M3/M2/_0_  (.A1(\V1/V1/V4/A2/M3/s1 ),
    .A2(\V1/V1/V4/A2/c2 ),
    .ZN(\V1/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M3/M2/_1_  (.A(\V1/V1/V4/A2/M3/s1 ),
    .B(\V1/V1/V4/A2/c2 ),
    .Z(\V1/V1/V4/s2 [2]));
 OR2_X1 \V1/V1/V4/A2/M3/_0_  (.A1(\V1/V1/V4/A2/M3/c1 ),
    .A2(\V1/V1/V4/A2/M3/c2 ),
    .ZN(\V1/V1/V4/A2/c3 ));
 AND2_X1 \V1/V1/V4/A2/M4/M1/_0_  (.A1(\V1/V1/V4/s1 [3]),
    .A2(net4),
    .ZN(\V1/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A2/M4/M1/_1_  (.A(\V1/V1/V4/s1 [3]),
    .B(net4),
    .Z(\V1/V1/V4/A2/M4/s1 ));
 AND2_X1 \V1/V1/V4/A2/M4/M2/_0_  (.A1(\V1/V1/V4/A2/M4/s1 ),
    .A2(\V1/V1/V4/A2/c3 ),
    .ZN(\V1/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A2/M4/M2/_1_  (.A(\V1/V1/V4/A2/M4/s1 ),
    .B(\V1/V1/V4/A2/c3 ),
    .Z(\V1/V1/V4/s2 [3]));
 OR2_X1 \V1/V1/V4/A2/M4/_0_  (.A1(\V1/V1/V4/A2/M4/c1 ),
    .A2(\V1/V1/V4/A2/M4/c2 ),
    .ZN(\V1/V1/V4/c2 ));
 AND2_X1 \V1/V1/V4/A3/M1/M1/_0_  (.A1(\V1/V1/V4/v4 [0]),
    .A2(\V1/V1/V4/s2 [2]),
    .ZN(\V1/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M1/M1/_1_  (.A(\V1/V1/V4/v4 [0]),
    .B(\V1/V1/V4/s2 [2]),
    .Z(\V1/V1/V4/A3/M1/s1 ));
 AND2_X1 \V1/V1/V4/A3/M1/M2/_0_  (.A1(\V1/V1/V4/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M1/M2/_1_  (.A(\V1/V1/V4/A3/M1/s1 ),
    .B(net4),
    .Z(\V1/V1/v4 [4]));
 OR2_X1 \V1/V1/V4/A3/M1/_0_  (.A1(\V1/V1/V4/A3/M1/c1 ),
    .A2(\V1/V1/V4/A3/M1/c2 ),
    .ZN(\V1/V1/V4/A3/c1 ));
 AND2_X1 \V1/V1/V4/A3/M2/M1/_0_  (.A1(\V1/V1/V4/v4 [1]),
    .A2(\V1/V1/V4/s2 [3]),
    .ZN(\V1/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M2/M1/_1_  (.A(\V1/V1/V4/v4 [1]),
    .B(\V1/V1/V4/s2 [3]),
    .Z(\V1/V1/V4/A3/M2/s1 ));
 AND2_X1 \V1/V1/V4/A3/M2/M2/_0_  (.A1(\V1/V1/V4/A3/M2/s1 ),
    .A2(\V1/V1/V4/A3/c1 ),
    .ZN(\V1/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M2/M2/_1_  (.A(\V1/V1/V4/A3/M2/s1 ),
    .B(\V1/V1/V4/A3/c1 ),
    .Z(\V1/V1/v4 [5]));
 OR2_X1 \V1/V1/V4/A3/M2/_0_  (.A1(\V1/V1/V4/A3/M2/c1 ),
    .A2(\V1/V1/V4/A3/M2/c2 ),
    .ZN(\V1/V1/V4/A3/c2 ));
 AND2_X1 \V1/V1/V4/A3/M3/M1/_0_  (.A1(\V1/V1/V4/v4 [2]),
    .A2(\V1/V1/V4/c3 ),
    .ZN(\V1/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M3/M1/_1_  (.A(\V1/V1/V4/v4 [2]),
    .B(\V1/V1/V4/c3 ),
    .Z(\V1/V1/V4/A3/M3/s1 ));
 AND2_X1 \V1/V1/V4/A3/M3/M2/_0_  (.A1(\V1/V1/V4/A3/M3/s1 ),
    .A2(\V1/V1/V4/A3/c2 ),
    .ZN(\V1/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M3/M2/_1_  (.A(\V1/V1/V4/A3/M3/s1 ),
    .B(\V1/V1/V4/A3/c2 ),
    .Z(\V1/V1/v4 [6]));
 OR2_X1 \V1/V1/V4/A3/M3/_0_  (.A1(\V1/V1/V4/A3/M3/c1 ),
    .A2(\V1/V1/V4/A3/M3/c2 ),
    .ZN(\V1/V1/V4/A3/c3 ));
 AND2_X1 \V1/V1/V4/A3/M4/M1/_0_  (.A1(\V1/V1/V4/v4 [3]),
    .A2(net4),
    .ZN(\V1/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V1/V4/A3/M4/M1/_1_  (.A(\V1/V1/V4/v4 [3]),
    .B(net4),
    .Z(\V1/V1/V4/A3/M4/s1 ));
 AND2_X1 \V1/V1/V4/A3/M4/M2/_0_  (.A1(\V1/V1/V4/A3/M4/s1 ),
    .A2(\V1/V1/V4/A3/c3 ),
    .ZN(\V1/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V1/V4/A3/M4/M2/_1_  (.A(\V1/V1/V4/A3/M4/s1 ),
    .B(\V1/V1/V4/A3/c3 ),
    .Z(\V1/V1/v4 [7]));
 OR2_X1 \V1/V1/V4/A3/M4/_0_  (.A1(\V1/V1/V4/A3/M4/c1 ),
    .A2(\V1/V1/V4/A3/M4/c2 ),
    .ZN(\V1/V1/V4/overflow ));
 AND2_X1 \V1/V1/V4/V1/HA1/_0_  (.A1(\V1/V1/V4/V1/w2 ),
    .A2(\V1/V1/V4/V1/w1 ),
    .ZN(\V1/V1/V4/V1/w4 ));
 XOR2_X2 \V1/V1/V4/V1/HA1/_1_  (.A(\V1/V1/V4/V1/w2 ),
    .B(\V1/V1/V4/V1/w1 ),
    .Z(\V1/V1/v4 [1]));
 AND2_X1 \V1/V1/V4/V1/HA2/_0_  (.A1(\V1/V1/V4/V1/w4 ),
    .A2(\V1/V1/V4/V1/w3 ),
    .ZN(\V1/V1/V4/v1 [3]));
 XOR2_X2 \V1/V1/V4/V1/HA2/_1_  (.A(\V1/V1/V4/V1/w4 ),
    .B(\V1/V1/V4/V1/w3 ),
    .Z(\V1/V1/V4/v1 [2]));
 AND2_X1 \V1/V1/V4/V1/_0_  (.A1(A[4]),
    .A2(B[4]),
    .ZN(\V1/V1/v4 [0]));
 AND2_X1 \V1/V1/V4/V1/_1_  (.A1(A[4]),
    .A2(B[5]),
    .ZN(\V1/V1/V4/V1/w1 ));
 AND2_X1 \V1/V1/V4/V1/_2_  (.A1(B[4]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V1/w2 ));
 AND2_X1 \V1/V1/V4/V1/_3_  (.A1(B[5]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V1/w3 ));
 AND2_X1 \V1/V1/V4/V2/HA1/_0_  (.A1(\V1/V1/V4/V2/w2 ),
    .A2(\V1/V1/V4/V2/w1 ),
    .ZN(\V1/V1/V4/V2/w4 ));
 XOR2_X2 \V1/V1/V4/V2/HA1/_1_  (.A(\V1/V1/V4/V2/w2 ),
    .B(\V1/V1/V4/V2/w1 ),
    .Z(\V1/V1/V4/v2 [1]));
 AND2_X1 \V1/V1/V4/V2/HA2/_0_  (.A1(\V1/V1/V4/V2/w4 ),
    .A2(\V1/V1/V4/V2/w3 ),
    .ZN(\V1/V1/V4/v2 [3]));
 XOR2_X2 \V1/V1/V4/V2/HA2/_1_  (.A(\V1/V1/V4/V2/w4 ),
    .B(\V1/V1/V4/V2/w3 ),
    .Z(\V1/V1/V4/v2 [2]));
 AND2_X1 \V1/V1/V4/V2/_0_  (.A1(A[6]),
    .A2(B[4]),
    .ZN(\V1/V1/V4/v2 [0]));
 AND2_X1 \V1/V1/V4/V2/_1_  (.A1(A[6]),
    .A2(B[5]),
    .ZN(\V1/V1/V4/V2/w1 ));
 AND2_X1 \V1/V1/V4/V2/_2_  (.A1(B[4]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V2/w2 ));
 AND2_X1 \V1/V1/V4/V2/_3_  (.A1(B[5]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V2/w3 ));
 AND2_X1 \V1/V1/V4/V3/HA1/_0_  (.A1(\V1/V1/V4/V3/w2 ),
    .A2(\V1/V1/V4/V3/w1 ),
    .ZN(\V1/V1/V4/V3/w4 ));
 XOR2_X2 \V1/V1/V4/V3/HA1/_1_  (.A(\V1/V1/V4/V3/w2 ),
    .B(\V1/V1/V4/V3/w1 ),
    .Z(\V1/V1/V4/v3 [1]));
 AND2_X1 \V1/V1/V4/V3/HA2/_0_  (.A1(\V1/V1/V4/V3/w4 ),
    .A2(\V1/V1/V4/V3/w3 ),
    .ZN(\V1/V1/V4/v3 [3]));
 XOR2_X2 \V1/V1/V4/V3/HA2/_1_  (.A(\V1/V1/V4/V3/w4 ),
    .B(\V1/V1/V4/V3/w3 ),
    .Z(\V1/V1/V4/v3 [2]));
 AND2_X1 \V1/V1/V4/V3/_0_  (.A1(A[4]),
    .A2(B[6]),
    .ZN(\V1/V1/V4/v3 [0]));
 AND2_X1 \V1/V1/V4/V3/_1_  (.A1(A[4]),
    .A2(B[7]),
    .ZN(\V1/V1/V4/V3/w1 ));
 AND2_X1 \V1/V1/V4/V3/_2_  (.A1(B[6]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V3/w2 ));
 AND2_X1 \V1/V1/V4/V3/_3_  (.A1(B[7]),
    .A2(A[5]),
    .ZN(\V1/V1/V4/V3/w3 ));
 AND2_X1 \V1/V1/V4/V4/HA1/_0_  (.A1(\V1/V1/V4/V4/w2 ),
    .A2(\V1/V1/V4/V4/w1 ),
    .ZN(\V1/V1/V4/V4/w4 ));
 XOR2_X2 \V1/V1/V4/V4/HA1/_1_  (.A(\V1/V1/V4/V4/w2 ),
    .B(\V1/V1/V4/V4/w1 ),
    .Z(\V1/V1/V4/v4 [1]));
 AND2_X1 \V1/V1/V4/V4/HA2/_0_  (.A1(\V1/V1/V4/V4/w4 ),
    .A2(\V1/V1/V4/V4/w3 ),
    .ZN(\V1/V1/V4/v4 [3]));
 XOR2_X2 \V1/V1/V4/V4/HA2/_1_  (.A(\V1/V1/V4/V4/w4 ),
    .B(\V1/V1/V4/V4/w3 ),
    .Z(\V1/V1/V4/v4 [2]));
 AND2_X1 \V1/V1/V4/V4/_0_  (.A1(A[6]),
    .A2(B[6]),
    .ZN(\V1/V1/V4/v4 [0]));
 AND2_X1 \V1/V1/V4/V4/_1_  (.A1(A[6]),
    .A2(B[7]),
    .ZN(\V1/V1/V4/V4/w1 ));
 AND2_X1 \V1/V1/V4/V4/_2_  (.A1(B[6]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V4/w2 ));
 AND2_X1 \V1/V1/V4/V4/_3_  (.A1(B[7]),
    .A2(A[7]),
    .ZN(\V1/V1/V4/V4/w3 ));
 OR2_X1 \V1/V1/V4/_0_  (.A1(\V1/V1/V4/c1 ),
    .A2(\V1/V1/V4/c2 ),
    .ZN(\V1/V1/V4/c3 ));
 OR2_X1 \V1/V1/_0_  (.A1(\V1/V1/c1 ),
    .A2(\V1/V1/c2 ),
    .ZN(\V1/V1/c3 ));
 AND2_X1 \V1/V2/A1/A1/M1/M1/_0_  (.A1(\V1/V2/v2 [0]),
    .A2(\V1/V2/v3 [0]),
    .ZN(\V1/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M1/M1/_1_  (.A(\V1/V2/v2 [0]),
    .B(\V1/V2/v3 [0]),
    .Z(\V1/V2/A1/A1/M1/s1 ));
 AND2_X1 \V1/V2/A1/A1/M1/M2/_0_  (.A1(\V1/V2/A1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M1/M2/_1_  (.A(\V1/V2/A1/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/s1 [0]));
 OR2_X1 \V1/V2/A1/A1/M1/_0_  (.A1(\V1/V2/A1/A1/M1/c1 ),
    .A2(\V1/V2/A1/A1/M1/c2 ),
    .ZN(\V1/V2/A1/A1/c1 ));
 AND2_X1 \V1/V2/A1/A1/M2/M1/_0_  (.A1(\V1/V2/v2 [1]),
    .A2(\V1/V2/v3 [1]),
    .ZN(\V1/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M2/M1/_1_  (.A(\V1/V2/v2 [1]),
    .B(\V1/V2/v3 [1]),
    .Z(\V1/V2/A1/A1/M2/s1 ));
 AND2_X1 \V1/V2/A1/A1/M2/M2/_0_  (.A1(\V1/V2/A1/A1/M2/s1 ),
    .A2(\V1/V2/A1/A1/c1 ),
    .ZN(\V1/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M2/M2/_1_  (.A(\V1/V2/A1/A1/M2/s1 ),
    .B(\V1/V2/A1/A1/c1 ),
    .Z(\V1/V2/s1 [1]));
 OR2_X1 \V1/V2/A1/A1/M2/_0_  (.A1(\V1/V2/A1/A1/M2/c1 ),
    .A2(\V1/V2/A1/A1/M2/c2 ),
    .ZN(\V1/V2/A1/A1/c2 ));
 AND2_X1 \V1/V2/A1/A1/M3/M1/_0_  (.A1(\V1/V2/v2 [2]),
    .A2(\V1/V2/v3 [2]),
    .ZN(\V1/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M3/M1/_1_  (.A(\V1/V2/v2 [2]),
    .B(\V1/V2/v3 [2]),
    .Z(\V1/V2/A1/A1/M3/s1 ));
 AND2_X1 \V1/V2/A1/A1/M3/M2/_0_  (.A1(\V1/V2/A1/A1/M3/s1 ),
    .A2(\V1/V2/A1/A1/c2 ),
    .ZN(\V1/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M3/M2/_1_  (.A(\V1/V2/A1/A1/M3/s1 ),
    .B(\V1/V2/A1/A1/c2 ),
    .Z(\V1/V2/s1 [2]));
 OR2_X1 \V1/V2/A1/A1/M3/_0_  (.A1(\V1/V2/A1/A1/M3/c1 ),
    .A2(\V1/V2/A1/A1/M3/c2 ),
    .ZN(\V1/V2/A1/A1/c3 ));
 AND2_X1 \V1/V2/A1/A1/M4/M1/_0_  (.A1(\V1/V2/v2 [3]),
    .A2(\V1/V2/v3 [3]),
    .ZN(\V1/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A1/A1/M4/M1/_1_  (.A(\V1/V2/v2 [3]),
    .B(\V1/V2/v3 [3]),
    .Z(\V1/V2/A1/A1/M4/s1 ));
 AND2_X1 \V1/V2/A1/A1/M4/M2/_0_  (.A1(\V1/V2/A1/A1/M4/s1 ),
    .A2(\V1/V2/A1/A1/c3 ),
    .ZN(\V1/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A1/A1/M4/M2/_1_  (.A(\V1/V2/A1/A1/M4/s1 ),
    .B(\V1/V2/A1/A1/c3 ),
    .Z(\V1/V2/s1 [3]));
 OR2_X1 \V1/V2/A1/A1/M4/_0_  (.A1(\V1/V2/A1/A1/M4/c1 ),
    .A2(\V1/V2/A1/A1/M4/c2 ),
    .ZN(\V1/V2/A1/c1 ));
 AND2_X1 \V1/V2/A1/A2/M1/M1/_0_  (.A1(\V1/V2/v2 [4]),
    .A2(\V1/V2/v3 [4]),
    .ZN(\V1/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M1/M1/_1_  (.A(\V1/V2/v2 [4]),
    .B(\V1/V2/v3 [4]),
    .Z(\V1/V2/A1/A2/M1/s1 ));
 AND2_X1 \V1/V2/A1/A2/M1/M2/_0_  (.A1(\V1/V2/A1/A2/M1/s1 ),
    .A2(\V1/V2/A1/c1 ),
    .ZN(\V1/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M1/M2/_1_  (.A(\V1/V2/A1/A2/M1/s1 ),
    .B(\V1/V2/A1/c1 ),
    .Z(\V1/V2/s1 [4]));
 OR2_X1 \V1/V2/A1/A2/M1/_0_  (.A1(\V1/V2/A1/A2/M1/c1 ),
    .A2(\V1/V2/A1/A2/M1/c2 ),
    .ZN(\V1/V2/A1/A2/c1 ));
 AND2_X1 \V1/V2/A1/A2/M2/M1/_0_  (.A1(\V1/V2/v2 [5]),
    .A2(\V1/V2/v3 [5]),
    .ZN(\V1/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M2/M1/_1_  (.A(\V1/V2/v2 [5]),
    .B(\V1/V2/v3 [5]),
    .Z(\V1/V2/A1/A2/M2/s1 ));
 AND2_X1 \V1/V2/A1/A2/M2/M2/_0_  (.A1(\V1/V2/A1/A2/M2/s1 ),
    .A2(\V1/V2/A1/A2/c1 ),
    .ZN(\V1/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M2/M2/_1_  (.A(\V1/V2/A1/A2/M2/s1 ),
    .B(\V1/V2/A1/A2/c1 ),
    .Z(\V1/V2/s1 [5]));
 OR2_X1 \V1/V2/A1/A2/M2/_0_  (.A1(\V1/V2/A1/A2/M2/c1 ),
    .A2(\V1/V2/A1/A2/M2/c2 ),
    .ZN(\V1/V2/A1/A2/c2 ));
 AND2_X1 \V1/V2/A1/A2/M3/M1/_0_  (.A1(\V1/V2/v2 [6]),
    .A2(\V1/V2/v3 [6]),
    .ZN(\V1/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M3/M1/_1_  (.A(\V1/V2/v2 [6]),
    .B(\V1/V2/v3 [6]),
    .Z(\V1/V2/A1/A2/M3/s1 ));
 AND2_X1 \V1/V2/A1/A2/M3/M2/_0_  (.A1(\V1/V2/A1/A2/M3/s1 ),
    .A2(\V1/V2/A1/A2/c2 ),
    .ZN(\V1/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M3/M2/_1_  (.A(\V1/V2/A1/A2/M3/s1 ),
    .B(\V1/V2/A1/A2/c2 ),
    .Z(\V1/V2/s1 [6]));
 OR2_X1 \V1/V2/A1/A2/M3/_0_  (.A1(\V1/V2/A1/A2/M3/c1 ),
    .A2(\V1/V2/A1/A2/M3/c2 ),
    .ZN(\V1/V2/A1/A2/c3 ));
 AND2_X1 \V1/V2/A1/A2/M4/M1/_0_  (.A1(\V1/V2/v2 [7]),
    .A2(\V1/V2/v3 [7]),
    .ZN(\V1/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A1/A2/M4/M1/_1_  (.A(\V1/V2/v2 [7]),
    .B(\V1/V2/v3 [7]),
    .Z(\V1/V2/A1/A2/M4/s1 ));
 AND2_X1 \V1/V2/A1/A2/M4/M2/_0_  (.A1(\V1/V2/A1/A2/M4/s1 ),
    .A2(\V1/V2/A1/A2/c3 ),
    .ZN(\V1/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A1/A2/M4/M2/_1_  (.A(\V1/V2/A1/A2/M4/s1 ),
    .B(\V1/V2/A1/A2/c3 ),
    .Z(\V1/V2/s1 [7]));
 OR2_X1 \V1/V2/A1/A2/M4/_0_  (.A1(\V1/V2/A1/A2/M4/c1 ),
    .A2(\V1/V2/A1/A2/M4/c2 ),
    .ZN(\V1/V2/c1 ));
 AND2_X1 \V1/V2/A2/A1/M1/M1/_0_  (.A1(\V1/V2/s1 [0]),
    .A2(\V1/V2/v1 [4]),
    .ZN(\V1/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M1/M1/_1_  (.A(\V1/V2/s1 [0]),
    .B(\V1/V2/v1 [4]),
    .Z(\V1/V2/A2/A1/M1/s1 ));
 AND2_X1 \V1/V2/A2/A1/M1/M2/_0_  (.A1(\V1/V2/A2/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M1/M2/_1_  (.A(\V1/V2/A2/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/v2 [4]));
 OR2_X1 \V1/V2/A2/A1/M1/_0_  (.A1(\V1/V2/A2/A1/M1/c1 ),
    .A2(\V1/V2/A2/A1/M1/c2 ),
    .ZN(\V1/V2/A2/A1/c1 ));
 AND2_X1 \V1/V2/A2/A1/M2/M1/_0_  (.A1(\V1/V2/s1 [1]),
    .A2(\V1/V2/v1 [5]),
    .ZN(\V1/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M2/M1/_1_  (.A(\V1/V2/s1 [1]),
    .B(\V1/V2/v1 [5]),
    .Z(\V1/V2/A2/A1/M2/s1 ));
 AND2_X1 \V1/V2/A2/A1/M2/M2/_0_  (.A1(\V1/V2/A2/A1/M2/s1 ),
    .A2(\V1/V2/A2/A1/c1 ),
    .ZN(\V1/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M2/M2/_1_  (.A(\V1/V2/A2/A1/M2/s1 ),
    .B(\V1/V2/A2/A1/c1 ),
    .Z(\V1/v2 [5]));
 OR2_X1 \V1/V2/A2/A1/M2/_0_  (.A1(\V1/V2/A2/A1/M2/c1 ),
    .A2(\V1/V2/A2/A1/M2/c2 ),
    .ZN(\V1/V2/A2/A1/c2 ));
 AND2_X1 \V1/V2/A2/A1/M3/M1/_0_  (.A1(\V1/V2/s1 [2]),
    .A2(\V1/V2/v1 [6]),
    .ZN(\V1/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M3/M1/_1_  (.A(\V1/V2/s1 [2]),
    .B(\V1/V2/v1 [6]),
    .Z(\V1/V2/A2/A1/M3/s1 ));
 AND2_X1 \V1/V2/A2/A1/M3/M2/_0_  (.A1(\V1/V2/A2/A1/M3/s1 ),
    .A2(\V1/V2/A2/A1/c2 ),
    .ZN(\V1/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M3/M2/_1_  (.A(\V1/V2/A2/A1/M3/s1 ),
    .B(\V1/V2/A2/A1/c2 ),
    .Z(\V1/v2 [6]));
 OR2_X1 \V1/V2/A2/A1/M3/_0_  (.A1(\V1/V2/A2/A1/M3/c1 ),
    .A2(\V1/V2/A2/A1/M3/c2 ),
    .ZN(\V1/V2/A2/A1/c3 ));
 AND2_X1 \V1/V2/A2/A1/M4/M1/_0_  (.A1(\V1/V2/s1 [3]),
    .A2(\V1/V2/v1 [7]),
    .ZN(\V1/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A2/A1/M4/M1/_1_  (.A(\V1/V2/s1 [3]),
    .B(\V1/V2/v1 [7]),
    .Z(\V1/V2/A2/A1/M4/s1 ));
 AND2_X1 \V1/V2/A2/A1/M4/M2/_0_  (.A1(\V1/V2/A2/A1/M4/s1 ),
    .A2(\V1/V2/A2/A1/c3 ),
    .ZN(\V1/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A2/A1/M4/M2/_1_  (.A(\V1/V2/A2/A1/M4/s1 ),
    .B(\V1/V2/A2/A1/c3 ),
    .Z(\V1/v2 [7]));
 OR2_X1 \V1/V2/A2/A1/M4/_0_  (.A1(\V1/V2/A2/A1/M4/c1 ),
    .A2(\V1/V2/A2/A1/M4/c2 ),
    .ZN(\V1/V2/A2/c1 ));
 AND2_X1 \V1/V2/A2/A2/M1/M1/_0_  (.A1(\V1/V2/s1 [4]),
    .A2(net3),
    .ZN(\V1/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M1/M1/_1_  (.A(\V1/V2/s1 [4]),
    .B(net3),
    .Z(\V1/V2/A2/A2/M1/s1 ));
 AND2_X1 \V1/V2/A2/A2/M1/M2/_0_  (.A1(\V1/V2/A2/A2/M1/s1 ),
    .A2(\V1/V2/A2/c1 ),
    .ZN(\V1/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M1/M2/_1_  (.A(\V1/V2/A2/A2/M1/s1 ),
    .B(\V1/V2/A2/c1 ),
    .Z(\V1/V2/s2 [4]));
 OR2_X1 \V1/V2/A2/A2/M1/_0_  (.A1(\V1/V2/A2/A2/M1/c1 ),
    .A2(\V1/V2/A2/A2/M1/c2 ),
    .ZN(\V1/V2/A2/A2/c1 ));
 AND2_X1 \V1/V2/A2/A2/M2/M1/_0_  (.A1(\V1/V2/s1 [5]),
    .A2(net3),
    .ZN(\V1/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M2/M1/_1_  (.A(\V1/V2/s1 [5]),
    .B(net3),
    .Z(\V1/V2/A2/A2/M2/s1 ));
 AND2_X1 \V1/V2/A2/A2/M2/M2/_0_  (.A1(\V1/V2/A2/A2/M2/s1 ),
    .A2(\V1/V2/A2/A2/c1 ),
    .ZN(\V1/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M2/M2/_1_  (.A(\V1/V2/A2/A2/M2/s1 ),
    .B(\V1/V2/A2/A2/c1 ),
    .Z(\V1/V2/s2 [5]));
 OR2_X1 \V1/V2/A2/A2/M2/_0_  (.A1(\V1/V2/A2/A2/M2/c1 ),
    .A2(\V1/V2/A2/A2/M2/c2 ),
    .ZN(\V1/V2/A2/A2/c2 ));
 AND2_X1 \V1/V2/A2/A2/M3/M1/_0_  (.A1(\V1/V2/s1 [6]),
    .A2(net3),
    .ZN(\V1/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M3/M1/_1_  (.A(\V1/V2/s1 [6]),
    .B(net3),
    .Z(\V1/V2/A2/A2/M3/s1 ));
 AND2_X1 \V1/V2/A2/A2/M3/M2/_0_  (.A1(\V1/V2/A2/A2/M3/s1 ),
    .A2(\V1/V2/A2/A2/c2 ),
    .ZN(\V1/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M3/M2/_1_  (.A(\V1/V2/A2/A2/M3/s1 ),
    .B(\V1/V2/A2/A2/c2 ),
    .Z(\V1/V2/s2 [6]));
 OR2_X1 \V1/V2/A2/A2/M3/_0_  (.A1(\V1/V2/A2/A2/M3/c1 ),
    .A2(\V1/V2/A2/A2/M3/c2 ),
    .ZN(\V1/V2/A2/A2/c3 ));
 AND2_X1 \V1/V2/A2/A2/M4/M1/_0_  (.A1(\V1/V2/s1 [7]),
    .A2(net3),
    .ZN(\V1/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A2/A2/M4/M1/_1_  (.A(\V1/V2/s1 [7]),
    .B(net3),
    .Z(\V1/V2/A2/A2/M4/s1 ));
 AND2_X1 \V1/V2/A2/A2/M4/M2/_0_  (.A1(\V1/V2/A2/A2/M4/s1 ),
    .A2(\V1/V2/A2/A2/c3 ),
    .ZN(\V1/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A2/A2/M4/M2/_1_  (.A(\V1/V2/A2/A2/M4/s1 ),
    .B(\V1/V2/A2/A2/c3 ),
    .Z(\V1/V2/s2 [7]));
 OR2_X1 \V1/V2/A2/A2/M4/_0_  (.A1(\V1/V2/A2/A2/M4/c1 ),
    .A2(\V1/V2/A2/A2/M4/c2 ),
    .ZN(\V1/V2/c2 ));
 AND2_X1 \V1/V2/A3/A1/M1/M1/_0_  (.A1(\V1/V2/v4 [0]),
    .A2(\V1/V2/s2 [4]),
    .ZN(\V1/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M1/M1/_1_  (.A(\V1/V2/v4 [0]),
    .B(\V1/V2/s2 [4]),
    .Z(\V1/V2/A3/A1/M1/s1 ));
 AND2_X1 \V1/V2/A3/A1/M1/M2/_0_  (.A1(\V1/V2/A3/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M1/M2/_1_  (.A(\V1/V2/A3/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/v2 [8]));
 OR2_X1 \V1/V2/A3/A1/M1/_0_  (.A1(\V1/V2/A3/A1/M1/c1 ),
    .A2(\V1/V2/A3/A1/M1/c2 ),
    .ZN(\V1/V2/A3/A1/c1 ));
 AND2_X1 \V1/V2/A3/A1/M2/M1/_0_  (.A1(\V1/V2/v4 [1]),
    .A2(\V1/V2/s2 [5]),
    .ZN(\V1/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M2/M1/_1_  (.A(\V1/V2/v4 [1]),
    .B(\V1/V2/s2 [5]),
    .Z(\V1/V2/A3/A1/M2/s1 ));
 AND2_X1 \V1/V2/A3/A1/M2/M2/_0_  (.A1(\V1/V2/A3/A1/M2/s1 ),
    .A2(\V1/V2/A3/A1/c1 ),
    .ZN(\V1/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M2/M2/_1_  (.A(\V1/V2/A3/A1/M2/s1 ),
    .B(\V1/V2/A3/A1/c1 ),
    .Z(\V1/v2 [9]));
 OR2_X1 \V1/V2/A3/A1/M2/_0_  (.A1(\V1/V2/A3/A1/M2/c1 ),
    .A2(\V1/V2/A3/A1/M2/c2 ),
    .ZN(\V1/V2/A3/A1/c2 ));
 AND2_X1 \V1/V2/A3/A1/M3/M1/_0_  (.A1(\V1/V2/v4 [2]),
    .A2(\V1/V2/s2 [6]),
    .ZN(\V1/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M3/M1/_1_  (.A(\V1/V2/v4 [2]),
    .B(\V1/V2/s2 [6]),
    .Z(\V1/V2/A3/A1/M3/s1 ));
 AND2_X1 \V1/V2/A3/A1/M3/M2/_0_  (.A1(\V1/V2/A3/A1/M3/s1 ),
    .A2(\V1/V2/A3/A1/c2 ),
    .ZN(\V1/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M3/M2/_1_  (.A(\V1/V2/A3/A1/M3/s1 ),
    .B(\V1/V2/A3/A1/c2 ),
    .Z(\V1/v2 [10]));
 OR2_X1 \V1/V2/A3/A1/M3/_0_  (.A1(\V1/V2/A3/A1/M3/c1 ),
    .A2(\V1/V2/A3/A1/M3/c2 ),
    .ZN(\V1/V2/A3/A1/c3 ));
 AND2_X1 \V1/V2/A3/A1/M4/M1/_0_  (.A1(\V1/V2/v4 [3]),
    .A2(\V1/V2/s2 [7]),
    .ZN(\V1/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V2/A3/A1/M4/M1/_1_  (.A(\V1/V2/v4 [3]),
    .B(\V1/V2/s2 [7]),
    .Z(\V1/V2/A3/A1/M4/s1 ));
 AND2_X1 \V1/V2/A3/A1/M4/M2/_0_  (.A1(\V1/V2/A3/A1/M4/s1 ),
    .A2(\V1/V2/A3/A1/c3 ),
    .ZN(\V1/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V2/A3/A1/M4/M2/_1_  (.A(\V1/V2/A3/A1/M4/s1 ),
    .B(\V1/V2/A3/A1/c3 ),
    .Z(\V1/v2 [11]));
 OR2_X1 \V1/V2/A3/A1/M4/_0_  (.A1(\V1/V2/A3/A1/M4/c1 ),
    .A2(\V1/V2/A3/A1/M4/c2 ),
    .ZN(\V1/V2/A3/c1 ));
 AND2_X1 \V1/V2/A3/A2/M1/M1/_0_  (.A1(\V1/V2/v4 [4]),
    .A2(\V1/V2/c3 ),
    .ZN(\V1/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M1/M1/_1_  (.A(\V1/V2/v4 [4]),
    .B(\V1/V2/c3 ),
    .Z(\V1/V2/A3/A2/M1/s1 ));
 AND2_X1 \V1/V2/A3/A2/M1/M2/_0_  (.A1(\V1/V2/A3/A2/M1/s1 ),
    .A2(\V1/V2/A3/c1 ),
    .ZN(\V1/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M1/M2/_1_  (.A(\V1/V2/A3/A2/M1/s1 ),
    .B(\V1/V2/A3/c1 ),
    .Z(\V1/v2 [12]));
 OR2_X1 \V1/V2/A3/A2/M1/_0_  (.A1(\V1/V2/A3/A2/M1/c1 ),
    .A2(\V1/V2/A3/A2/M1/c2 ),
    .ZN(\V1/V2/A3/A2/c1 ));
 AND2_X1 \V1/V2/A3/A2/M2/M1/_0_  (.A1(\V1/V2/v4 [5]),
    .A2(net3),
    .ZN(\V1/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M2/M1/_1_  (.A(\V1/V2/v4 [5]),
    .B(net3),
    .Z(\V1/V2/A3/A2/M2/s1 ));
 AND2_X1 \V1/V2/A3/A2/M2/M2/_0_  (.A1(\V1/V2/A3/A2/M2/s1 ),
    .A2(\V1/V2/A3/A2/c1 ),
    .ZN(\V1/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M2/M2/_1_  (.A(\V1/V2/A3/A2/M2/s1 ),
    .B(\V1/V2/A3/A2/c1 ),
    .Z(\V1/v2 [13]));
 OR2_X1 \V1/V2/A3/A2/M2/_0_  (.A1(\V1/V2/A3/A2/M2/c1 ),
    .A2(\V1/V2/A3/A2/M2/c2 ),
    .ZN(\V1/V2/A3/A2/c2 ));
 AND2_X1 \V1/V2/A3/A2/M3/M1/_0_  (.A1(\V1/V2/v4 [6]),
    .A2(net3),
    .ZN(\V1/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M3/M1/_1_  (.A(\V1/V2/v4 [6]),
    .B(net3),
    .Z(\V1/V2/A3/A2/M3/s1 ));
 AND2_X1 \V1/V2/A3/A2/M3/M2/_0_  (.A1(\V1/V2/A3/A2/M3/s1 ),
    .A2(\V1/V2/A3/A2/c2 ),
    .ZN(\V1/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M3/M2/_1_  (.A(\V1/V2/A3/A2/M3/s1 ),
    .B(\V1/V2/A3/A2/c2 ),
    .Z(\V1/v2 [14]));
 OR2_X1 \V1/V2/A3/A2/M3/_0_  (.A1(\V1/V2/A3/A2/M3/c1 ),
    .A2(\V1/V2/A3/A2/M3/c2 ),
    .ZN(\V1/V2/A3/A2/c3 ));
 AND2_X1 \V1/V2/A3/A2/M4/M1/_0_  (.A1(\V1/V2/v4 [7]),
    .A2(net3),
    .ZN(\V1/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V2/A3/A2/M4/M1/_1_  (.A(\V1/V2/v4 [7]),
    .B(net3),
    .Z(\V1/V2/A3/A2/M4/s1 ));
 AND2_X1 \V1/V2/A3/A2/M4/M2/_0_  (.A1(\V1/V2/A3/A2/M4/s1 ),
    .A2(\V1/V2/A3/A2/c3 ),
    .ZN(\V1/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V2/A3/A2/M4/M2/_1_  (.A(\V1/V2/A3/A2/M4/s1 ),
    .B(\V1/V2/A3/A2/c3 ),
    .Z(\V1/v2 [15]));
 OR2_X1 \V1/V2/A3/A2/M4/_0_  (.A1(\V1/V2/A3/A2/M4/c1 ),
    .A2(\V1/V2/A3/A2/M4/c2 ),
    .ZN(\V1/V2/overflow ));
 AND2_X1 \V1/V2/V1/A1/M1/M1/_0_  (.A1(\V1/V2/V1/v2 [0]),
    .A2(\V1/V2/V1/v3 [0]),
    .ZN(\V1/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M1/M1/_1_  (.A(\V1/V2/V1/v2 [0]),
    .B(\V1/V2/V1/v3 [0]),
    .Z(\V1/V2/V1/A1/M1/s1 ));
 AND2_X1 \V1/V2/V1/A1/M1/M2/_0_  (.A1(\V1/V2/V1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M1/M2/_1_  (.A(\V1/V2/V1/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/V1/s1 [0]));
 OR2_X1 \V1/V2/V1/A1/M1/_0_  (.A1(\V1/V2/V1/A1/M1/c1 ),
    .A2(\V1/V2/V1/A1/M1/c2 ),
    .ZN(\V1/V2/V1/A1/c1 ));
 AND2_X1 \V1/V2/V1/A1/M2/M1/_0_  (.A1(\V1/V2/V1/v2 [1]),
    .A2(\V1/V2/V1/v3 [1]),
    .ZN(\V1/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M2/M1/_1_  (.A(\V1/V2/V1/v2 [1]),
    .B(\V1/V2/V1/v3 [1]),
    .Z(\V1/V2/V1/A1/M2/s1 ));
 AND2_X1 \V1/V2/V1/A1/M2/M2/_0_  (.A1(\V1/V2/V1/A1/M2/s1 ),
    .A2(\V1/V2/V1/A1/c1 ),
    .ZN(\V1/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M2/M2/_1_  (.A(\V1/V2/V1/A1/M2/s1 ),
    .B(\V1/V2/V1/A1/c1 ),
    .Z(\V1/V2/V1/s1 [1]));
 OR2_X1 \V1/V2/V1/A1/M2/_0_  (.A1(\V1/V2/V1/A1/M2/c1 ),
    .A2(\V1/V2/V1/A1/M2/c2 ),
    .ZN(\V1/V2/V1/A1/c2 ));
 AND2_X1 \V1/V2/V1/A1/M3/M1/_0_  (.A1(\V1/V2/V1/v2 [2]),
    .A2(\V1/V2/V1/v3 [2]),
    .ZN(\V1/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M3/M1/_1_  (.A(\V1/V2/V1/v2 [2]),
    .B(\V1/V2/V1/v3 [2]),
    .Z(\V1/V2/V1/A1/M3/s1 ));
 AND2_X1 \V1/V2/V1/A1/M3/M2/_0_  (.A1(\V1/V2/V1/A1/M3/s1 ),
    .A2(\V1/V2/V1/A1/c2 ),
    .ZN(\V1/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M3/M2/_1_  (.A(\V1/V2/V1/A1/M3/s1 ),
    .B(\V1/V2/V1/A1/c2 ),
    .Z(\V1/V2/V1/s1 [2]));
 OR2_X1 \V1/V2/V1/A1/M3/_0_  (.A1(\V1/V2/V1/A1/M3/c1 ),
    .A2(\V1/V2/V1/A1/M3/c2 ),
    .ZN(\V1/V2/V1/A1/c3 ));
 AND2_X1 \V1/V2/V1/A1/M4/M1/_0_  (.A1(\V1/V2/V1/v2 [3]),
    .A2(\V1/V2/V1/v3 [3]),
    .ZN(\V1/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A1/M4/M1/_1_  (.A(\V1/V2/V1/v2 [3]),
    .B(\V1/V2/V1/v3 [3]),
    .Z(\V1/V2/V1/A1/M4/s1 ));
 AND2_X1 \V1/V2/V1/A1/M4/M2/_0_  (.A1(\V1/V2/V1/A1/M4/s1 ),
    .A2(\V1/V2/V1/A1/c3 ),
    .ZN(\V1/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A1/M4/M2/_1_  (.A(\V1/V2/V1/A1/M4/s1 ),
    .B(\V1/V2/V1/A1/c3 ),
    .Z(\V1/V2/V1/s1 [3]));
 OR2_X1 \V1/V2/V1/A1/M4/_0_  (.A1(\V1/V2/V1/A1/M4/c1 ),
    .A2(\V1/V2/V1/A1/M4/c2 ),
    .ZN(\V1/V2/V1/c1 ));
 AND2_X1 \V1/V2/V1/A2/M1/M1/_0_  (.A1(\V1/V2/V1/s1 [0]),
    .A2(\V1/V2/V1/v1 [2]),
    .ZN(\V1/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M1/M1/_1_  (.A(\V1/V2/V1/s1 [0]),
    .B(\V1/V2/V1/v1 [2]),
    .Z(\V1/V2/V1/A2/M1/s1 ));
 AND2_X1 \V1/V2/V1/A2/M1/M2/_0_  (.A1(\V1/V2/V1/A2/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M1/M2/_1_  (.A(\V1/V2/V1/A2/M1/s1 ),
    .B(net4),
    .Z(\V1/v2 [2]));
 OR2_X1 \V1/V2/V1/A2/M1/_0_  (.A1(\V1/V2/V1/A2/M1/c1 ),
    .A2(\V1/V2/V1/A2/M1/c2 ),
    .ZN(\V1/V2/V1/A2/c1 ));
 AND2_X1 \V1/V2/V1/A2/M2/M1/_0_  (.A1(\V1/V2/V1/s1 [1]),
    .A2(\V1/V2/V1/v1 [3]),
    .ZN(\V1/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M2/M1/_1_  (.A(\V1/V2/V1/s1 [1]),
    .B(\V1/V2/V1/v1 [3]),
    .Z(\V1/V2/V1/A2/M2/s1 ));
 AND2_X1 \V1/V2/V1/A2/M2/M2/_0_  (.A1(\V1/V2/V1/A2/M2/s1 ),
    .A2(\V1/V2/V1/A2/c1 ),
    .ZN(\V1/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M2/M2/_1_  (.A(\V1/V2/V1/A2/M2/s1 ),
    .B(\V1/V2/V1/A2/c1 ),
    .Z(\V1/v2 [3]));
 OR2_X1 \V1/V2/V1/A2/M2/_0_  (.A1(\V1/V2/V1/A2/M2/c1 ),
    .A2(\V1/V2/V1/A2/M2/c2 ),
    .ZN(\V1/V2/V1/A2/c2 ));
 AND2_X1 \V1/V2/V1/A2/M3/M1/_0_  (.A1(\V1/V2/V1/s1 [2]),
    .A2(net3),
    .ZN(\V1/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M3/M1/_1_  (.A(\V1/V2/V1/s1 [2]),
    .B(net3),
    .Z(\V1/V2/V1/A2/M3/s1 ));
 AND2_X1 \V1/V2/V1/A2/M3/M2/_0_  (.A1(\V1/V2/V1/A2/M3/s1 ),
    .A2(\V1/V2/V1/A2/c2 ),
    .ZN(\V1/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M3/M2/_1_  (.A(\V1/V2/V1/A2/M3/s1 ),
    .B(\V1/V2/V1/A2/c2 ),
    .Z(\V1/V2/V1/s2 [2]));
 OR2_X1 \V1/V2/V1/A2/M3/_0_  (.A1(\V1/V2/V1/A2/M3/c1 ),
    .A2(\V1/V2/V1/A2/M3/c2 ),
    .ZN(\V1/V2/V1/A2/c3 ));
 AND2_X1 \V1/V2/V1/A2/M4/M1/_0_  (.A1(\V1/V2/V1/s1 [3]),
    .A2(net3),
    .ZN(\V1/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A2/M4/M1/_1_  (.A(\V1/V2/V1/s1 [3]),
    .B(net3),
    .Z(\V1/V2/V1/A2/M4/s1 ));
 AND2_X1 \V1/V2/V1/A2/M4/M2/_0_  (.A1(\V1/V2/V1/A2/M4/s1 ),
    .A2(\V1/V2/V1/A2/c3 ),
    .ZN(\V1/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A2/M4/M2/_1_  (.A(\V1/V2/V1/A2/M4/s1 ),
    .B(\V1/V2/V1/A2/c3 ),
    .Z(\V1/V2/V1/s2 [3]));
 OR2_X1 \V1/V2/V1/A2/M4/_0_  (.A1(\V1/V2/V1/A2/M4/c1 ),
    .A2(\V1/V2/V1/A2/M4/c2 ),
    .ZN(\V1/V2/V1/c2 ));
 AND2_X1 \V1/V2/V1/A3/M1/M1/_0_  (.A1(\V1/V2/V1/v4 [0]),
    .A2(\V1/V2/V1/s2 [2]),
    .ZN(\V1/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M1/M1/_1_  (.A(\V1/V2/V1/v4 [0]),
    .B(\V1/V2/V1/s2 [2]),
    .Z(\V1/V2/V1/A3/M1/s1 ));
 AND2_X1 \V1/V2/V1/A3/M1/M2/_0_  (.A1(\V1/V2/V1/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M1/M2/_1_  (.A(\V1/V2/V1/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v1 [4]));
 OR2_X1 \V1/V2/V1/A3/M1/_0_  (.A1(\V1/V2/V1/A3/M1/c1 ),
    .A2(\V1/V2/V1/A3/M1/c2 ),
    .ZN(\V1/V2/V1/A3/c1 ));
 AND2_X1 \V1/V2/V1/A3/M2/M1/_0_  (.A1(\V1/V2/V1/v4 [1]),
    .A2(\V1/V2/V1/s2 [3]),
    .ZN(\V1/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M2/M1/_1_  (.A(\V1/V2/V1/v4 [1]),
    .B(\V1/V2/V1/s2 [3]),
    .Z(\V1/V2/V1/A3/M2/s1 ));
 AND2_X1 \V1/V2/V1/A3/M2/M2/_0_  (.A1(\V1/V2/V1/A3/M2/s1 ),
    .A2(\V1/V2/V1/A3/c1 ),
    .ZN(\V1/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M2/M2/_1_  (.A(\V1/V2/V1/A3/M2/s1 ),
    .B(\V1/V2/V1/A3/c1 ),
    .Z(\V1/V2/v1 [5]));
 OR2_X1 \V1/V2/V1/A3/M2/_0_  (.A1(\V1/V2/V1/A3/M2/c1 ),
    .A2(\V1/V2/V1/A3/M2/c2 ),
    .ZN(\V1/V2/V1/A3/c2 ));
 AND2_X1 \V1/V2/V1/A3/M3/M1/_0_  (.A1(\V1/V2/V1/v4 [2]),
    .A2(\V1/V2/V1/c3 ),
    .ZN(\V1/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M3/M1/_1_  (.A(\V1/V2/V1/v4 [2]),
    .B(\V1/V2/V1/c3 ),
    .Z(\V1/V2/V1/A3/M3/s1 ));
 AND2_X1 \V1/V2/V1/A3/M3/M2/_0_  (.A1(\V1/V2/V1/A3/M3/s1 ),
    .A2(\V1/V2/V1/A3/c2 ),
    .ZN(\V1/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M3/M2/_1_  (.A(\V1/V2/V1/A3/M3/s1 ),
    .B(\V1/V2/V1/A3/c2 ),
    .Z(\V1/V2/v1 [6]));
 OR2_X1 \V1/V2/V1/A3/M3/_0_  (.A1(\V1/V2/V1/A3/M3/c1 ),
    .A2(\V1/V2/V1/A3/M3/c2 ),
    .ZN(\V1/V2/V1/A3/c3 ));
 AND2_X1 \V1/V2/V1/A3/M4/M1/_0_  (.A1(\V1/V2/V1/v4 [3]),
    .A2(net3),
    .ZN(\V1/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V1/A3/M4/M1/_1_  (.A(\V1/V2/V1/v4 [3]),
    .B(net3),
    .Z(\V1/V2/V1/A3/M4/s1 ));
 AND2_X1 \V1/V2/V1/A3/M4/M2/_0_  (.A1(\V1/V2/V1/A3/M4/s1 ),
    .A2(\V1/V2/V1/A3/c3 ),
    .ZN(\V1/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V1/A3/M4/M2/_1_  (.A(\V1/V2/V1/A3/M4/s1 ),
    .B(\V1/V2/V1/A3/c3 ),
    .Z(\V1/V2/v1 [7]));
 OR2_X1 \V1/V2/V1/A3/M4/_0_  (.A1(\V1/V2/V1/A3/M4/c1 ),
    .A2(\V1/V2/V1/A3/M4/c2 ),
    .ZN(\V1/V2/V1/overflow ));
 AND2_X1 \V1/V2/V1/V1/HA1/_0_  (.A1(\V1/V2/V1/V1/w2 ),
    .A2(\V1/V2/V1/V1/w1 ),
    .ZN(\V1/V2/V1/V1/w4 ));
 XOR2_X2 \V1/V2/V1/V1/HA1/_1_  (.A(\V1/V2/V1/V1/w2 ),
    .B(\V1/V2/V1/V1/w1 ),
    .Z(\V1/v2 [1]));
 AND2_X1 \V1/V2/V1/V1/HA2/_0_  (.A1(\V1/V2/V1/V1/w4 ),
    .A2(\V1/V2/V1/V1/w3 ),
    .ZN(\V1/V2/V1/v1 [3]));
 XOR2_X2 \V1/V2/V1/V1/HA2/_1_  (.A(\V1/V2/V1/V1/w4 ),
    .B(\V1/V2/V1/V1/w3 ),
    .Z(\V1/V2/V1/v1 [2]));
 AND2_X1 \V1/V2/V1/V1/_0_  (.A1(net25),
    .A2(net23),
    .ZN(\V1/v2 [0]));
 AND2_X1 \V1/V2/V1/V1/_1_  (.A1(net25),
    .A2(B[1]),
    .ZN(\V1/V2/V1/V1/w1 ));
 AND2_X1 \V1/V2/V1/V1/_2_  (.A1(net23),
    .A2(net24),
    .ZN(\V1/V2/V1/V1/w2 ));
 AND2_X1 \V1/V2/V1/V1/_3_  (.A1(B[1]),
    .A2(net24),
    .ZN(\V1/V2/V1/V1/w3 ));
 AND2_X1 \V1/V2/V1/V2/HA1/_0_  (.A1(\V1/V2/V1/V2/w2 ),
    .A2(\V1/V2/V1/V2/w1 ),
    .ZN(\V1/V2/V1/V2/w4 ));
 XOR2_X2 \V1/V2/V1/V2/HA1/_1_  (.A(\V1/V2/V1/V2/w2 ),
    .B(\V1/V2/V1/V2/w1 ),
    .Z(\V1/V2/V1/v2 [1]));
 AND2_X1 \V1/V2/V1/V2/HA2/_0_  (.A1(\V1/V2/V1/V2/w4 ),
    .A2(\V1/V2/V1/V2/w3 ),
    .ZN(\V1/V2/V1/v2 [3]));
 XOR2_X2 \V1/V2/V1/V2/HA2/_1_  (.A(\V1/V2/V1/V2/w4 ),
    .B(\V1/V2/V1/V2/w3 ),
    .Z(\V1/V2/V1/v2 [2]));
 AND2_X1 \V1/V2/V1/V2/_0_  (.A1(net47),
    .A2(B[0]),
    .ZN(\V1/V2/V1/v2 [0]));
 AND2_X1 \V1/V2/V1/V2/_1_  (.A1(net47),
    .A2(B[1]),
    .ZN(\V1/V2/V1/V2/w1 ));
 AND2_X1 \V1/V2/V1/V2/_2_  (.A1(B[0]),
    .A2(net46),
    .ZN(\V1/V2/V1/V2/w2 ));
 AND2_X1 \V1/V2/V1/V2/_3_  (.A1(B[1]),
    .A2(net46),
    .ZN(\V1/V2/V1/V2/w3 ));
 AND2_X1 \V1/V2/V1/V3/HA1/_0_  (.A1(\V1/V2/V1/V3/w2 ),
    .A2(\V1/V2/V1/V3/w1 ),
    .ZN(\V1/V2/V1/V3/w4 ));
 XOR2_X2 \V1/V2/V1/V3/HA1/_1_  (.A(\V1/V2/V1/V3/w2 ),
    .B(\V1/V2/V1/V3/w1 ),
    .Z(\V1/V2/V1/v3 [1]));
 AND2_X1 \V1/V2/V1/V3/HA2/_0_  (.A1(\V1/V2/V1/V3/w4 ),
    .A2(\V1/V2/V1/V3/w3 ),
    .ZN(\V1/V2/V1/v3 [3]));
 XOR2_X2 \V1/V2/V1/V3/HA2/_1_  (.A(\V1/V2/V1/V3/w4 ),
    .B(\V1/V2/V1/V3/w3 ),
    .Z(\V1/V2/V1/v3 [2]));
 AND2_X1 \V1/V2/V1/V3/_0_  (.A1(net25),
    .A2(B[2]),
    .ZN(\V1/V2/V1/v3 [0]));
 AND2_X1 \V1/V2/V1/V3/_1_  (.A1(net25),
    .A2(B[3]),
    .ZN(\V1/V2/V1/V3/w1 ));
 AND2_X1 \V1/V2/V1/V3/_2_  (.A1(B[2]),
    .A2(net24),
    .ZN(\V1/V2/V1/V3/w2 ));
 AND2_X1 \V1/V2/V1/V3/_3_  (.A1(B[3]),
    .A2(net24),
    .ZN(\V1/V2/V1/V3/w3 ));
 AND2_X1 \V1/V2/V1/V4/HA1/_0_  (.A1(\V1/V2/V1/V4/w2 ),
    .A2(\V1/V2/V1/V4/w1 ),
    .ZN(\V1/V2/V1/V4/w4 ));
 XOR2_X2 \V1/V2/V1/V4/HA1/_1_  (.A(\V1/V2/V1/V4/w2 ),
    .B(\V1/V2/V1/V4/w1 ),
    .Z(\V1/V2/V1/v4 [1]));
 AND2_X1 \V1/V2/V1/V4/HA2/_0_  (.A1(\V1/V2/V1/V4/w4 ),
    .A2(\V1/V2/V1/V4/w3 ),
    .ZN(\V1/V2/V1/v4 [3]));
 XOR2_X2 \V1/V2/V1/V4/HA2/_1_  (.A(\V1/V2/V1/V4/w4 ),
    .B(\V1/V2/V1/V4/w3 ),
    .Z(\V1/V2/V1/v4 [2]));
 AND2_X1 \V1/V2/V1/V4/_0_  (.A1(net47),
    .A2(B[2]),
    .ZN(\V1/V2/V1/v4 [0]));
 AND2_X1 \V1/V2/V1/V4/_1_  (.A1(net47),
    .A2(B[3]),
    .ZN(\V1/V2/V1/V4/w1 ));
 AND2_X1 \V1/V2/V1/V4/_2_  (.A1(B[2]),
    .A2(net46),
    .ZN(\V1/V2/V1/V4/w2 ));
 AND2_X1 \V1/V2/V1/V4/_3_  (.A1(B[3]),
    .A2(net46),
    .ZN(\V1/V2/V1/V4/w3 ));
 OR2_X1 \V1/V2/V1/_0_  (.A1(\V1/V2/V1/c1 ),
    .A2(\V1/V2/V1/c2 ),
    .ZN(\V1/V2/V1/c3 ));
 AND2_X1 \V1/V2/V2/A1/M1/M1/_0_  (.A1(\V1/V2/V2/v2 [0]),
    .A2(\V1/V2/V2/v3 [0]),
    .ZN(\V1/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M1/M1/_1_  (.A(\V1/V2/V2/v2 [0]),
    .B(\V1/V2/V2/v3 [0]),
    .Z(\V1/V2/V2/A1/M1/s1 ));
 AND2_X1 \V1/V2/V2/A1/M1/M2/_0_  (.A1(\V1/V2/V2/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M1/M2/_1_  (.A(\V1/V2/V2/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/V2/s1 [0]));
 OR2_X1 \V1/V2/V2/A1/M1/_0_  (.A1(\V1/V2/V2/A1/M1/c1 ),
    .A2(\V1/V2/V2/A1/M1/c2 ),
    .ZN(\V1/V2/V2/A1/c1 ));
 AND2_X1 \V1/V2/V2/A1/M2/M1/_0_  (.A1(\V1/V2/V2/v2 [1]),
    .A2(\V1/V2/V2/v3 [1]),
    .ZN(\V1/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M2/M1/_1_  (.A(\V1/V2/V2/v2 [1]),
    .B(\V1/V2/V2/v3 [1]),
    .Z(\V1/V2/V2/A1/M2/s1 ));
 AND2_X1 \V1/V2/V2/A1/M2/M2/_0_  (.A1(\V1/V2/V2/A1/M2/s1 ),
    .A2(\V1/V2/V2/A1/c1 ),
    .ZN(\V1/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M2/M2/_1_  (.A(\V1/V2/V2/A1/M2/s1 ),
    .B(\V1/V2/V2/A1/c1 ),
    .Z(\V1/V2/V2/s1 [1]));
 OR2_X1 \V1/V2/V2/A1/M2/_0_  (.A1(\V1/V2/V2/A1/M2/c1 ),
    .A2(\V1/V2/V2/A1/M2/c2 ),
    .ZN(\V1/V2/V2/A1/c2 ));
 AND2_X1 \V1/V2/V2/A1/M3/M1/_0_  (.A1(\V1/V2/V2/v2 [2]),
    .A2(\V1/V2/V2/v3 [2]),
    .ZN(\V1/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M3/M1/_1_  (.A(\V1/V2/V2/v2 [2]),
    .B(\V1/V2/V2/v3 [2]),
    .Z(\V1/V2/V2/A1/M3/s1 ));
 AND2_X1 \V1/V2/V2/A1/M3/M2/_0_  (.A1(\V1/V2/V2/A1/M3/s1 ),
    .A2(\V1/V2/V2/A1/c2 ),
    .ZN(\V1/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M3/M2/_1_  (.A(\V1/V2/V2/A1/M3/s1 ),
    .B(\V1/V2/V2/A1/c2 ),
    .Z(\V1/V2/V2/s1 [2]));
 OR2_X1 \V1/V2/V2/A1/M3/_0_  (.A1(\V1/V2/V2/A1/M3/c1 ),
    .A2(\V1/V2/V2/A1/M3/c2 ),
    .ZN(\V1/V2/V2/A1/c3 ));
 AND2_X1 \V1/V2/V2/A1/M4/M1/_0_  (.A1(\V1/V2/V2/v2 [3]),
    .A2(\V1/V2/V2/v3 [3]),
    .ZN(\V1/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A1/M4/M1/_1_  (.A(\V1/V2/V2/v2 [3]),
    .B(\V1/V2/V2/v3 [3]),
    .Z(\V1/V2/V2/A1/M4/s1 ));
 AND2_X1 \V1/V2/V2/A1/M4/M2/_0_  (.A1(\V1/V2/V2/A1/M4/s1 ),
    .A2(\V1/V2/V2/A1/c3 ),
    .ZN(\V1/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A1/M4/M2/_1_  (.A(\V1/V2/V2/A1/M4/s1 ),
    .B(\V1/V2/V2/A1/c3 ),
    .Z(\V1/V2/V2/s1 [3]));
 OR2_X1 \V1/V2/V2/A1/M4/_0_  (.A1(\V1/V2/V2/A1/M4/c1 ),
    .A2(\V1/V2/V2/A1/M4/c2 ),
    .ZN(\V1/V2/V2/c1 ));
 AND2_X1 \V1/V2/V2/A2/M1/M1/_0_  (.A1(\V1/V2/V2/s1 [0]),
    .A2(\V1/V2/V2/v1 [2]),
    .ZN(\V1/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M1/M1/_1_  (.A(\V1/V2/V2/s1 [0]),
    .B(\V1/V2/V2/v1 [2]),
    .Z(\V1/V2/V2/A2/M1/s1 ));
 AND2_X1 \V1/V2/V2/A2/M1/M2/_0_  (.A1(\V1/V2/V2/A2/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M1/M2/_1_  (.A(\V1/V2/V2/A2/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v2 [2]));
 OR2_X1 \V1/V2/V2/A2/M1/_0_  (.A1(\V1/V2/V2/A2/M1/c1 ),
    .A2(\V1/V2/V2/A2/M1/c2 ),
    .ZN(\V1/V2/V2/A2/c1 ));
 AND2_X1 \V1/V2/V2/A2/M2/M1/_0_  (.A1(\V1/V2/V2/s1 [1]),
    .A2(\V1/V2/V2/v1 [3]),
    .ZN(\V1/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M2/M1/_1_  (.A(\V1/V2/V2/s1 [1]),
    .B(\V1/V2/V2/v1 [3]),
    .Z(\V1/V2/V2/A2/M2/s1 ));
 AND2_X1 \V1/V2/V2/A2/M2/M2/_0_  (.A1(\V1/V2/V2/A2/M2/s1 ),
    .A2(\V1/V2/V2/A2/c1 ),
    .ZN(\V1/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M2/M2/_1_  (.A(\V1/V2/V2/A2/M2/s1 ),
    .B(\V1/V2/V2/A2/c1 ),
    .Z(\V1/V2/v2 [3]));
 OR2_X1 \V1/V2/V2/A2/M2/_0_  (.A1(\V1/V2/V2/A2/M2/c1 ),
    .A2(\V1/V2/V2/A2/M2/c2 ),
    .ZN(\V1/V2/V2/A2/c2 ));
 AND2_X1 \V1/V2/V2/A2/M3/M1/_0_  (.A1(\V1/V2/V2/s1 [2]),
    .A2(net3),
    .ZN(\V1/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M3/M1/_1_  (.A(\V1/V2/V2/s1 [2]),
    .B(net3),
    .Z(\V1/V2/V2/A2/M3/s1 ));
 AND2_X1 \V1/V2/V2/A2/M3/M2/_0_  (.A1(\V1/V2/V2/A2/M3/s1 ),
    .A2(\V1/V2/V2/A2/c2 ),
    .ZN(\V1/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M3/M2/_1_  (.A(\V1/V2/V2/A2/M3/s1 ),
    .B(\V1/V2/V2/A2/c2 ),
    .Z(\V1/V2/V2/s2 [2]));
 OR2_X1 \V1/V2/V2/A2/M3/_0_  (.A1(\V1/V2/V2/A2/M3/c1 ),
    .A2(\V1/V2/V2/A2/M3/c2 ),
    .ZN(\V1/V2/V2/A2/c3 ));
 AND2_X1 \V1/V2/V2/A2/M4/M1/_0_  (.A1(\V1/V2/V2/s1 [3]),
    .A2(net3),
    .ZN(\V1/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A2/M4/M1/_1_  (.A(\V1/V2/V2/s1 [3]),
    .B(net3),
    .Z(\V1/V2/V2/A2/M4/s1 ));
 AND2_X1 \V1/V2/V2/A2/M4/M2/_0_  (.A1(\V1/V2/V2/A2/M4/s1 ),
    .A2(\V1/V2/V2/A2/c3 ),
    .ZN(\V1/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A2/M4/M2/_1_  (.A(\V1/V2/V2/A2/M4/s1 ),
    .B(\V1/V2/V2/A2/c3 ),
    .Z(\V1/V2/V2/s2 [3]));
 OR2_X1 \V1/V2/V2/A2/M4/_0_  (.A1(\V1/V2/V2/A2/M4/c1 ),
    .A2(\V1/V2/V2/A2/M4/c2 ),
    .ZN(\V1/V2/V2/c2 ));
 AND2_X1 \V1/V2/V2/A3/M1/M1/_0_  (.A1(\V1/V2/V2/v4 [0]),
    .A2(\V1/V2/V2/s2 [2]),
    .ZN(\V1/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M1/M1/_1_  (.A(\V1/V2/V2/v4 [0]),
    .B(\V1/V2/V2/s2 [2]),
    .Z(\V1/V2/V2/A3/M1/s1 ));
 AND2_X1 \V1/V2/V2/A3/M1/M2/_0_  (.A1(\V1/V2/V2/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M1/M2/_1_  (.A(\V1/V2/V2/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v2 [4]));
 OR2_X1 \V1/V2/V2/A3/M1/_0_  (.A1(\V1/V2/V2/A3/M1/c1 ),
    .A2(\V1/V2/V2/A3/M1/c2 ),
    .ZN(\V1/V2/V2/A3/c1 ));
 AND2_X1 \V1/V2/V2/A3/M2/M1/_0_  (.A1(\V1/V2/V2/v4 [1]),
    .A2(\V1/V2/V2/s2 [3]),
    .ZN(\V1/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M2/M1/_1_  (.A(\V1/V2/V2/v4 [1]),
    .B(\V1/V2/V2/s2 [3]),
    .Z(\V1/V2/V2/A3/M2/s1 ));
 AND2_X1 \V1/V2/V2/A3/M2/M2/_0_  (.A1(\V1/V2/V2/A3/M2/s1 ),
    .A2(\V1/V2/V2/A3/c1 ),
    .ZN(\V1/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M2/M2/_1_  (.A(\V1/V2/V2/A3/M2/s1 ),
    .B(\V1/V2/V2/A3/c1 ),
    .Z(\V1/V2/v2 [5]));
 OR2_X1 \V1/V2/V2/A3/M2/_0_  (.A1(\V1/V2/V2/A3/M2/c1 ),
    .A2(\V1/V2/V2/A3/M2/c2 ),
    .ZN(\V1/V2/V2/A3/c2 ));
 AND2_X1 \V1/V2/V2/A3/M3/M1/_0_  (.A1(\V1/V2/V2/v4 [2]),
    .A2(\V1/V2/V2/c3 ),
    .ZN(\V1/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M3/M1/_1_  (.A(\V1/V2/V2/v4 [2]),
    .B(\V1/V2/V2/c3 ),
    .Z(\V1/V2/V2/A3/M3/s1 ));
 AND2_X1 \V1/V2/V2/A3/M3/M2/_0_  (.A1(\V1/V2/V2/A3/M3/s1 ),
    .A2(\V1/V2/V2/A3/c2 ),
    .ZN(\V1/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M3/M2/_1_  (.A(\V1/V2/V2/A3/M3/s1 ),
    .B(\V1/V2/V2/A3/c2 ),
    .Z(\V1/V2/v2 [6]));
 OR2_X1 \V1/V2/V2/A3/M3/_0_  (.A1(\V1/V2/V2/A3/M3/c1 ),
    .A2(\V1/V2/V2/A3/M3/c2 ),
    .ZN(\V1/V2/V2/A3/c3 ));
 AND2_X1 \V1/V2/V2/A3/M4/M1/_0_  (.A1(\V1/V2/V2/v4 [3]),
    .A2(net3),
    .ZN(\V1/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V2/A3/M4/M1/_1_  (.A(\V1/V2/V2/v4 [3]),
    .B(net3),
    .Z(\V1/V2/V2/A3/M4/s1 ));
 AND2_X1 \V1/V2/V2/A3/M4/M2/_0_  (.A1(\V1/V2/V2/A3/M4/s1 ),
    .A2(\V1/V2/V2/A3/c3 ),
    .ZN(\V1/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V2/A3/M4/M2/_1_  (.A(\V1/V2/V2/A3/M4/s1 ),
    .B(\V1/V2/V2/A3/c3 ),
    .Z(\V1/V2/v2 [7]));
 OR2_X1 \V1/V2/V2/A3/M4/_0_  (.A1(\V1/V2/V2/A3/M4/c1 ),
    .A2(\V1/V2/V2/A3/M4/c2 ),
    .ZN(\V1/V2/V2/overflow ));
 AND2_X1 \V1/V2/V2/V1/HA1/_0_  (.A1(\V1/V2/V2/V1/w2 ),
    .A2(\V1/V2/V2/V1/w1 ),
    .ZN(\V1/V2/V2/V1/w4 ));
 XOR2_X2 \V1/V2/V2/V1/HA1/_1_  (.A(\V1/V2/V2/V1/w2 ),
    .B(\V1/V2/V2/V1/w1 ),
    .Z(\V1/V2/v2 [1]));
 AND2_X1 \V1/V2/V2/V1/HA2/_0_  (.A1(\V1/V2/V2/V1/w4 ),
    .A2(\V1/V2/V2/V1/w3 ),
    .ZN(\V1/V2/V2/v1 [3]));
 XOR2_X2 \V1/V2/V2/V1/HA2/_1_  (.A(\V1/V2/V2/V1/w4 ),
    .B(\V1/V2/V2/V1/w3 ),
    .Z(\V1/V2/V2/v1 [2]));
 AND2_X1 \V1/V2/V2/V1/_0_  (.A1(net45),
    .A2(B[0]),
    .ZN(\V1/V2/v2 [0]));
 AND2_X1 \V1/V2/V2/V1/_1_  (.A1(net45),
    .A2(B[1]),
    .ZN(\V1/V2/V2/V1/w1 ));
 AND2_X1 \V1/V2/V2/V1/_2_  (.A1(B[0]),
    .A2(net44),
    .ZN(\V1/V2/V2/V1/w2 ));
 AND2_X1 \V1/V2/V2/V1/_3_  (.A1(B[1]),
    .A2(net44),
    .ZN(\V1/V2/V2/V1/w3 ));
 AND2_X1 \V1/V2/V2/V2/HA1/_0_  (.A1(\V1/V2/V2/V2/w2 ),
    .A2(\V1/V2/V2/V2/w1 ),
    .ZN(\V1/V2/V2/V2/w4 ));
 XOR2_X2 \V1/V2/V2/V2/HA1/_1_  (.A(\V1/V2/V2/V2/w2 ),
    .B(\V1/V2/V2/V2/w1 ),
    .Z(\V1/V2/V2/v2 [1]));
 AND2_X1 \V1/V2/V2/V2/HA2/_0_  (.A1(\V1/V2/V2/V2/w4 ),
    .A2(\V1/V2/V2/V2/w3 ),
    .ZN(\V1/V2/V2/v2 [3]));
 XOR2_X2 \V1/V2/V2/V2/HA2/_1_  (.A(\V1/V2/V2/V2/w4 ),
    .B(\V1/V2/V2/V2/w3 ),
    .Z(\V1/V2/V2/v2 [2]));
 AND2_X1 \V1/V2/V2/V2/_0_  (.A1(net43),
    .A2(B[0]),
    .ZN(\V1/V2/V2/v2 [0]));
 AND2_X1 \V1/V2/V2/V2/_1_  (.A1(net43),
    .A2(B[1]),
    .ZN(\V1/V2/V2/V2/w1 ));
 AND2_X1 \V1/V2/V2/V2/_2_  (.A1(B[0]),
    .A2(net42),
    .ZN(\V1/V2/V2/V2/w2 ));
 AND2_X1 \V1/V2/V2/V2/_3_  (.A1(B[1]),
    .A2(net42),
    .ZN(\V1/V2/V2/V2/w3 ));
 AND2_X1 \V1/V2/V2/V3/HA1/_0_  (.A1(\V1/V2/V2/V3/w2 ),
    .A2(\V1/V2/V2/V3/w1 ),
    .ZN(\V1/V2/V2/V3/w4 ));
 XOR2_X2 \V1/V2/V2/V3/HA1/_1_  (.A(\V1/V2/V2/V3/w2 ),
    .B(\V1/V2/V2/V3/w1 ),
    .Z(\V1/V2/V2/v3 [1]));
 AND2_X1 \V1/V2/V2/V3/HA2/_0_  (.A1(\V1/V2/V2/V3/w4 ),
    .A2(\V1/V2/V2/V3/w3 ),
    .ZN(\V1/V2/V2/v3 [3]));
 XOR2_X2 \V1/V2/V2/V3/HA2/_1_  (.A(\V1/V2/V2/V3/w4 ),
    .B(\V1/V2/V2/V3/w3 ),
    .Z(\V1/V2/V2/v3 [2]));
 AND2_X1 \V1/V2/V2/V3/_0_  (.A1(net45),
    .A2(B[2]),
    .ZN(\V1/V2/V2/v3 [0]));
 AND2_X1 \V1/V2/V2/V3/_1_  (.A1(net45),
    .A2(B[3]),
    .ZN(\V1/V2/V2/V3/w1 ));
 AND2_X1 \V1/V2/V2/V3/_2_  (.A1(B[2]),
    .A2(net44),
    .ZN(\V1/V2/V2/V3/w2 ));
 AND2_X1 \V1/V2/V2/V3/_3_  (.A1(B[3]),
    .A2(net44),
    .ZN(\V1/V2/V2/V3/w3 ));
 AND2_X1 \V1/V2/V2/V4/HA1/_0_  (.A1(\V1/V2/V2/V4/w2 ),
    .A2(\V1/V2/V2/V4/w1 ),
    .ZN(\V1/V2/V2/V4/w4 ));
 XOR2_X2 \V1/V2/V2/V4/HA1/_1_  (.A(\V1/V2/V2/V4/w2 ),
    .B(\V1/V2/V2/V4/w1 ),
    .Z(\V1/V2/V2/v4 [1]));
 AND2_X1 \V1/V2/V2/V4/HA2/_0_  (.A1(\V1/V2/V2/V4/w4 ),
    .A2(\V1/V2/V2/V4/w3 ),
    .ZN(\V1/V2/V2/v4 [3]));
 XOR2_X2 \V1/V2/V2/V4/HA2/_1_  (.A(\V1/V2/V2/V4/w4 ),
    .B(\V1/V2/V2/V4/w3 ),
    .Z(\V1/V2/V2/v4 [2]));
 AND2_X1 \V1/V2/V2/V4/_0_  (.A1(net43),
    .A2(B[2]),
    .ZN(\V1/V2/V2/v4 [0]));
 AND2_X1 \V1/V2/V2/V4/_1_  (.A1(net43),
    .A2(B[3]),
    .ZN(\V1/V2/V2/V4/w1 ));
 AND2_X1 \V1/V2/V2/V4/_2_  (.A1(B[2]),
    .A2(net42),
    .ZN(\V1/V2/V2/V4/w2 ));
 AND2_X1 \V1/V2/V2/V4/_3_  (.A1(B[3]),
    .A2(net42),
    .ZN(\V1/V2/V2/V4/w3 ));
 OR2_X1 \V1/V2/V2/_0_  (.A1(\V1/V2/V2/c1 ),
    .A2(\V1/V2/V2/c2 ),
    .ZN(\V1/V2/V2/c3 ));
 AND2_X1 \V1/V2/V3/A1/M1/M1/_0_  (.A1(\V1/V2/V3/v2 [0]),
    .A2(\V1/V2/V3/v3 [0]),
    .ZN(\V1/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M1/M1/_1_  (.A(\V1/V2/V3/v2 [0]),
    .B(\V1/V2/V3/v3 [0]),
    .Z(\V1/V2/V3/A1/M1/s1 ));
 AND2_X1 \V1/V2/V3/A1/M1/M2/_0_  (.A1(\V1/V2/V3/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M1/M2/_1_  (.A(\V1/V2/V3/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/V3/s1 [0]));
 OR2_X1 \V1/V2/V3/A1/M1/_0_  (.A1(\V1/V2/V3/A1/M1/c1 ),
    .A2(\V1/V2/V3/A1/M1/c2 ),
    .ZN(\V1/V2/V3/A1/c1 ));
 AND2_X1 \V1/V2/V3/A1/M2/M1/_0_  (.A1(\V1/V2/V3/v2 [1]),
    .A2(\V1/V2/V3/v3 [1]),
    .ZN(\V1/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M2/M1/_1_  (.A(\V1/V2/V3/v2 [1]),
    .B(\V1/V2/V3/v3 [1]),
    .Z(\V1/V2/V3/A1/M2/s1 ));
 AND2_X1 \V1/V2/V3/A1/M2/M2/_0_  (.A1(\V1/V2/V3/A1/M2/s1 ),
    .A2(\V1/V2/V3/A1/c1 ),
    .ZN(\V1/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M2/M2/_1_  (.A(\V1/V2/V3/A1/M2/s1 ),
    .B(\V1/V2/V3/A1/c1 ),
    .Z(\V1/V2/V3/s1 [1]));
 OR2_X1 \V1/V2/V3/A1/M2/_0_  (.A1(\V1/V2/V3/A1/M2/c1 ),
    .A2(\V1/V2/V3/A1/M2/c2 ),
    .ZN(\V1/V2/V3/A1/c2 ));
 AND2_X1 \V1/V2/V3/A1/M3/M1/_0_  (.A1(\V1/V2/V3/v2 [2]),
    .A2(\V1/V2/V3/v3 [2]),
    .ZN(\V1/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M3/M1/_1_  (.A(\V1/V2/V3/v2 [2]),
    .B(\V1/V2/V3/v3 [2]),
    .Z(\V1/V2/V3/A1/M3/s1 ));
 AND2_X1 \V1/V2/V3/A1/M3/M2/_0_  (.A1(\V1/V2/V3/A1/M3/s1 ),
    .A2(\V1/V2/V3/A1/c2 ),
    .ZN(\V1/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M3/M2/_1_  (.A(\V1/V2/V3/A1/M3/s1 ),
    .B(\V1/V2/V3/A1/c2 ),
    .Z(\V1/V2/V3/s1 [2]));
 OR2_X1 \V1/V2/V3/A1/M3/_0_  (.A1(\V1/V2/V3/A1/M3/c1 ),
    .A2(\V1/V2/V3/A1/M3/c2 ),
    .ZN(\V1/V2/V3/A1/c3 ));
 AND2_X1 \V1/V2/V3/A1/M4/M1/_0_  (.A1(\V1/V2/V3/v2 [3]),
    .A2(\V1/V2/V3/v3 [3]),
    .ZN(\V1/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A1/M4/M1/_1_  (.A(\V1/V2/V3/v2 [3]),
    .B(\V1/V2/V3/v3 [3]),
    .Z(\V1/V2/V3/A1/M4/s1 ));
 AND2_X1 \V1/V2/V3/A1/M4/M2/_0_  (.A1(\V1/V2/V3/A1/M4/s1 ),
    .A2(\V1/V2/V3/A1/c3 ),
    .ZN(\V1/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A1/M4/M2/_1_  (.A(\V1/V2/V3/A1/M4/s1 ),
    .B(\V1/V2/V3/A1/c3 ),
    .Z(\V1/V2/V3/s1 [3]));
 OR2_X1 \V1/V2/V3/A1/M4/_0_  (.A1(\V1/V2/V3/A1/M4/c1 ),
    .A2(\V1/V2/V3/A1/M4/c2 ),
    .ZN(\V1/V2/V3/c1 ));
 AND2_X1 \V1/V2/V3/A2/M1/M1/_0_  (.A1(\V1/V2/V3/s1 [0]),
    .A2(\V1/V2/V3/v1 [2]),
    .ZN(\V1/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M1/M1/_1_  (.A(\V1/V2/V3/s1 [0]),
    .B(\V1/V2/V3/v1 [2]),
    .Z(\V1/V2/V3/A2/M1/s1 ));
 AND2_X1 \V1/V2/V3/A2/M1/M2/_0_  (.A1(\V1/V2/V3/A2/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M1/M2/_1_  (.A(\V1/V2/V3/A2/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v3 [2]));
 OR2_X1 \V1/V2/V3/A2/M1/_0_  (.A1(\V1/V2/V3/A2/M1/c1 ),
    .A2(\V1/V2/V3/A2/M1/c2 ),
    .ZN(\V1/V2/V3/A2/c1 ));
 AND2_X1 \V1/V2/V3/A2/M2/M1/_0_  (.A1(\V1/V2/V3/s1 [1]),
    .A2(\V1/V2/V3/v1 [3]),
    .ZN(\V1/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M2/M1/_1_  (.A(\V1/V2/V3/s1 [1]),
    .B(\V1/V2/V3/v1 [3]),
    .Z(\V1/V2/V3/A2/M2/s1 ));
 AND2_X1 \V1/V2/V3/A2/M2/M2/_0_  (.A1(\V1/V2/V3/A2/M2/s1 ),
    .A2(\V1/V2/V3/A2/c1 ),
    .ZN(\V1/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M2/M2/_1_  (.A(\V1/V2/V3/A2/M2/s1 ),
    .B(\V1/V2/V3/A2/c1 ),
    .Z(\V1/V2/v3 [3]));
 OR2_X1 \V1/V2/V3/A2/M2/_0_  (.A1(\V1/V2/V3/A2/M2/c1 ),
    .A2(\V1/V2/V3/A2/M2/c2 ),
    .ZN(\V1/V2/V3/A2/c2 ));
 AND2_X1 \V1/V2/V3/A2/M3/M1/_0_  (.A1(\V1/V2/V3/s1 [2]),
    .A2(net3),
    .ZN(\V1/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M3/M1/_1_  (.A(\V1/V2/V3/s1 [2]),
    .B(net3),
    .Z(\V1/V2/V3/A2/M3/s1 ));
 AND2_X1 \V1/V2/V3/A2/M3/M2/_0_  (.A1(\V1/V2/V3/A2/M3/s1 ),
    .A2(\V1/V2/V3/A2/c2 ),
    .ZN(\V1/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M3/M2/_1_  (.A(\V1/V2/V3/A2/M3/s1 ),
    .B(\V1/V2/V3/A2/c2 ),
    .Z(\V1/V2/V3/s2 [2]));
 OR2_X1 \V1/V2/V3/A2/M3/_0_  (.A1(\V1/V2/V3/A2/M3/c1 ),
    .A2(\V1/V2/V3/A2/M3/c2 ),
    .ZN(\V1/V2/V3/A2/c3 ));
 AND2_X1 \V1/V2/V3/A2/M4/M1/_0_  (.A1(\V1/V2/V3/s1 [3]),
    .A2(net3),
    .ZN(\V1/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A2/M4/M1/_1_  (.A(\V1/V2/V3/s1 [3]),
    .B(net3),
    .Z(\V1/V2/V3/A2/M4/s1 ));
 AND2_X1 \V1/V2/V3/A2/M4/M2/_0_  (.A1(\V1/V2/V3/A2/M4/s1 ),
    .A2(\V1/V2/V3/A2/c3 ),
    .ZN(\V1/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A2/M4/M2/_1_  (.A(\V1/V2/V3/A2/M4/s1 ),
    .B(\V1/V2/V3/A2/c3 ),
    .Z(\V1/V2/V3/s2 [3]));
 OR2_X1 \V1/V2/V3/A2/M4/_0_  (.A1(\V1/V2/V3/A2/M4/c1 ),
    .A2(\V1/V2/V3/A2/M4/c2 ),
    .ZN(\V1/V2/V3/c2 ));
 AND2_X1 \V1/V2/V3/A3/M1/M1/_0_  (.A1(\V1/V2/V3/v4 [0]),
    .A2(\V1/V2/V3/s2 [2]),
    .ZN(\V1/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M1/M1/_1_  (.A(\V1/V2/V3/v4 [0]),
    .B(\V1/V2/V3/s2 [2]),
    .Z(\V1/V2/V3/A3/M1/s1 ));
 AND2_X1 \V1/V2/V3/A3/M1/M2/_0_  (.A1(\V1/V2/V3/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M1/M2/_1_  (.A(\V1/V2/V3/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v3 [4]));
 OR2_X1 \V1/V2/V3/A3/M1/_0_  (.A1(\V1/V2/V3/A3/M1/c1 ),
    .A2(\V1/V2/V3/A3/M1/c2 ),
    .ZN(\V1/V2/V3/A3/c1 ));
 AND2_X1 \V1/V2/V3/A3/M2/M1/_0_  (.A1(\V1/V2/V3/v4 [1]),
    .A2(\V1/V2/V3/s2 [3]),
    .ZN(\V1/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M2/M1/_1_  (.A(\V1/V2/V3/v4 [1]),
    .B(\V1/V2/V3/s2 [3]),
    .Z(\V1/V2/V3/A3/M2/s1 ));
 AND2_X1 \V1/V2/V3/A3/M2/M2/_0_  (.A1(\V1/V2/V3/A3/M2/s1 ),
    .A2(\V1/V2/V3/A3/c1 ),
    .ZN(\V1/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M2/M2/_1_  (.A(\V1/V2/V3/A3/M2/s1 ),
    .B(\V1/V2/V3/A3/c1 ),
    .Z(\V1/V2/v3 [5]));
 OR2_X1 \V1/V2/V3/A3/M2/_0_  (.A1(\V1/V2/V3/A3/M2/c1 ),
    .A2(\V1/V2/V3/A3/M2/c2 ),
    .ZN(\V1/V2/V3/A3/c2 ));
 AND2_X1 \V1/V2/V3/A3/M3/M1/_0_  (.A1(\V1/V2/V3/v4 [2]),
    .A2(\V1/V2/V3/c3 ),
    .ZN(\V1/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M3/M1/_1_  (.A(\V1/V2/V3/v4 [2]),
    .B(\V1/V2/V3/c3 ),
    .Z(\V1/V2/V3/A3/M3/s1 ));
 AND2_X1 \V1/V2/V3/A3/M3/M2/_0_  (.A1(\V1/V2/V3/A3/M3/s1 ),
    .A2(\V1/V2/V3/A3/c2 ),
    .ZN(\V1/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M3/M2/_1_  (.A(\V1/V2/V3/A3/M3/s1 ),
    .B(\V1/V2/V3/A3/c2 ),
    .Z(\V1/V2/v3 [6]));
 OR2_X1 \V1/V2/V3/A3/M3/_0_  (.A1(\V1/V2/V3/A3/M3/c1 ),
    .A2(\V1/V2/V3/A3/M3/c2 ),
    .ZN(\V1/V2/V3/A3/c3 ));
 AND2_X1 \V1/V2/V3/A3/M4/M1/_0_  (.A1(\V1/V2/V3/v4 [3]),
    .A2(net3),
    .ZN(\V1/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V3/A3/M4/M1/_1_  (.A(\V1/V2/V3/v4 [3]),
    .B(net3),
    .Z(\V1/V2/V3/A3/M4/s1 ));
 AND2_X1 \V1/V2/V3/A3/M4/M2/_0_  (.A1(\V1/V2/V3/A3/M4/s1 ),
    .A2(\V1/V2/V3/A3/c3 ),
    .ZN(\V1/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V3/A3/M4/M2/_1_  (.A(\V1/V2/V3/A3/M4/s1 ),
    .B(\V1/V2/V3/A3/c3 ),
    .Z(\V1/V2/v3 [7]));
 OR2_X1 \V1/V2/V3/A3/M4/_0_  (.A1(\V1/V2/V3/A3/M4/c1 ),
    .A2(\V1/V2/V3/A3/M4/c2 ),
    .ZN(\V1/V2/V3/overflow ));
 AND2_X1 \V1/V2/V3/V1/HA1/_0_  (.A1(\V1/V2/V3/V1/w2 ),
    .A2(\V1/V2/V3/V1/w1 ),
    .ZN(\V1/V2/V3/V1/w4 ));
 XOR2_X2 \V1/V2/V3/V1/HA1/_1_  (.A(\V1/V2/V3/V1/w2 ),
    .B(\V1/V2/V3/V1/w1 ),
    .Z(\V1/V2/v3 [1]));
 AND2_X1 \V1/V2/V3/V1/HA2/_0_  (.A1(\V1/V2/V3/V1/w4 ),
    .A2(\V1/V2/V3/V1/w3 ),
    .ZN(\V1/V2/V3/v1 [3]));
 XOR2_X2 \V1/V2/V3/V1/HA2/_1_  (.A(\V1/V2/V3/V1/w4 ),
    .B(\V1/V2/V3/V1/w3 ),
    .Z(\V1/V2/V3/v1 [2]));
 AND2_X1 \V1/V2/V3/V1/_0_  (.A1(net25),
    .A2(B[4]),
    .ZN(\V1/V2/v3 [0]));
 AND2_X1 \V1/V2/V3/V1/_1_  (.A1(net25),
    .A2(B[5]),
    .ZN(\V1/V2/V3/V1/w1 ));
 AND2_X1 \V1/V2/V3/V1/_2_  (.A1(B[4]),
    .A2(net24),
    .ZN(\V1/V2/V3/V1/w2 ));
 AND2_X1 \V1/V2/V3/V1/_3_  (.A1(B[5]),
    .A2(net24),
    .ZN(\V1/V2/V3/V1/w3 ));
 AND2_X1 \V1/V2/V3/V2/HA1/_0_  (.A1(\V1/V2/V3/V2/w2 ),
    .A2(\V1/V2/V3/V2/w1 ),
    .ZN(\V1/V2/V3/V2/w4 ));
 XOR2_X2 \V1/V2/V3/V2/HA1/_1_  (.A(\V1/V2/V3/V2/w2 ),
    .B(\V1/V2/V3/V2/w1 ),
    .Z(\V1/V2/V3/v2 [1]));
 AND2_X1 \V1/V2/V3/V2/HA2/_0_  (.A1(\V1/V2/V3/V2/w4 ),
    .A2(\V1/V2/V3/V2/w3 ),
    .ZN(\V1/V2/V3/v2 [3]));
 XOR2_X2 \V1/V2/V3/V2/HA2/_1_  (.A(\V1/V2/V3/V2/w4 ),
    .B(\V1/V2/V3/V2/w3 ),
    .Z(\V1/V2/V3/v2 [2]));
 AND2_X1 \V1/V2/V3/V2/_0_  (.A1(net47),
    .A2(B[4]),
    .ZN(\V1/V2/V3/v2 [0]));
 AND2_X1 \V1/V2/V3/V2/_1_  (.A1(net47),
    .A2(B[5]),
    .ZN(\V1/V2/V3/V2/w1 ));
 AND2_X1 \V1/V2/V3/V2/_2_  (.A1(B[4]),
    .A2(net46),
    .ZN(\V1/V2/V3/V2/w2 ));
 AND2_X1 \V1/V2/V3/V2/_3_  (.A1(B[5]),
    .A2(net46),
    .ZN(\V1/V2/V3/V2/w3 ));
 AND2_X1 \V1/V2/V3/V3/HA1/_0_  (.A1(\V1/V2/V3/V3/w2 ),
    .A2(\V1/V2/V3/V3/w1 ),
    .ZN(\V1/V2/V3/V3/w4 ));
 XOR2_X2 \V1/V2/V3/V3/HA1/_1_  (.A(\V1/V2/V3/V3/w2 ),
    .B(\V1/V2/V3/V3/w1 ),
    .Z(\V1/V2/V3/v3 [1]));
 AND2_X1 \V1/V2/V3/V3/HA2/_0_  (.A1(\V1/V2/V3/V3/w4 ),
    .A2(\V1/V2/V3/V3/w3 ),
    .ZN(\V1/V2/V3/v3 [3]));
 XOR2_X2 \V1/V2/V3/V3/HA2/_1_  (.A(\V1/V2/V3/V3/w4 ),
    .B(\V1/V2/V3/V3/w3 ),
    .Z(\V1/V2/V3/v3 [2]));
 AND2_X1 \V1/V2/V3/V3/_0_  (.A1(net25),
    .A2(B[6]),
    .ZN(\V1/V2/V3/v3 [0]));
 AND2_X1 \V1/V2/V3/V3/_1_  (.A1(net25),
    .A2(B[7]),
    .ZN(\V1/V2/V3/V3/w1 ));
 AND2_X1 \V1/V2/V3/V3/_2_  (.A1(B[6]),
    .A2(net24),
    .ZN(\V1/V2/V3/V3/w2 ));
 AND2_X1 \V1/V2/V3/V3/_3_  (.A1(B[7]),
    .A2(net24),
    .ZN(\V1/V2/V3/V3/w3 ));
 AND2_X1 \V1/V2/V3/V4/HA1/_0_  (.A1(\V1/V2/V3/V4/w2 ),
    .A2(\V1/V2/V3/V4/w1 ),
    .ZN(\V1/V2/V3/V4/w4 ));
 XOR2_X2 \V1/V2/V3/V4/HA1/_1_  (.A(\V1/V2/V3/V4/w2 ),
    .B(\V1/V2/V3/V4/w1 ),
    .Z(\V1/V2/V3/v4 [1]));
 AND2_X1 \V1/V2/V3/V4/HA2/_0_  (.A1(\V1/V2/V3/V4/w4 ),
    .A2(\V1/V2/V3/V4/w3 ),
    .ZN(\V1/V2/V3/v4 [3]));
 XOR2_X2 \V1/V2/V3/V4/HA2/_1_  (.A(\V1/V2/V3/V4/w4 ),
    .B(\V1/V2/V3/V4/w3 ),
    .Z(\V1/V2/V3/v4 [2]));
 AND2_X1 \V1/V2/V3/V4/_0_  (.A1(net47),
    .A2(B[6]),
    .ZN(\V1/V2/V3/v4 [0]));
 AND2_X1 \V1/V2/V3/V4/_1_  (.A1(net47),
    .A2(B[7]),
    .ZN(\V1/V2/V3/V4/w1 ));
 AND2_X1 \V1/V2/V3/V4/_2_  (.A1(B[6]),
    .A2(net46),
    .ZN(\V1/V2/V3/V4/w2 ));
 AND2_X1 \V1/V2/V3/V4/_3_  (.A1(B[7]),
    .A2(net46),
    .ZN(\V1/V2/V3/V4/w3 ));
 OR2_X1 \V1/V2/V3/_0_  (.A1(\V1/V2/V3/c1 ),
    .A2(\V1/V2/V3/c2 ),
    .ZN(\V1/V2/V3/c3 ));
 AND2_X1 \V1/V2/V4/A1/M1/M1/_0_  (.A1(\V1/V2/V4/v2 [0]),
    .A2(\V1/V2/V4/v3 [0]),
    .ZN(\V1/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M1/M1/_1_  (.A(\V1/V2/V4/v2 [0]),
    .B(\V1/V2/V4/v3 [0]),
    .Z(\V1/V2/V4/A1/M1/s1 ));
 AND2_X1 \V1/V2/V4/A1/M1/M2/_0_  (.A1(\V1/V2/V4/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M1/M2/_1_  (.A(\V1/V2/V4/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/V4/s1 [0]));
 OR2_X1 \V1/V2/V4/A1/M1/_0_  (.A1(\V1/V2/V4/A1/M1/c1 ),
    .A2(\V1/V2/V4/A1/M1/c2 ),
    .ZN(\V1/V2/V4/A1/c1 ));
 AND2_X1 \V1/V2/V4/A1/M2/M1/_0_  (.A1(\V1/V2/V4/v2 [1]),
    .A2(\V1/V2/V4/v3 [1]),
    .ZN(\V1/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M2/M1/_1_  (.A(\V1/V2/V4/v2 [1]),
    .B(\V1/V2/V4/v3 [1]),
    .Z(\V1/V2/V4/A1/M2/s1 ));
 AND2_X1 \V1/V2/V4/A1/M2/M2/_0_  (.A1(\V1/V2/V4/A1/M2/s1 ),
    .A2(\V1/V2/V4/A1/c1 ),
    .ZN(\V1/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M2/M2/_1_  (.A(\V1/V2/V4/A1/M2/s1 ),
    .B(\V1/V2/V4/A1/c1 ),
    .Z(\V1/V2/V4/s1 [1]));
 OR2_X1 \V1/V2/V4/A1/M2/_0_  (.A1(\V1/V2/V4/A1/M2/c1 ),
    .A2(\V1/V2/V4/A1/M2/c2 ),
    .ZN(\V1/V2/V4/A1/c2 ));
 AND2_X1 \V1/V2/V4/A1/M3/M1/_0_  (.A1(\V1/V2/V4/v2 [2]),
    .A2(\V1/V2/V4/v3 [2]),
    .ZN(\V1/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M3/M1/_1_  (.A(\V1/V2/V4/v2 [2]),
    .B(\V1/V2/V4/v3 [2]),
    .Z(\V1/V2/V4/A1/M3/s1 ));
 AND2_X1 \V1/V2/V4/A1/M3/M2/_0_  (.A1(\V1/V2/V4/A1/M3/s1 ),
    .A2(\V1/V2/V4/A1/c2 ),
    .ZN(\V1/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M3/M2/_1_  (.A(\V1/V2/V4/A1/M3/s1 ),
    .B(\V1/V2/V4/A1/c2 ),
    .Z(\V1/V2/V4/s1 [2]));
 OR2_X1 \V1/V2/V4/A1/M3/_0_  (.A1(\V1/V2/V4/A1/M3/c1 ),
    .A2(\V1/V2/V4/A1/M3/c2 ),
    .ZN(\V1/V2/V4/A1/c3 ));
 AND2_X1 \V1/V2/V4/A1/M4/M1/_0_  (.A1(\V1/V2/V4/v2 [3]),
    .A2(\V1/V2/V4/v3 [3]),
    .ZN(\V1/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A1/M4/M1/_1_  (.A(\V1/V2/V4/v2 [3]),
    .B(\V1/V2/V4/v3 [3]),
    .Z(\V1/V2/V4/A1/M4/s1 ));
 AND2_X1 \V1/V2/V4/A1/M4/M2/_0_  (.A1(\V1/V2/V4/A1/M4/s1 ),
    .A2(\V1/V2/V4/A1/c3 ),
    .ZN(\V1/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A1/M4/M2/_1_  (.A(\V1/V2/V4/A1/M4/s1 ),
    .B(\V1/V2/V4/A1/c3 ),
    .Z(\V1/V2/V4/s1 [3]));
 OR2_X1 \V1/V2/V4/A1/M4/_0_  (.A1(\V1/V2/V4/A1/M4/c1 ),
    .A2(\V1/V2/V4/A1/M4/c2 ),
    .ZN(\V1/V2/V4/c1 ));
 AND2_X1 \V1/V2/V4/A2/M1/M1/_0_  (.A1(\V1/V2/V4/s1 [0]),
    .A2(\V1/V2/V4/v1 [2]),
    .ZN(\V1/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M1/M1/_1_  (.A(\V1/V2/V4/s1 [0]),
    .B(\V1/V2/V4/v1 [2]),
    .Z(\V1/V2/V4/A2/M1/s1 ));
 AND2_X1 \V1/V2/V4/A2/M1/M2/_0_  (.A1(\V1/V2/V4/A2/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M1/M2/_1_  (.A(\V1/V2/V4/A2/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v4 [2]));
 OR2_X1 \V1/V2/V4/A2/M1/_0_  (.A1(\V1/V2/V4/A2/M1/c1 ),
    .A2(\V1/V2/V4/A2/M1/c2 ),
    .ZN(\V1/V2/V4/A2/c1 ));
 AND2_X1 \V1/V2/V4/A2/M2/M1/_0_  (.A1(\V1/V2/V4/s1 [1]),
    .A2(\V1/V2/V4/v1 [3]),
    .ZN(\V1/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M2/M1/_1_  (.A(\V1/V2/V4/s1 [1]),
    .B(\V1/V2/V4/v1 [3]),
    .Z(\V1/V2/V4/A2/M2/s1 ));
 AND2_X1 \V1/V2/V4/A2/M2/M2/_0_  (.A1(\V1/V2/V4/A2/M2/s1 ),
    .A2(\V1/V2/V4/A2/c1 ),
    .ZN(\V1/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M2/M2/_1_  (.A(\V1/V2/V4/A2/M2/s1 ),
    .B(\V1/V2/V4/A2/c1 ),
    .Z(\V1/V2/v4 [3]));
 OR2_X1 \V1/V2/V4/A2/M2/_0_  (.A1(\V1/V2/V4/A2/M2/c1 ),
    .A2(\V1/V2/V4/A2/M2/c2 ),
    .ZN(\V1/V2/V4/A2/c2 ));
 AND2_X1 \V1/V2/V4/A2/M3/M1/_0_  (.A1(\V1/V2/V4/s1 [2]),
    .A2(net3),
    .ZN(\V1/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M3/M1/_1_  (.A(\V1/V2/V4/s1 [2]),
    .B(net3),
    .Z(\V1/V2/V4/A2/M3/s1 ));
 AND2_X1 \V1/V2/V4/A2/M3/M2/_0_  (.A1(\V1/V2/V4/A2/M3/s1 ),
    .A2(\V1/V2/V4/A2/c2 ),
    .ZN(\V1/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M3/M2/_1_  (.A(\V1/V2/V4/A2/M3/s1 ),
    .B(\V1/V2/V4/A2/c2 ),
    .Z(\V1/V2/V4/s2 [2]));
 OR2_X1 \V1/V2/V4/A2/M3/_0_  (.A1(\V1/V2/V4/A2/M3/c1 ),
    .A2(\V1/V2/V4/A2/M3/c2 ),
    .ZN(\V1/V2/V4/A2/c3 ));
 AND2_X1 \V1/V2/V4/A2/M4/M1/_0_  (.A1(\V1/V2/V4/s1 [3]),
    .A2(net3),
    .ZN(\V1/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A2/M4/M1/_1_  (.A(\V1/V2/V4/s1 [3]),
    .B(net3),
    .Z(\V1/V2/V4/A2/M4/s1 ));
 AND2_X1 \V1/V2/V4/A2/M4/M2/_0_  (.A1(\V1/V2/V4/A2/M4/s1 ),
    .A2(\V1/V2/V4/A2/c3 ),
    .ZN(\V1/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A2/M4/M2/_1_  (.A(\V1/V2/V4/A2/M4/s1 ),
    .B(\V1/V2/V4/A2/c3 ),
    .Z(\V1/V2/V4/s2 [3]));
 OR2_X1 \V1/V2/V4/A2/M4/_0_  (.A1(\V1/V2/V4/A2/M4/c1 ),
    .A2(\V1/V2/V4/A2/M4/c2 ),
    .ZN(\V1/V2/V4/c2 ));
 AND2_X1 \V1/V2/V4/A3/M1/M1/_0_  (.A1(\V1/V2/V4/v4 [0]),
    .A2(\V1/V2/V4/s2 [2]),
    .ZN(\V1/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M1/M1/_1_  (.A(\V1/V2/V4/v4 [0]),
    .B(\V1/V2/V4/s2 [2]),
    .Z(\V1/V2/V4/A3/M1/s1 ));
 AND2_X1 \V1/V2/V4/A3/M1/M2/_0_  (.A1(\V1/V2/V4/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M1/M2/_1_  (.A(\V1/V2/V4/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V2/v4 [4]));
 OR2_X1 \V1/V2/V4/A3/M1/_0_  (.A1(\V1/V2/V4/A3/M1/c1 ),
    .A2(\V1/V2/V4/A3/M1/c2 ),
    .ZN(\V1/V2/V4/A3/c1 ));
 AND2_X1 \V1/V2/V4/A3/M2/M1/_0_  (.A1(\V1/V2/V4/v4 [1]),
    .A2(\V1/V2/V4/s2 [3]),
    .ZN(\V1/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M2/M1/_1_  (.A(\V1/V2/V4/v4 [1]),
    .B(\V1/V2/V4/s2 [3]),
    .Z(\V1/V2/V4/A3/M2/s1 ));
 AND2_X1 \V1/V2/V4/A3/M2/M2/_0_  (.A1(\V1/V2/V4/A3/M2/s1 ),
    .A2(\V1/V2/V4/A3/c1 ),
    .ZN(\V1/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M2/M2/_1_  (.A(\V1/V2/V4/A3/M2/s1 ),
    .B(\V1/V2/V4/A3/c1 ),
    .Z(\V1/V2/v4 [5]));
 OR2_X1 \V1/V2/V4/A3/M2/_0_  (.A1(\V1/V2/V4/A3/M2/c1 ),
    .A2(\V1/V2/V4/A3/M2/c2 ),
    .ZN(\V1/V2/V4/A3/c2 ));
 AND2_X1 \V1/V2/V4/A3/M3/M1/_0_  (.A1(\V1/V2/V4/v4 [2]),
    .A2(\V1/V2/V4/c3 ),
    .ZN(\V1/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M3/M1/_1_  (.A(\V1/V2/V4/v4 [2]),
    .B(\V1/V2/V4/c3 ),
    .Z(\V1/V2/V4/A3/M3/s1 ));
 AND2_X1 \V1/V2/V4/A3/M3/M2/_0_  (.A1(\V1/V2/V4/A3/M3/s1 ),
    .A2(\V1/V2/V4/A3/c2 ),
    .ZN(\V1/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M3/M2/_1_  (.A(\V1/V2/V4/A3/M3/s1 ),
    .B(\V1/V2/V4/A3/c2 ),
    .Z(\V1/V2/v4 [6]));
 OR2_X1 \V1/V2/V4/A3/M3/_0_  (.A1(\V1/V2/V4/A3/M3/c1 ),
    .A2(\V1/V2/V4/A3/M3/c2 ),
    .ZN(\V1/V2/V4/A3/c3 ));
 AND2_X1 \V1/V2/V4/A3/M4/M1/_0_  (.A1(\V1/V2/V4/v4 [3]),
    .A2(net3),
    .ZN(\V1/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V2/V4/A3/M4/M1/_1_  (.A(\V1/V2/V4/v4 [3]),
    .B(net3),
    .Z(\V1/V2/V4/A3/M4/s1 ));
 AND2_X1 \V1/V2/V4/A3/M4/M2/_0_  (.A1(\V1/V2/V4/A3/M4/s1 ),
    .A2(\V1/V2/V4/A3/c3 ),
    .ZN(\V1/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V2/V4/A3/M4/M2/_1_  (.A(\V1/V2/V4/A3/M4/s1 ),
    .B(\V1/V2/V4/A3/c3 ),
    .Z(\V1/V2/v4 [7]));
 OR2_X1 \V1/V2/V4/A3/M4/_0_  (.A1(\V1/V2/V4/A3/M4/c1 ),
    .A2(\V1/V2/V4/A3/M4/c2 ),
    .ZN(\V1/V2/V4/overflow ));
 AND2_X1 \V1/V2/V4/V1/HA1/_0_  (.A1(\V1/V2/V4/V1/w2 ),
    .A2(\V1/V2/V4/V1/w1 ),
    .ZN(\V1/V2/V4/V1/w4 ));
 XOR2_X2 \V1/V2/V4/V1/HA1/_1_  (.A(\V1/V2/V4/V1/w2 ),
    .B(\V1/V2/V4/V1/w1 ),
    .Z(\V1/V2/v4 [1]));
 AND2_X1 \V1/V2/V4/V1/HA2/_0_  (.A1(\V1/V2/V4/V1/w4 ),
    .A2(\V1/V2/V4/V1/w3 ),
    .ZN(\V1/V2/V4/v1 [3]));
 XOR2_X2 \V1/V2/V4/V1/HA2/_1_  (.A(\V1/V2/V4/V1/w4 ),
    .B(\V1/V2/V4/V1/w3 ),
    .Z(\V1/V2/V4/v1 [2]));
 AND2_X1 \V1/V2/V4/V1/_0_  (.A1(net45),
    .A2(B[4]),
    .ZN(\V1/V2/v4 [0]));
 AND2_X1 \V1/V2/V4/V1/_1_  (.A1(net45),
    .A2(B[5]),
    .ZN(\V1/V2/V4/V1/w1 ));
 AND2_X1 \V1/V2/V4/V1/_2_  (.A1(B[4]),
    .A2(net44),
    .ZN(\V1/V2/V4/V1/w2 ));
 AND2_X1 \V1/V2/V4/V1/_3_  (.A1(B[5]),
    .A2(net44),
    .ZN(\V1/V2/V4/V1/w3 ));
 AND2_X1 \V1/V2/V4/V2/HA1/_0_  (.A1(\V1/V2/V4/V2/w2 ),
    .A2(\V1/V2/V4/V2/w1 ),
    .ZN(\V1/V2/V4/V2/w4 ));
 XOR2_X2 \V1/V2/V4/V2/HA1/_1_  (.A(\V1/V2/V4/V2/w2 ),
    .B(\V1/V2/V4/V2/w1 ),
    .Z(\V1/V2/V4/v2 [1]));
 AND2_X1 \V1/V2/V4/V2/HA2/_0_  (.A1(\V1/V2/V4/V2/w4 ),
    .A2(\V1/V2/V4/V2/w3 ),
    .ZN(\V1/V2/V4/v2 [3]));
 XOR2_X2 \V1/V2/V4/V2/HA2/_1_  (.A(\V1/V2/V4/V2/w4 ),
    .B(\V1/V2/V4/V2/w3 ),
    .Z(\V1/V2/V4/v2 [2]));
 AND2_X1 \V1/V2/V4/V2/_0_  (.A1(net43),
    .A2(B[4]),
    .ZN(\V1/V2/V4/v2 [0]));
 AND2_X1 \V1/V2/V4/V2/_1_  (.A1(net43),
    .A2(B[5]),
    .ZN(\V1/V2/V4/V2/w1 ));
 AND2_X1 \V1/V2/V4/V2/_2_  (.A1(B[4]),
    .A2(net42),
    .ZN(\V1/V2/V4/V2/w2 ));
 AND2_X1 \V1/V2/V4/V2/_3_  (.A1(B[5]),
    .A2(net42),
    .ZN(\V1/V2/V4/V2/w3 ));
 AND2_X1 \V1/V2/V4/V3/HA1/_0_  (.A1(\V1/V2/V4/V3/w2 ),
    .A2(\V1/V2/V4/V3/w1 ),
    .ZN(\V1/V2/V4/V3/w4 ));
 XOR2_X2 \V1/V2/V4/V3/HA1/_1_  (.A(\V1/V2/V4/V3/w2 ),
    .B(\V1/V2/V4/V3/w1 ),
    .Z(\V1/V2/V4/v3 [1]));
 AND2_X1 \V1/V2/V4/V3/HA2/_0_  (.A1(\V1/V2/V4/V3/w4 ),
    .A2(\V1/V2/V4/V3/w3 ),
    .ZN(\V1/V2/V4/v3 [3]));
 XOR2_X2 \V1/V2/V4/V3/HA2/_1_  (.A(\V1/V2/V4/V3/w4 ),
    .B(\V1/V2/V4/V3/w3 ),
    .Z(\V1/V2/V4/v3 [2]));
 AND2_X1 \V1/V2/V4/V3/_0_  (.A1(net45),
    .A2(B[6]),
    .ZN(\V1/V2/V4/v3 [0]));
 AND2_X1 \V1/V2/V4/V3/_1_  (.A1(net45),
    .A2(B[7]),
    .ZN(\V1/V2/V4/V3/w1 ));
 AND2_X1 \V1/V2/V4/V3/_2_  (.A1(B[6]),
    .A2(net44),
    .ZN(\V1/V2/V4/V3/w2 ));
 AND2_X1 \V1/V2/V4/V3/_3_  (.A1(B[7]),
    .A2(net44),
    .ZN(\V1/V2/V4/V3/w3 ));
 AND2_X1 \V1/V2/V4/V4/HA1/_0_  (.A1(\V1/V2/V4/V4/w2 ),
    .A2(\V1/V2/V4/V4/w1 ),
    .ZN(\V1/V2/V4/V4/w4 ));
 XOR2_X2 \V1/V2/V4/V4/HA1/_1_  (.A(\V1/V2/V4/V4/w2 ),
    .B(\V1/V2/V4/V4/w1 ),
    .Z(\V1/V2/V4/v4 [1]));
 AND2_X1 \V1/V2/V4/V4/HA2/_0_  (.A1(\V1/V2/V4/V4/w4 ),
    .A2(\V1/V2/V4/V4/w3 ),
    .ZN(\V1/V2/V4/v4 [3]));
 XOR2_X2 \V1/V2/V4/V4/HA2/_1_  (.A(\V1/V2/V4/V4/w4 ),
    .B(\V1/V2/V4/V4/w3 ),
    .Z(\V1/V2/V4/v4 [2]));
 AND2_X1 \V1/V2/V4/V4/_0_  (.A1(net43),
    .A2(B[6]),
    .ZN(\V1/V2/V4/v4 [0]));
 AND2_X1 \V1/V2/V4/V4/_1_  (.A1(net43),
    .A2(B[7]),
    .ZN(\V1/V2/V4/V4/w1 ));
 AND2_X1 \V1/V2/V4/V4/_2_  (.A1(B[6]),
    .A2(net42),
    .ZN(\V1/V2/V4/V4/w2 ));
 AND2_X1 \V1/V2/V4/V4/_3_  (.A1(B[7]),
    .A2(net42),
    .ZN(\V1/V2/V4/V4/w3 ));
 OR2_X1 \V1/V2/V4/_0_  (.A1(\V1/V2/V4/c1 ),
    .A2(\V1/V2/V4/c2 ),
    .ZN(\V1/V2/V4/c3 ));
 OR2_X1 \V1/V2/_0_  (.A1(\V1/V2/c1 ),
    .A2(\V1/V2/c2 ),
    .ZN(\V1/V2/c3 ));
 AND2_X1 \V1/V3/A1/A1/M1/M1/_0_  (.A1(\V1/V3/v2 [0]),
    .A2(\V1/V3/v3 [0]),
    .ZN(\V1/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M1/M1/_1_  (.A(\V1/V3/v2 [0]),
    .B(\V1/V3/v3 [0]),
    .Z(\V1/V3/A1/A1/M1/s1 ));
 AND2_X1 \V1/V3/A1/A1/M1/M2/_0_  (.A1(\V1/V3/A1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M1/M2/_1_  (.A(\V1/V3/A1/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V3/s1 [0]));
 OR2_X1 \V1/V3/A1/A1/M1/_0_  (.A1(\V1/V3/A1/A1/M1/c1 ),
    .A2(\V1/V3/A1/A1/M1/c2 ),
    .ZN(\V1/V3/A1/A1/c1 ));
 AND2_X1 \V1/V3/A1/A1/M2/M1/_0_  (.A1(\V1/V3/v2 [1]),
    .A2(\V1/V3/v3 [1]),
    .ZN(\V1/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M2/M1/_1_  (.A(\V1/V3/v2 [1]),
    .B(\V1/V3/v3 [1]),
    .Z(\V1/V3/A1/A1/M2/s1 ));
 AND2_X1 \V1/V3/A1/A1/M2/M2/_0_  (.A1(\V1/V3/A1/A1/M2/s1 ),
    .A2(\V1/V3/A1/A1/c1 ),
    .ZN(\V1/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M2/M2/_1_  (.A(\V1/V3/A1/A1/M2/s1 ),
    .B(\V1/V3/A1/A1/c1 ),
    .Z(\V1/V3/s1 [1]));
 OR2_X1 \V1/V3/A1/A1/M2/_0_  (.A1(\V1/V3/A1/A1/M2/c1 ),
    .A2(\V1/V3/A1/A1/M2/c2 ),
    .ZN(\V1/V3/A1/A1/c2 ));
 AND2_X1 \V1/V3/A1/A1/M3/M1/_0_  (.A1(\V1/V3/v2 [2]),
    .A2(\V1/V3/v3 [2]),
    .ZN(\V1/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M3/M1/_1_  (.A(\V1/V3/v2 [2]),
    .B(\V1/V3/v3 [2]),
    .Z(\V1/V3/A1/A1/M3/s1 ));
 AND2_X1 \V1/V3/A1/A1/M3/M2/_0_  (.A1(\V1/V3/A1/A1/M3/s1 ),
    .A2(\V1/V3/A1/A1/c2 ),
    .ZN(\V1/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M3/M2/_1_  (.A(\V1/V3/A1/A1/M3/s1 ),
    .B(\V1/V3/A1/A1/c2 ),
    .Z(\V1/V3/s1 [2]));
 OR2_X1 \V1/V3/A1/A1/M3/_0_  (.A1(\V1/V3/A1/A1/M3/c1 ),
    .A2(\V1/V3/A1/A1/M3/c2 ),
    .ZN(\V1/V3/A1/A1/c3 ));
 AND2_X1 \V1/V3/A1/A1/M4/M1/_0_  (.A1(\V1/V3/v2 [3]),
    .A2(\V1/V3/v3 [3]),
    .ZN(\V1/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A1/A1/M4/M1/_1_  (.A(\V1/V3/v2 [3]),
    .B(\V1/V3/v3 [3]),
    .Z(\V1/V3/A1/A1/M4/s1 ));
 AND2_X1 \V1/V3/A1/A1/M4/M2/_0_  (.A1(\V1/V3/A1/A1/M4/s1 ),
    .A2(\V1/V3/A1/A1/c3 ),
    .ZN(\V1/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A1/A1/M4/M2/_1_  (.A(\V1/V3/A1/A1/M4/s1 ),
    .B(\V1/V3/A1/A1/c3 ),
    .Z(\V1/V3/s1 [3]));
 OR2_X1 \V1/V3/A1/A1/M4/_0_  (.A1(\V1/V3/A1/A1/M4/c1 ),
    .A2(\V1/V3/A1/A1/M4/c2 ),
    .ZN(\V1/V3/A1/c1 ));
 AND2_X1 \V1/V3/A1/A2/M1/M1/_0_  (.A1(\V1/V3/v2 [4]),
    .A2(\V1/V3/v3 [4]),
    .ZN(\V1/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M1/M1/_1_  (.A(\V1/V3/v2 [4]),
    .B(\V1/V3/v3 [4]),
    .Z(\V1/V3/A1/A2/M1/s1 ));
 AND2_X1 \V1/V3/A1/A2/M1/M2/_0_  (.A1(\V1/V3/A1/A2/M1/s1 ),
    .A2(\V1/V3/A1/c1 ),
    .ZN(\V1/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M1/M2/_1_  (.A(\V1/V3/A1/A2/M1/s1 ),
    .B(\V1/V3/A1/c1 ),
    .Z(\V1/V3/s1 [4]));
 OR2_X1 \V1/V3/A1/A2/M1/_0_  (.A1(\V1/V3/A1/A2/M1/c1 ),
    .A2(\V1/V3/A1/A2/M1/c2 ),
    .ZN(\V1/V3/A1/A2/c1 ));
 AND2_X1 \V1/V3/A1/A2/M2/M1/_0_  (.A1(\V1/V3/v2 [5]),
    .A2(\V1/V3/v3 [5]),
    .ZN(\V1/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M2/M1/_1_  (.A(\V1/V3/v2 [5]),
    .B(\V1/V3/v3 [5]),
    .Z(\V1/V3/A1/A2/M2/s1 ));
 AND2_X1 \V1/V3/A1/A2/M2/M2/_0_  (.A1(\V1/V3/A1/A2/M2/s1 ),
    .A2(\V1/V3/A1/A2/c1 ),
    .ZN(\V1/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M2/M2/_1_  (.A(\V1/V3/A1/A2/M2/s1 ),
    .B(\V1/V3/A1/A2/c1 ),
    .Z(\V1/V3/s1 [5]));
 OR2_X1 \V1/V3/A1/A2/M2/_0_  (.A1(\V1/V3/A1/A2/M2/c1 ),
    .A2(\V1/V3/A1/A2/M2/c2 ),
    .ZN(\V1/V3/A1/A2/c2 ));
 AND2_X1 \V1/V3/A1/A2/M3/M1/_0_  (.A1(\V1/V3/v2 [6]),
    .A2(\V1/V3/v3 [6]),
    .ZN(\V1/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M3/M1/_1_  (.A(\V1/V3/v2 [6]),
    .B(\V1/V3/v3 [6]),
    .Z(\V1/V3/A1/A2/M3/s1 ));
 AND2_X1 \V1/V3/A1/A2/M3/M2/_0_  (.A1(\V1/V3/A1/A2/M3/s1 ),
    .A2(\V1/V3/A1/A2/c2 ),
    .ZN(\V1/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M3/M2/_1_  (.A(\V1/V3/A1/A2/M3/s1 ),
    .B(\V1/V3/A1/A2/c2 ),
    .Z(\V1/V3/s1 [6]));
 OR2_X1 \V1/V3/A1/A2/M3/_0_  (.A1(\V1/V3/A1/A2/M3/c1 ),
    .A2(\V1/V3/A1/A2/M3/c2 ),
    .ZN(\V1/V3/A1/A2/c3 ));
 AND2_X1 \V1/V3/A1/A2/M4/M1/_0_  (.A1(\V1/V3/v2 [7]),
    .A2(\V1/V3/v3 [7]),
    .ZN(\V1/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A1/A2/M4/M1/_1_  (.A(\V1/V3/v2 [7]),
    .B(\V1/V3/v3 [7]),
    .Z(\V1/V3/A1/A2/M4/s1 ));
 AND2_X1 \V1/V3/A1/A2/M4/M2/_0_  (.A1(\V1/V3/A1/A2/M4/s1 ),
    .A2(\V1/V3/A1/A2/c3 ),
    .ZN(\V1/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A1/A2/M4/M2/_1_  (.A(\V1/V3/A1/A2/M4/s1 ),
    .B(\V1/V3/A1/A2/c3 ),
    .Z(\V1/V3/s1 [7]));
 OR2_X1 \V1/V3/A1/A2/M4/_0_  (.A1(\V1/V3/A1/A2/M4/c1 ),
    .A2(\V1/V3/A1/A2/M4/c2 ),
    .ZN(\V1/V3/c1 ));
 AND2_X1 \V1/V3/A2/A1/M1/M1/_0_  (.A1(\V1/V3/s1 [0]),
    .A2(\V1/V3/v1 [4]),
    .ZN(\V1/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M1/M1/_1_  (.A(\V1/V3/s1 [0]),
    .B(\V1/V3/v1 [4]),
    .Z(\V1/V3/A2/A1/M1/s1 ));
 AND2_X1 \V1/V3/A2/A1/M1/M2/_0_  (.A1(\V1/V3/A2/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M1/M2/_1_  (.A(\V1/V3/A2/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/v3 [4]));
 OR2_X1 \V1/V3/A2/A1/M1/_0_  (.A1(\V1/V3/A2/A1/M1/c1 ),
    .A2(\V1/V3/A2/A1/M1/c2 ),
    .ZN(\V1/V3/A2/A1/c1 ));
 AND2_X1 \V1/V3/A2/A1/M2/M1/_0_  (.A1(\V1/V3/s1 [1]),
    .A2(\V1/V3/v1 [5]),
    .ZN(\V1/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M2/M1/_1_  (.A(\V1/V3/s1 [1]),
    .B(\V1/V3/v1 [5]),
    .Z(\V1/V3/A2/A1/M2/s1 ));
 AND2_X1 \V1/V3/A2/A1/M2/M2/_0_  (.A1(\V1/V3/A2/A1/M2/s1 ),
    .A2(\V1/V3/A2/A1/c1 ),
    .ZN(\V1/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M2/M2/_1_  (.A(\V1/V3/A2/A1/M2/s1 ),
    .B(\V1/V3/A2/A1/c1 ),
    .Z(\V1/v3 [5]));
 OR2_X1 \V1/V3/A2/A1/M2/_0_  (.A1(\V1/V3/A2/A1/M2/c1 ),
    .A2(\V1/V3/A2/A1/M2/c2 ),
    .ZN(\V1/V3/A2/A1/c2 ));
 AND2_X1 \V1/V3/A2/A1/M3/M1/_0_  (.A1(\V1/V3/s1 [2]),
    .A2(\V1/V3/v1 [6]),
    .ZN(\V1/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M3/M1/_1_  (.A(\V1/V3/s1 [2]),
    .B(\V1/V3/v1 [6]),
    .Z(\V1/V3/A2/A1/M3/s1 ));
 AND2_X1 \V1/V3/A2/A1/M3/M2/_0_  (.A1(\V1/V3/A2/A1/M3/s1 ),
    .A2(\V1/V3/A2/A1/c2 ),
    .ZN(\V1/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M3/M2/_1_  (.A(\V1/V3/A2/A1/M3/s1 ),
    .B(\V1/V3/A2/A1/c2 ),
    .Z(\V1/v3 [6]));
 OR2_X1 \V1/V3/A2/A1/M3/_0_  (.A1(\V1/V3/A2/A1/M3/c1 ),
    .A2(\V1/V3/A2/A1/M3/c2 ),
    .ZN(\V1/V3/A2/A1/c3 ));
 AND2_X1 \V1/V3/A2/A1/M4/M1/_0_  (.A1(\V1/V3/s1 [3]),
    .A2(\V1/V3/v1 [7]),
    .ZN(\V1/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A2/A1/M4/M1/_1_  (.A(\V1/V3/s1 [3]),
    .B(\V1/V3/v1 [7]),
    .Z(\V1/V3/A2/A1/M4/s1 ));
 AND2_X1 \V1/V3/A2/A1/M4/M2/_0_  (.A1(\V1/V3/A2/A1/M4/s1 ),
    .A2(\V1/V3/A2/A1/c3 ),
    .ZN(\V1/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A2/A1/M4/M2/_1_  (.A(\V1/V3/A2/A1/M4/s1 ),
    .B(\V1/V3/A2/A1/c3 ),
    .Z(\V1/v3 [7]));
 OR2_X1 \V1/V3/A2/A1/M4/_0_  (.A1(\V1/V3/A2/A1/M4/c1 ),
    .A2(\V1/V3/A2/A1/M4/c2 ),
    .ZN(\V1/V3/A2/c1 ));
 AND2_X1 \V1/V3/A2/A2/M1/M1/_0_  (.A1(\V1/V3/s1 [4]),
    .A2(net3),
    .ZN(\V1/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M1/M1/_1_  (.A(\V1/V3/s1 [4]),
    .B(net3),
    .Z(\V1/V3/A2/A2/M1/s1 ));
 AND2_X1 \V1/V3/A2/A2/M1/M2/_0_  (.A1(\V1/V3/A2/A2/M1/s1 ),
    .A2(\V1/V3/A2/c1 ),
    .ZN(\V1/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M1/M2/_1_  (.A(\V1/V3/A2/A2/M1/s1 ),
    .B(\V1/V3/A2/c1 ),
    .Z(\V1/V3/s2 [4]));
 OR2_X1 \V1/V3/A2/A2/M1/_0_  (.A1(\V1/V3/A2/A2/M1/c1 ),
    .A2(\V1/V3/A2/A2/M1/c2 ),
    .ZN(\V1/V3/A2/A2/c1 ));
 AND2_X1 \V1/V3/A2/A2/M2/M1/_0_  (.A1(\V1/V3/s1 [5]),
    .A2(net3),
    .ZN(\V1/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M2/M1/_1_  (.A(\V1/V3/s1 [5]),
    .B(net3),
    .Z(\V1/V3/A2/A2/M2/s1 ));
 AND2_X1 \V1/V3/A2/A2/M2/M2/_0_  (.A1(\V1/V3/A2/A2/M2/s1 ),
    .A2(\V1/V3/A2/A2/c1 ),
    .ZN(\V1/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M2/M2/_1_  (.A(\V1/V3/A2/A2/M2/s1 ),
    .B(\V1/V3/A2/A2/c1 ),
    .Z(\V1/V3/s2 [5]));
 OR2_X1 \V1/V3/A2/A2/M2/_0_  (.A1(\V1/V3/A2/A2/M2/c1 ),
    .A2(\V1/V3/A2/A2/M2/c2 ),
    .ZN(\V1/V3/A2/A2/c2 ));
 AND2_X1 \V1/V3/A2/A2/M3/M1/_0_  (.A1(\V1/V3/s1 [6]),
    .A2(net3),
    .ZN(\V1/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M3/M1/_1_  (.A(\V1/V3/s1 [6]),
    .B(net3),
    .Z(\V1/V3/A2/A2/M3/s1 ));
 AND2_X1 \V1/V3/A2/A2/M3/M2/_0_  (.A1(\V1/V3/A2/A2/M3/s1 ),
    .A2(\V1/V3/A2/A2/c2 ),
    .ZN(\V1/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M3/M2/_1_  (.A(\V1/V3/A2/A2/M3/s1 ),
    .B(\V1/V3/A2/A2/c2 ),
    .Z(\V1/V3/s2 [6]));
 OR2_X1 \V1/V3/A2/A2/M3/_0_  (.A1(\V1/V3/A2/A2/M3/c1 ),
    .A2(\V1/V3/A2/A2/M3/c2 ),
    .ZN(\V1/V3/A2/A2/c3 ));
 AND2_X1 \V1/V3/A2/A2/M4/M1/_0_  (.A1(\V1/V3/s1 [7]),
    .A2(net3),
    .ZN(\V1/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A2/A2/M4/M1/_1_  (.A(\V1/V3/s1 [7]),
    .B(net3),
    .Z(\V1/V3/A2/A2/M4/s1 ));
 AND2_X1 \V1/V3/A2/A2/M4/M2/_0_  (.A1(\V1/V3/A2/A2/M4/s1 ),
    .A2(\V1/V3/A2/A2/c3 ),
    .ZN(\V1/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A2/A2/M4/M2/_1_  (.A(\V1/V3/A2/A2/M4/s1 ),
    .B(\V1/V3/A2/A2/c3 ),
    .Z(\V1/V3/s2 [7]));
 OR2_X1 \V1/V3/A2/A2/M4/_0_  (.A1(\V1/V3/A2/A2/M4/c1 ),
    .A2(\V1/V3/A2/A2/M4/c2 ),
    .ZN(\V1/V3/c2 ));
 AND2_X1 \V1/V3/A3/A1/M1/M1/_0_  (.A1(\V1/V3/v4 [0]),
    .A2(\V1/V3/s2 [4]),
    .ZN(\V1/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M1/M1/_1_  (.A(\V1/V3/v4 [0]),
    .B(\V1/V3/s2 [4]),
    .Z(\V1/V3/A3/A1/M1/s1 ));
 AND2_X1 \V1/V3/A3/A1/M1/M2/_0_  (.A1(\V1/V3/A3/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M1/M2/_1_  (.A(\V1/V3/A3/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/v3 [8]));
 OR2_X1 \V1/V3/A3/A1/M1/_0_  (.A1(\V1/V3/A3/A1/M1/c1 ),
    .A2(\V1/V3/A3/A1/M1/c2 ),
    .ZN(\V1/V3/A3/A1/c1 ));
 AND2_X1 \V1/V3/A3/A1/M2/M1/_0_  (.A1(\V1/V3/v4 [1]),
    .A2(\V1/V3/s2 [5]),
    .ZN(\V1/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M2/M1/_1_  (.A(\V1/V3/v4 [1]),
    .B(\V1/V3/s2 [5]),
    .Z(\V1/V3/A3/A1/M2/s1 ));
 AND2_X1 \V1/V3/A3/A1/M2/M2/_0_  (.A1(\V1/V3/A3/A1/M2/s1 ),
    .A2(\V1/V3/A3/A1/c1 ),
    .ZN(\V1/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M2/M2/_1_  (.A(\V1/V3/A3/A1/M2/s1 ),
    .B(\V1/V3/A3/A1/c1 ),
    .Z(\V1/v3 [9]));
 OR2_X1 \V1/V3/A3/A1/M2/_0_  (.A1(\V1/V3/A3/A1/M2/c1 ),
    .A2(\V1/V3/A3/A1/M2/c2 ),
    .ZN(\V1/V3/A3/A1/c2 ));
 AND2_X1 \V1/V3/A3/A1/M3/M1/_0_  (.A1(\V1/V3/v4 [2]),
    .A2(\V1/V3/s2 [6]),
    .ZN(\V1/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M3/M1/_1_  (.A(\V1/V3/v4 [2]),
    .B(\V1/V3/s2 [6]),
    .Z(\V1/V3/A3/A1/M3/s1 ));
 AND2_X1 \V1/V3/A3/A1/M3/M2/_0_  (.A1(\V1/V3/A3/A1/M3/s1 ),
    .A2(\V1/V3/A3/A1/c2 ),
    .ZN(\V1/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M3/M2/_1_  (.A(\V1/V3/A3/A1/M3/s1 ),
    .B(\V1/V3/A3/A1/c2 ),
    .Z(\V1/v3 [10]));
 OR2_X1 \V1/V3/A3/A1/M3/_0_  (.A1(\V1/V3/A3/A1/M3/c1 ),
    .A2(\V1/V3/A3/A1/M3/c2 ),
    .ZN(\V1/V3/A3/A1/c3 ));
 AND2_X1 \V1/V3/A3/A1/M4/M1/_0_  (.A1(\V1/V3/v4 [3]),
    .A2(\V1/V3/s2 [7]),
    .ZN(\V1/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V3/A3/A1/M4/M1/_1_  (.A(\V1/V3/v4 [3]),
    .B(\V1/V3/s2 [7]),
    .Z(\V1/V3/A3/A1/M4/s1 ));
 AND2_X1 \V1/V3/A3/A1/M4/M2/_0_  (.A1(\V1/V3/A3/A1/M4/s1 ),
    .A2(\V1/V3/A3/A1/c3 ),
    .ZN(\V1/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V3/A3/A1/M4/M2/_1_  (.A(\V1/V3/A3/A1/M4/s1 ),
    .B(\V1/V3/A3/A1/c3 ),
    .Z(\V1/v3 [11]));
 OR2_X1 \V1/V3/A3/A1/M4/_0_  (.A1(\V1/V3/A3/A1/M4/c1 ),
    .A2(\V1/V3/A3/A1/M4/c2 ),
    .ZN(\V1/V3/A3/c1 ));
 AND2_X1 \V1/V3/A3/A2/M1/M1/_0_  (.A1(\V1/V3/v4 [4]),
    .A2(\V1/V3/c3 ),
    .ZN(\V1/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M1/M1/_1_  (.A(\V1/V3/v4 [4]),
    .B(\V1/V3/c3 ),
    .Z(\V1/V3/A3/A2/M1/s1 ));
 AND2_X1 \V1/V3/A3/A2/M1/M2/_0_  (.A1(\V1/V3/A3/A2/M1/s1 ),
    .A2(\V1/V3/A3/c1 ),
    .ZN(\V1/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M1/M2/_1_  (.A(\V1/V3/A3/A2/M1/s1 ),
    .B(\V1/V3/A3/c1 ),
    .Z(\V1/v3 [12]));
 OR2_X1 \V1/V3/A3/A2/M1/_0_  (.A1(\V1/V3/A3/A2/M1/c1 ),
    .A2(\V1/V3/A3/A2/M1/c2 ),
    .ZN(\V1/V3/A3/A2/c1 ));
 AND2_X1 \V1/V3/A3/A2/M2/M1/_0_  (.A1(\V1/V3/v4 [5]),
    .A2(net3),
    .ZN(\V1/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M2/M1/_1_  (.A(\V1/V3/v4 [5]),
    .B(net3),
    .Z(\V1/V3/A3/A2/M2/s1 ));
 AND2_X1 \V1/V3/A3/A2/M2/M2/_0_  (.A1(\V1/V3/A3/A2/M2/s1 ),
    .A2(\V1/V3/A3/A2/c1 ),
    .ZN(\V1/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M2/M2/_1_  (.A(\V1/V3/A3/A2/M2/s1 ),
    .B(\V1/V3/A3/A2/c1 ),
    .Z(\V1/v3 [13]));
 OR2_X1 \V1/V3/A3/A2/M2/_0_  (.A1(\V1/V3/A3/A2/M2/c1 ),
    .A2(\V1/V3/A3/A2/M2/c2 ),
    .ZN(\V1/V3/A3/A2/c2 ));
 AND2_X1 \V1/V3/A3/A2/M3/M1/_0_  (.A1(\V1/V3/v4 [6]),
    .A2(net3),
    .ZN(\V1/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M3/M1/_1_  (.A(\V1/V3/v4 [6]),
    .B(net3),
    .Z(\V1/V3/A3/A2/M3/s1 ));
 AND2_X1 \V1/V3/A3/A2/M3/M2/_0_  (.A1(\V1/V3/A3/A2/M3/s1 ),
    .A2(\V1/V3/A3/A2/c2 ),
    .ZN(\V1/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M3/M2/_1_  (.A(\V1/V3/A3/A2/M3/s1 ),
    .B(\V1/V3/A3/A2/c2 ),
    .Z(\V1/v3 [14]));
 OR2_X1 \V1/V3/A3/A2/M3/_0_  (.A1(\V1/V3/A3/A2/M3/c1 ),
    .A2(\V1/V3/A3/A2/M3/c2 ),
    .ZN(\V1/V3/A3/A2/c3 ));
 AND2_X1 \V1/V3/A3/A2/M4/M1/_0_  (.A1(\V1/V3/v4 [7]),
    .A2(net3),
    .ZN(\V1/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V3/A3/A2/M4/M1/_1_  (.A(\V1/V3/v4 [7]),
    .B(net3),
    .Z(\V1/V3/A3/A2/M4/s1 ));
 AND2_X1 \V1/V3/A3/A2/M4/M2/_0_  (.A1(\V1/V3/A3/A2/M4/s1 ),
    .A2(\V1/V3/A3/A2/c3 ),
    .ZN(\V1/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V3/A3/A2/M4/M2/_1_  (.A(\V1/V3/A3/A2/M4/s1 ),
    .B(\V1/V3/A3/A2/c3 ),
    .Z(\V1/v3 [15]));
 OR2_X1 \V1/V3/A3/A2/M4/_0_  (.A1(\V1/V3/A3/A2/M4/c1 ),
    .A2(\V1/V3/A3/A2/M4/c2 ),
    .ZN(\V1/V3/overflow ));
 AND2_X1 \V1/V3/V1/A1/M1/M1/_0_  (.A1(\V1/V3/V1/v2 [0]),
    .A2(\V1/V3/V1/v3 [0]),
    .ZN(\V1/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M1/M1/_1_  (.A(\V1/V3/V1/v2 [0]),
    .B(\V1/V3/V1/v3 [0]),
    .Z(\V1/V3/V1/A1/M1/s1 ));
 AND2_X1 \V1/V3/V1/A1/M1/M2/_0_  (.A1(\V1/V3/V1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M1/M2/_1_  (.A(\V1/V3/V1/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V3/V1/s1 [0]));
 OR2_X1 \V1/V3/V1/A1/M1/_0_  (.A1(\V1/V3/V1/A1/M1/c1 ),
    .A2(\V1/V3/V1/A1/M1/c2 ),
    .ZN(\V1/V3/V1/A1/c1 ));
 AND2_X1 \V1/V3/V1/A1/M2/M1/_0_  (.A1(\V1/V3/V1/v2 [1]),
    .A2(\V1/V3/V1/v3 [1]),
    .ZN(\V1/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M2/M1/_1_  (.A(\V1/V3/V1/v2 [1]),
    .B(\V1/V3/V1/v3 [1]),
    .Z(\V1/V3/V1/A1/M2/s1 ));
 AND2_X1 \V1/V3/V1/A1/M2/M2/_0_  (.A1(\V1/V3/V1/A1/M2/s1 ),
    .A2(\V1/V3/V1/A1/c1 ),
    .ZN(\V1/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M2/M2/_1_  (.A(\V1/V3/V1/A1/M2/s1 ),
    .B(\V1/V3/V1/A1/c1 ),
    .Z(\V1/V3/V1/s1 [1]));
 OR2_X1 \V1/V3/V1/A1/M2/_0_  (.A1(\V1/V3/V1/A1/M2/c1 ),
    .A2(\V1/V3/V1/A1/M2/c2 ),
    .ZN(\V1/V3/V1/A1/c2 ));
 AND2_X1 \V1/V3/V1/A1/M3/M1/_0_  (.A1(\V1/V3/V1/v2 [2]),
    .A2(\V1/V3/V1/v3 [2]),
    .ZN(\V1/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M3/M1/_1_  (.A(\V1/V3/V1/v2 [2]),
    .B(\V1/V3/V1/v3 [2]),
    .Z(\V1/V3/V1/A1/M3/s1 ));
 AND2_X1 \V1/V3/V1/A1/M3/M2/_0_  (.A1(\V1/V3/V1/A1/M3/s1 ),
    .A2(\V1/V3/V1/A1/c2 ),
    .ZN(\V1/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M3/M2/_1_  (.A(\V1/V3/V1/A1/M3/s1 ),
    .B(\V1/V3/V1/A1/c2 ),
    .Z(\V1/V3/V1/s1 [2]));
 OR2_X1 \V1/V3/V1/A1/M3/_0_  (.A1(\V1/V3/V1/A1/M3/c1 ),
    .A2(\V1/V3/V1/A1/M3/c2 ),
    .ZN(\V1/V3/V1/A1/c3 ));
 AND2_X1 \V1/V3/V1/A1/M4/M1/_0_  (.A1(\V1/V3/V1/v2 [3]),
    .A2(\V1/V3/V1/v3 [3]),
    .ZN(\V1/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A1/M4/M1/_1_  (.A(\V1/V3/V1/v2 [3]),
    .B(\V1/V3/V1/v3 [3]),
    .Z(\V1/V3/V1/A1/M4/s1 ));
 AND2_X1 \V1/V3/V1/A1/M4/M2/_0_  (.A1(\V1/V3/V1/A1/M4/s1 ),
    .A2(\V1/V3/V1/A1/c3 ),
    .ZN(\V1/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A1/M4/M2/_1_  (.A(\V1/V3/V1/A1/M4/s1 ),
    .B(\V1/V3/V1/A1/c3 ),
    .Z(\V1/V3/V1/s1 [3]));
 OR2_X1 \V1/V3/V1/A1/M4/_0_  (.A1(\V1/V3/V1/A1/M4/c1 ),
    .A2(\V1/V3/V1/A1/M4/c2 ),
    .ZN(\V1/V3/V1/c1 ));
 AND2_X1 \V1/V3/V1/A2/M1/M1/_0_  (.A1(\V1/V3/V1/s1 [0]),
    .A2(\V1/V3/V1/v1 [2]),
    .ZN(\V1/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M1/M1/_1_  (.A(\V1/V3/V1/s1 [0]),
    .B(\V1/V3/V1/v1 [2]),
    .Z(\V1/V3/V1/A2/M1/s1 ));
 AND2_X1 \V1/V3/V1/A2/M1/M2/_0_  (.A1(\V1/V3/V1/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M1/M2/_1_  (.A(\V1/V3/V1/A2/M1/s1 ),
    .B(net4),
    .Z(\V1/v3 [2]));
 OR2_X1 \V1/V3/V1/A2/M1/_0_  (.A1(\V1/V3/V1/A2/M1/c1 ),
    .A2(\V1/V3/V1/A2/M1/c2 ),
    .ZN(\V1/V3/V1/A2/c1 ));
 AND2_X1 \V1/V3/V1/A2/M2/M1/_0_  (.A1(\V1/V3/V1/s1 [1]),
    .A2(\V1/V3/V1/v1 [3]),
    .ZN(\V1/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M2/M1/_1_  (.A(\V1/V3/V1/s1 [1]),
    .B(\V1/V3/V1/v1 [3]),
    .Z(\V1/V3/V1/A2/M2/s1 ));
 AND2_X1 \V1/V3/V1/A2/M2/M2/_0_  (.A1(\V1/V3/V1/A2/M2/s1 ),
    .A2(\V1/V3/V1/A2/c1 ),
    .ZN(\V1/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M2/M2/_1_  (.A(\V1/V3/V1/A2/M2/s1 ),
    .B(\V1/V3/V1/A2/c1 ),
    .Z(\V1/v3 [3]));
 OR2_X1 \V1/V3/V1/A2/M2/_0_  (.A1(\V1/V3/V1/A2/M2/c1 ),
    .A2(\V1/V3/V1/A2/M2/c2 ),
    .ZN(\V1/V3/V1/A2/c2 ));
 AND2_X1 \V1/V3/V1/A2/M3/M1/_0_  (.A1(\V1/V3/V1/s1 [2]),
    .A2(net4),
    .ZN(\V1/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M3/M1/_1_  (.A(\V1/V3/V1/s1 [2]),
    .B(net4),
    .Z(\V1/V3/V1/A2/M3/s1 ));
 AND2_X1 \V1/V3/V1/A2/M3/M2/_0_  (.A1(\V1/V3/V1/A2/M3/s1 ),
    .A2(\V1/V3/V1/A2/c2 ),
    .ZN(\V1/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M3/M2/_1_  (.A(\V1/V3/V1/A2/M3/s1 ),
    .B(\V1/V3/V1/A2/c2 ),
    .Z(\V1/V3/V1/s2 [2]));
 OR2_X1 \V1/V3/V1/A2/M3/_0_  (.A1(\V1/V3/V1/A2/M3/c1 ),
    .A2(\V1/V3/V1/A2/M3/c2 ),
    .ZN(\V1/V3/V1/A2/c3 ));
 AND2_X1 \V1/V3/V1/A2/M4/M1/_0_  (.A1(\V1/V3/V1/s1 [3]),
    .A2(net4),
    .ZN(\V1/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A2/M4/M1/_1_  (.A(\V1/V3/V1/s1 [3]),
    .B(net4),
    .Z(\V1/V3/V1/A2/M4/s1 ));
 AND2_X1 \V1/V3/V1/A2/M4/M2/_0_  (.A1(\V1/V3/V1/A2/M4/s1 ),
    .A2(\V1/V3/V1/A2/c3 ),
    .ZN(\V1/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A2/M4/M2/_1_  (.A(\V1/V3/V1/A2/M4/s1 ),
    .B(\V1/V3/V1/A2/c3 ),
    .Z(\V1/V3/V1/s2 [3]));
 OR2_X1 \V1/V3/V1/A2/M4/_0_  (.A1(\V1/V3/V1/A2/M4/c1 ),
    .A2(\V1/V3/V1/A2/M4/c2 ),
    .ZN(\V1/V3/V1/c2 ));
 AND2_X1 \V1/V3/V1/A3/M1/M1/_0_  (.A1(\V1/V3/V1/v4 [0]),
    .A2(\V1/V3/V1/s2 [2]),
    .ZN(\V1/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M1/M1/_1_  (.A(\V1/V3/V1/v4 [0]),
    .B(\V1/V3/V1/s2 [2]),
    .Z(\V1/V3/V1/A3/M1/s1 ));
 AND2_X1 \V1/V3/V1/A3/M1/M2/_0_  (.A1(\V1/V3/V1/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M1/M2/_1_  (.A(\V1/V3/V1/A3/M1/s1 ),
    .B(net4),
    .Z(\V1/V3/v1 [4]));
 OR2_X1 \V1/V3/V1/A3/M1/_0_  (.A1(\V1/V3/V1/A3/M1/c1 ),
    .A2(\V1/V3/V1/A3/M1/c2 ),
    .ZN(\V1/V3/V1/A3/c1 ));
 AND2_X1 \V1/V3/V1/A3/M2/M1/_0_  (.A1(\V1/V3/V1/v4 [1]),
    .A2(\V1/V3/V1/s2 [3]),
    .ZN(\V1/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M2/M1/_1_  (.A(\V1/V3/V1/v4 [1]),
    .B(\V1/V3/V1/s2 [3]),
    .Z(\V1/V3/V1/A3/M2/s1 ));
 AND2_X1 \V1/V3/V1/A3/M2/M2/_0_  (.A1(\V1/V3/V1/A3/M2/s1 ),
    .A2(\V1/V3/V1/A3/c1 ),
    .ZN(\V1/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M2/M2/_1_  (.A(\V1/V3/V1/A3/M2/s1 ),
    .B(\V1/V3/V1/A3/c1 ),
    .Z(\V1/V3/v1 [5]));
 OR2_X1 \V1/V3/V1/A3/M2/_0_  (.A1(\V1/V3/V1/A3/M2/c1 ),
    .A2(\V1/V3/V1/A3/M2/c2 ),
    .ZN(\V1/V3/V1/A3/c2 ));
 AND2_X1 \V1/V3/V1/A3/M3/M1/_0_  (.A1(\V1/V3/V1/v4 [2]),
    .A2(\V1/V3/V1/c3 ),
    .ZN(\V1/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M3/M1/_1_  (.A(\V1/V3/V1/v4 [2]),
    .B(\V1/V3/V1/c3 ),
    .Z(\V1/V3/V1/A3/M3/s1 ));
 AND2_X1 \V1/V3/V1/A3/M3/M2/_0_  (.A1(\V1/V3/V1/A3/M3/s1 ),
    .A2(\V1/V3/V1/A3/c2 ),
    .ZN(\V1/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M3/M2/_1_  (.A(\V1/V3/V1/A3/M3/s1 ),
    .B(\V1/V3/V1/A3/c2 ),
    .Z(\V1/V3/v1 [6]));
 OR2_X1 \V1/V3/V1/A3/M3/_0_  (.A1(\V1/V3/V1/A3/M3/c1 ),
    .A2(\V1/V3/V1/A3/M3/c2 ),
    .ZN(\V1/V3/V1/A3/c3 ));
 AND2_X1 \V1/V3/V1/A3/M4/M1/_0_  (.A1(\V1/V3/V1/v4 [3]),
    .A2(net5),
    .ZN(\V1/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V1/A3/M4/M1/_1_  (.A(\V1/V3/V1/v4 [3]),
    .B(net5),
    .Z(\V1/V3/V1/A3/M4/s1 ));
 AND2_X1 \V1/V3/V1/A3/M4/M2/_0_  (.A1(\V1/V3/V1/A3/M4/s1 ),
    .A2(\V1/V3/V1/A3/c3 ),
    .ZN(\V1/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V1/A3/M4/M2/_1_  (.A(\V1/V3/V1/A3/M4/s1 ),
    .B(\V1/V3/V1/A3/c3 ),
    .Z(\V1/V3/v1 [7]));
 OR2_X1 \V1/V3/V1/A3/M4/_0_  (.A1(\V1/V3/V1/A3/M4/c1 ),
    .A2(\V1/V3/V1/A3/M4/c2 ),
    .ZN(\V1/V3/V1/overflow ));
 AND2_X1 \V1/V3/V1/V1/HA1/_0_  (.A1(\V1/V3/V1/V1/w2 ),
    .A2(\V1/V3/V1/V1/w1 ),
    .ZN(\V1/V3/V1/V1/w4 ));
 XOR2_X2 \V1/V3/V1/V1/HA1/_1_  (.A(\V1/V3/V1/V1/w2 ),
    .B(\V1/V3/V1/V1/w1 ),
    .Z(\V1/v3 [1]));
 AND2_X1 \V1/V3/V1/V1/HA2/_0_  (.A1(\V1/V3/V1/V1/w4 ),
    .A2(\V1/V3/V1/V1/w3 ),
    .ZN(\V1/V3/V1/v1 [3]));
 XOR2_X2 \V1/V3/V1/V1/HA2/_1_  (.A(\V1/V3/V1/V1/w4 ),
    .B(\V1/V3/V1/V1/w3 ),
    .Z(\V1/V3/V1/v1 [2]));
 AND2_X1 \V1/V3/V1/V1/_0_  (.A1(net48),
    .A2(net12),
    .ZN(\V1/v3 [0]));
 AND2_X1 \V1/V3/V1/V1/_1_  (.A1(net48),
    .A2(net11),
    .ZN(\V1/V3/V1/V1/w1 ));
 AND2_X1 \V1/V3/V1/V1/_2_  (.A1(net12),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V1/w2 ));
 AND2_X1 \V1/V3/V1/V1/_3_  (.A1(net11),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V1/w3 ));
 AND2_X1 \V1/V3/V1/V2/HA1/_0_  (.A1(\V1/V3/V1/V2/w2 ),
    .A2(\V1/V3/V1/V2/w1 ),
    .ZN(\V1/V3/V1/V2/w4 ));
 XOR2_X2 \V1/V3/V1/V2/HA1/_1_  (.A(\V1/V3/V1/V2/w2 ),
    .B(\V1/V3/V1/V2/w1 ),
    .Z(\V1/V3/V1/v2 [1]));
 AND2_X1 \V1/V3/V1/V2/HA2/_0_  (.A1(\V1/V3/V1/V2/w4 ),
    .A2(\V1/V3/V1/V2/w3 ),
    .ZN(\V1/V3/V1/v2 [3]));
 XOR2_X2 \V1/V3/V1/V2/HA2/_1_  (.A(\V1/V3/V1/V2/w4 ),
    .B(\V1/V3/V1/V2/w3 ),
    .Z(\V1/V3/V1/v2 [2]));
 AND2_X1 \V1/V3/V1/V2/_0_  (.A1(A[2]),
    .A2(net12),
    .ZN(\V1/V3/V1/v2 [0]));
 AND2_X1 \V1/V3/V1/V2/_1_  (.A1(A[2]),
    .A2(net11),
    .ZN(\V1/V3/V1/V2/w1 ));
 AND2_X1 \V1/V3/V1/V2/_2_  (.A1(net12),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V2/w2 ));
 AND2_X1 \V1/V3/V1/V2/_3_  (.A1(net11),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V2/w3 ));
 AND2_X1 \V1/V3/V1/V3/HA1/_0_  (.A1(\V1/V3/V1/V3/w2 ),
    .A2(\V1/V3/V1/V3/w1 ),
    .ZN(\V1/V3/V1/V3/w4 ));
 XOR2_X2 \V1/V3/V1/V3/HA1/_1_  (.A(\V1/V3/V1/V3/w2 ),
    .B(\V1/V3/V1/V3/w1 ),
    .Z(\V1/V3/V1/v3 [1]));
 AND2_X1 \V1/V3/V1/V3/HA2/_0_  (.A1(\V1/V3/V1/V3/w4 ),
    .A2(\V1/V3/V1/V3/w3 ),
    .ZN(\V1/V3/V1/v3 [3]));
 XOR2_X2 \V1/V3/V1/V3/HA2/_1_  (.A(\V1/V3/V1/V3/w4 ),
    .B(\V1/V3/V1/V3/w3 ),
    .Z(\V1/V3/V1/v3 [2]));
 AND2_X1 \V1/V3/V1/V3/_0_  (.A1(net48),
    .A2(B[10]),
    .ZN(\V1/V3/V1/v3 [0]));
 AND2_X1 \V1/V3/V1/V3/_1_  (.A1(net48),
    .A2(B[11]),
    .ZN(\V1/V3/V1/V3/w1 ));
 AND2_X1 \V1/V3/V1/V3/_2_  (.A1(B[10]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V3/w2 ));
 AND2_X1 \V1/V3/V1/V3/_3_  (.A1(B[11]),
    .A2(A[1]),
    .ZN(\V1/V3/V1/V3/w3 ));
 AND2_X1 \V1/V3/V1/V4/HA1/_0_  (.A1(\V1/V3/V1/V4/w2 ),
    .A2(\V1/V3/V1/V4/w1 ),
    .ZN(\V1/V3/V1/V4/w4 ));
 XOR2_X2 \V1/V3/V1/V4/HA1/_1_  (.A(\V1/V3/V1/V4/w2 ),
    .B(\V1/V3/V1/V4/w1 ),
    .Z(\V1/V3/V1/v4 [1]));
 AND2_X1 \V1/V3/V1/V4/HA2/_0_  (.A1(\V1/V3/V1/V4/w4 ),
    .A2(\V1/V3/V1/V4/w3 ),
    .ZN(\V1/V3/V1/v4 [3]));
 XOR2_X2 \V1/V3/V1/V4/HA2/_1_  (.A(\V1/V3/V1/V4/w4 ),
    .B(\V1/V3/V1/V4/w3 ),
    .Z(\V1/V3/V1/v4 [2]));
 AND2_X1 \V1/V3/V1/V4/_0_  (.A1(A[2]),
    .A2(B[10]),
    .ZN(\V1/V3/V1/v4 [0]));
 AND2_X1 \V1/V3/V1/V4/_1_  (.A1(A[2]),
    .A2(B[11]),
    .ZN(\V1/V3/V1/V4/w1 ));
 AND2_X1 \V1/V3/V1/V4/_2_  (.A1(B[10]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V4/w2 ));
 AND2_X1 \V1/V3/V1/V4/_3_  (.A1(B[11]),
    .A2(A[3]),
    .ZN(\V1/V3/V1/V4/w3 ));
 OR2_X1 \V1/V3/V1/_0_  (.A1(\V1/V3/V1/c1 ),
    .A2(\V1/V3/V1/c2 ),
    .ZN(\V1/V3/V1/c3 ));
 AND2_X1 \V1/V3/V2/A1/M1/M1/_0_  (.A1(\V1/V3/V2/v2 [0]),
    .A2(\V1/V3/V2/v3 [0]),
    .ZN(\V1/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M1/M1/_1_  (.A(\V1/V3/V2/v2 [0]),
    .B(\V1/V3/V2/v3 [0]),
    .Z(\V1/V3/V2/A1/M1/s1 ));
 AND2_X1 \V1/V3/V2/A1/M1/M2/_0_  (.A1(\V1/V3/V2/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M1/M2/_1_  (.A(\V1/V3/V2/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/V3/V2/s1 [0]));
 OR2_X1 \V1/V3/V2/A1/M1/_0_  (.A1(\V1/V3/V2/A1/M1/c1 ),
    .A2(\V1/V3/V2/A1/M1/c2 ),
    .ZN(\V1/V3/V2/A1/c1 ));
 AND2_X1 \V1/V3/V2/A1/M2/M1/_0_  (.A1(\V1/V3/V2/v2 [1]),
    .A2(\V1/V3/V2/v3 [1]),
    .ZN(\V1/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M2/M1/_1_  (.A(\V1/V3/V2/v2 [1]),
    .B(\V1/V3/V2/v3 [1]),
    .Z(\V1/V3/V2/A1/M2/s1 ));
 AND2_X1 \V1/V3/V2/A1/M2/M2/_0_  (.A1(\V1/V3/V2/A1/M2/s1 ),
    .A2(\V1/V3/V2/A1/c1 ),
    .ZN(\V1/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M2/M2/_1_  (.A(\V1/V3/V2/A1/M2/s1 ),
    .B(\V1/V3/V2/A1/c1 ),
    .Z(\V1/V3/V2/s1 [1]));
 OR2_X1 \V1/V3/V2/A1/M2/_0_  (.A1(\V1/V3/V2/A1/M2/c1 ),
    .A2(\V1/V3/V2/A1/M2/c2 ),
    .ZN(\V1/V3/V2/A1/c2 ));
 AND2_X1 \V1/V3/V2/A1/M3/M1/_0_  (.A1(\V1/V3/V2/v2 [2]),
    .A2(\V1/V3/V2/v3 [2]),
    .ZN(\V1/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M3/M1/_1_  (.A(\V1/V3/V2/v2 [2]),
    .B(\V1/V3/V2/v3 [2]),
    .Z(\V1/V3/V2/A1/M3/s1 ));
 AND2_X1 \V1/V3/V2/A1/M3/M2/_0_  (.A1(\V1/V3/V2/A1/M3/s1 ),
    .A2(\V1/V3/V2/A1/c2 ),
    .ZN(\V1/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M3/M2/_1_  (.A(\V1/V3/V2/A1/M3/s1 ),
    .B(\V1/V3/V2/A1/c2 ),
    .Z(\V1/V3/V2/s1 [2]));
 OR2_X1 \V1/V3/V2/A1/M3/_0_  (.A1(\V1/V3/V2/A1/M3/c1 ),
    .A2(\V1/V3/V2/A1/M3/c2 ),
    .ZN(\V1/V3/V2/A1/c3 ));
 AND2_X1 \V1/V3/V2/A1/M4/M1/_0_  (.A1(\V1/V3/V2/v2 [3]),
    .A2(\V1/V3/V2/v3 [3]),
    .ZN(\V1/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A1/M4/M1/_1_  (.A(\V1/V3/V2/v2 [3]),
    .B(\V1/V3/V2/v3 [3]),
    .Z(\V1/V3/V2/A1/M4/s1 ));
 AND2_X1 \V1/V3/V2/A1/M4/M2/_0_  (.A1(\V1/V3/V2/A1/M4/s1 ),
    .A2(\V1/V3/V2/A1/c3 ),
    .ZN(\V1/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A1/M4/M2/_1_  (.A(\V1/V3/V2/A1/M4/s1 ),
    .B(\V1/V3/V2/A1/c3 ),
    .Z(\V1/V3/V2/s1 [3]));
 OR2_X1 \V1/V3/V2/A1/M4/_0_  (.A1(\V1/V3/V2/A1/M4/c1 ),
    .A2(\V1/V3/V2/A1/M4/c2 ),
    .ZN(\V1/V3/V2/c1 ));
 AND2_X1 \V1/V3/V2/A2/M1/M1/_0_  (.A1(\V1/V3/V2/s1 [0]),
    .A2(\V1/V3/V2/v1 [2]),
    .ZN(\V1/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M1/M1/_1_  (.A(\V1/V3/V2/s1 [0]),
    .B(\V1/V3/V2/v1 [2]),
    .Z(\V1/V3/V2/A2/M1/s1 ));
 AND2_X1 \V1/V3/V2/A2/M1/M2/_0_  (.A1(\V1/V3/V2/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M1/M2/_1_  (.A(\V1/V3/V2/A2/M1/s1 ),
    .B(net5),
    .Z(\V1/V3/v2 [2]));
 OR2_X1 \V1/V3/V2/A2/M1/_0_  (.A1(\V1/V3/V2/A2/M1/c1 ),
    .A2(\V1/V3/V2/A2/M1/c2 ),
    .ZN(\V1/V3/V2/A2/c1 ));
 AND2_X1 \V1/V3/V2/A2/M2/M1/_0_  (.A1(\V1/V3/V2/s1 [1]),
    .A2(\V1/V3/V2/v1 [3]),
    .ZN(\V1/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M2/M1/_1_  (.A(\V1/V3/V2/s1 [1]),
    .B(\V1/V3/V2/v1 [3]),
    .Z(\V1/V3/V2/A2/M2/s1 ));
 AND2_X1 \V1/V3/V2/A2/M2/M2/_0_  (.A1(\V1/V3/V2/A2/M2/s1 ),
    .A2(\V1/V3/V2/A2/c1 ),
    .ZN(\V1/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M2/M2/_1_  (.A(\V1/V3/V2/A2/M2/s1 ),
    .B(\V1/V3/V2/A2/c1 ),
    .Z(\V1/V3/v2 [3]));
 OR2_X1 \V1/V3/V2/A2/M2/_0_  (.A1(\V1/V3/V2/A2/M2/c1 ),
    .A2(\V1/V3/V2/A2/M2/c2 ),
    .ZN(\V1/V3/V2/A2/c2 ));
 AND2_X1 \V1/V3/V2/A2/M3/M1/_0_  (.A1(\V1/V3/V2/s1 [2]),
    .A2(net5),
    .ZN(\V1/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M3/M1/_1_  (.A(\V1/V3/V2/s1 [2]),
    .B(net5),
    .Z(\V1/V3/V2/A2/M3/s1 ));
 AND2_X1 \V1/V3/V2/A2/M3/M2/_0_  (.A1(\V1/V3/V2/A2/M3/s1 ),
    .A2(\V1/V3/V2/A2/c2 ),
    .ZN(\V1/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M3/M2/_1_  (.A(\V1/V3/V2/A2/M3/s1 ),
    .B(\V1/V3/V2/A2/c2 ),
    .Z(\V1/V3/V2/s2 [2]));
 OR2_X1 \V1/V3/V2/A2/M3/_0_  (.A1(\V1/V3/V2/A2/M3/c1 ),
    .A2(\V1/V3/V2/A2/M3/c2 ),
    .ZN(\V1/V3/V2/A2/c3 ));
 AND2_X1 \V1/V3/V2/A2/M4/M1/_0_  (.A1(\V1/V3/V2/s1 [3]),
    .A2(net5),
    .ZN(\V1/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A2/M4/M1/_1_  (.A(\V1/V3/V2/s1 [3]),
    .B(net5),
    .Z(\V1/V3/V2/A2/M4/s1 ));
 AND2_X1 \V1/V3/V2/A2/M4/M2/_0_  (.A1(\V1/V3/V2/A2/M4/s1 ),
    .A2(\V1/V3/V2/A2/c3 ),
    .ZN(\V1/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A2/M4/M2/_1_  (.A(\V1/V3/V2/A2/M4/s1 ),
    .B(\V1/V3/V2/A2/c3 ),
    .Z(\V1/V3/V2/s2 [3]));
 OR2_X1 \V1/V3/V2/A2/M4/_0_  (.A1(\V1/V3/V2/A2/M4/c1 ),
    .A2(\V1/V3/V2/A2/M4/c2 ),
    .ZN(\V1/V3/V2/c2 ));
 AND2_X1 \V1/V3/V2/A3/M1/M1/_0_  (.A1(\V1/V3/V2/v4 [0]),
    .A2(\V1/V3/V2/s2 [2]),
    .ZN(\V1/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M1/M1/_1_  (.A(\V1/V3/V2/v4 [0]),
    .B(\V1/V3/V2/s2 [2]),
    .Z(\V1/V3/V2/A3/M1/s1 ));
 AND2_X1 \V1/V3/V2/A3/M1/M2/_0_  (.A1(\V1/V3/V2/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M1/M2/_1_  (.A(\V1/V3/V2/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V3/v2 [4]));
 OR2_X1 \V1/V3/V2/A3/M1/_0_  (.A1(\V1/V3/V2/A3/M1/c1 ),
    .A2(\V1/V3/V2/A3/M1/c2 ),
    .ZN(\V1/V3/V2/A3/c1 ));
 AND2_X1 \V1/V3/V2/A3/M2/M1/_0_  (.A1(\V1/V3/V2/v4 [1]),
    .A2(\V1/V3/V2/s2 [3]),
    .ZN(\V1/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M2/M1/_1_  (.A(\V1/V3/V2/v4 [1]),
    .B(\V1/V3/V2/s2 [3]),
    .Z(\V1/V3/V2/A3/M2/s1 ));
 AND2_X1 \V1/V3/V2/A3/M2/M2/_0_  (.A1(\V1/V3/V2/A3/M2/s1 ),
    .A2(\V1/V3/V2/A3/c1 ),
    .ZN(\V1/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M2/M2/_1_  (.A(\V1/V3/V2/A3/M2/s1 ),
    .B(\V1/V3/V2/A3/c1 ),
    .Z(\V1/V3/v2 [5]));
 OR2_X1 \V1/V3/V2/A3/M2/_0_  (.A1(\V1/V3/V2/A3/M2/c1 ),
    .A2(\V1/V3/V2/A3/M2/c2 ),
    .ZN(\V1/V3/V2/A3/c2 ));
 AND2_X1 \V1/V3/V2/A3/M3/M1/_0_  (.A1(\V1/V3/V2/v4 [2]),
    .A2(\V1/V3/V2/c3 ),
    .ZN(\V1/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M3/M1/_1_  (.A(\V1/V3/V2/v4 [2]),
    .B(\V1/V3/V2/c3 ),
    .Z(\V1/V3/V2/A3/M3/s1 ));
 AND2_X1 \V1/V3/V2/A3/M3/M2/_0_  (.A1(\V1/V3/V2/A3/M3/s1 ),
    .A2(\V1/V3/V2/A3/c2 ),
    .ZN(\V1/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M3/M2/_1_  (.A(\V1/V3/V2/A3/M3/s1 ),
    .B(\V1/V3/V2/A3/c2 ),
    .Z(\V1/V3/v2 [6]));
 OR2_X1 \V1/V3/V2/A3/M3/_0_  (.A1(\V1/V3/V2/A3/M3/c1 ),
    .A2(\V1/V3/V2/A3/M3/c2 ),
    .ZN(\V1/V3/V2/A3/c3 ));
 AND2_X1 \V1/V3/V2/A3/M4/M1/_0_  (.A1(\V1/V3/V2/v4 [3]),
    .A2(net5),
    .ZN(\V1/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V2/A3/M4/M1/_1_  (.A(\V1/V3/V2/v4 [3]),
    .B(net5),
    .Z(\V1/V3/V2/A3/M4/s1 ));
 AND2_X1 \V1/V3/V2/A3/M4/M2/_0_  (.A1(\V1/V3/V2/A3/M4/s1 ),
    .A2(\V1/V3/V2/A3/c3 ),
    .ZN(\V1/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V2/A3/M4/M2/_1_  (.A(\V1/V3/V2/A3/M4/s1 ),
    .B(\V1/V3/V2/A3/c3 ),
    .Z(\V1/V3/v2 [7]));
 OR2_X1 \V1/V3/V2/A3/M4/_0_  (.A1(\V1/V3/V2/A3/M4/c1 ),
    .A2(\V1/V3/V2/A3/M4/c2 ),
    .ZN(\V1/V3/V2/overflow ));
 AND2_X1 \V1/V3/V2/V1/HA1/_0_  (.A1(\V1/V3/V2/V1/w2 ),
    .A2(\V1/V3/V2/V1/w1 ),
    .ZN(\V1/V3/V2/V1/w4 ));
 XOR2_X2 \V1/V3/V2/V1/HA1/_1_  (.A(\V1/V3/V2/V1/w2 ),
    .B(\V1/V3/V2/V1/w1 ),
    .Z(\V1/V3/v2 [1]));
 AND2_X1 \V1/V3/V2/V1/HA2/_0_  (.A1(\V1/V3/V2/V1/w4 ),
    .A2(\V1/V3/V2/V1/w3 ),
    .ZN(\V1/V3/V2/v1 [3]));
 XOR2_X2 \V1/V3/V2/V1/HA2/_1_  (.A(\V1/V3/V2/V1/w4 ),
    .B(\V1/V3/V2/V1/w3 ),
    .Z(\V1/V3/V2/v1 [2]));
 AND2_X1 \V1/V3/V2/V1/_0_  (.A1(A[4]),
    .A2(net12),
    .ZN(\V1/V3/v2 [0]));
 AND2_X1 \V1/V3/V2/V1/_1_  (.A1(A[4]),
    .A2(net11),
    .ZN(\V1/V3/V2/V1/w1 ));
 AND2_X1 \V1/V3/V2/V1/_2_  (.A1(net12),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V1/w2 ));
 AND2_X1 \V1/V3/V2/V1/_3_  (.A1(net11),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V1/w3 ));
 AND2_X1 \V1/V3/V2/V2/HA1/_0_  (.A1(\V1/V3/V2/V2/w2 ),
    .A2(\V1/V3/V2/V2/w1 ),
    .ZN(\V1/V3/V2/V2/w4 ));
 XOR2_X2 \V1/V3/V2/V2/HA1/_1_  (.A(\V1/V3/V2/V2/w2 ),
    .B(\V1/V3/V2/V2/w1 ),
    .Z(\V1/V3/V2/v2 [1]));
 AND2_X1 \V1/V3/V2/V2/HA2/_0_  (.A1(\V1/V3/V2/V2/w4 ),
    .A2(\V1/V3/V2/V2/w3 ),
    .ZN(\V1/V3/V2/v2 [3]));
 XOR2_X2 \V1/V3/V2/V2/HA2/_1_  (.A(\V1/V3/V2/V2/w4 ),
    .B(\V1/V3/V2/V2/w3 ),
    .Z(\V1/V3/V2/v2 [2]));
 AND2_X1 \V1/V3/V2/V2/_0_  (.A1(A[6]),
    .A2(net12),
    .ZN(\V1/V3/V2/v2 [0]));
 AND2_X1 \V1/V3/V2/V2/_1_  (.A1(A[6]),
    .A2(net11),
    .ZN(\V1/V3/V2/V2/w1 ));
 AND2_X1 \V1/V3/V2/V2/_2_  (.A1(net12),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V2/w2 ));
 AND2_X1 \V1/V3/V2/V2/_3_  (.A1(net11),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V2/w3 ));
 AND2_X1 \V1/V3/V2/V3/HA1/_0_  (.A1(\V1/V3/V2/V3/w2 ),
    .A2(\V1/V3/V2/V3/w1 ),
    .ZN(\V1/V3/V2/V3/w4 ));
 XOR2_X2 \V1/V3/V2/V3/HA1/_1_  (.A(\V1/V3/V2/V3/w2 ),
    .B(\V1/V3/V2/V3/w1 ),
    .Z(\V1/V3/V2/v3 [1]));
 AND2_X1 \V1/V3/V2/V3/HA2/_0_  (.A1(\V1/V3/V2/V3/w4 ),
    .A2(\V1/V3/V2/V3/w3 ),
    .ZN(\V1/V3/V2/v3 [3]));
 XOR2_X2 \V1/V3/V2/V3/HA2/_1_  (.A(\V1/V3/V2/V3/w4 ),
    .B(\V1/V3/V2/V3/w3 ),
    .Z(\V1/V3/V2/v3 [2]));
 AND2_X1 \V1/V3/V2/V3/_0_  (.A1(A[4]),
    .A2(B[10]),
    .ZN(\V1/V3/V2/v3 [0]));
 AND2_X1 \V1/V3/V2/V3/_1_  (.A1(A[4]),
    .A2(B[11]),
    .ZN(\V1/V3/V2/V3/w1 ));
 AND2_X1 \V1/V3/V2/V3/_2_  (.A1(B[10]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V3/w2 ));
 AND2_X1 \V1/V3/V2/V3/_3_  (.A1(B[11]),
    .A2(A[5]),
    .ZN(\V1/V3/V2/V3/w3 ));
 AND2_X1 \V1/V3/V2/V4/HA1/_0_  (.A1(\V1/V3/V2/V4/w2 ),
    .A2(\V1/V3/V2/V4/w1 ),
    .ZN(\V1/V3/V2/V4/w4 ));
 XOR2_X2 \V1/V3/V2/V4/HA1/_1_  (.A(\V1/V3/V2/V4/w2 ),
    .B(\V1/V3/V2/V4/w1 ),
    .Z(\V1/V3/V2/v4 [1]));
 AND2_X1 \V1/V3/V2/V4/HA2/_0_  (.A1(\V1/V3/V2/V4/w4 ),
    .A2(\V1/V3/V2/V4/w3 ),
    .ZN(\V1/V3/V2/v4 [3]));
 XOR2_X2 \V1/V3/V2/V4/HA2/_1_  (.A(\V1/V3/V2/V4/w4 ),
    .B(\V1/V3/V2/V4/w3 ),
    .Z(\V1/V3/V2/v4 [2]));
 AND2_X1 \V1/V3/V2/V4/_0_  (.A1(A[6]),
    .A2(B[10]),
    .ZN(\V1/V3/V2/v4 [0]));
 AND2_X1 \V1/V3/V2/V4/_1_  (.A1(A[6]),
    .A2(B[11]),
    .ZN(\V1/V3/V2/V4/w1 ));
 AND2_X1 \V1/V3/V2/V4/_2_  (.A1(B[10]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V4/w2 ));
 AND2_X1 \V1/V3/V2/V4/_3_  (.A1(B[11]),
    .A2(A[7]),
    .ZN(\V1/V3/V2/V4/w3 ));
 OR2_X1 \V1/V3/V2/_0_  (.A1(\V1/V3/V2/c1 ),
    .A2(\V1/V3/V2/c2 ),
    .ZN(\V1/V3/V2/c3 ));
 AND2_X1 \V1/V3/V3/A1/M1/M1/_0_  (.A1(\V1/V3/V3/v2 [0]),
    .A2(\V1/V3/V3/v3 [0]),
    .ZN(\V1/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M1/M1/_1_  (.A(\V1/V3/V3/v2 [0]),
    .B(\V1/V3/V3/v3 [0]),
    .Z(\V1/V3/V3/A1/M1/s1 ));
 AND2_X1 \V1/V3/V3/A1/M1/M2/_0_  (.A1(\V1/V3/V3/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M1/M2/_1_  (.A(\V1/V3/V3/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/V3/V3/s1 [0]));
 OR2_X1 \V1/V3/V3/A1/M1/_0_  (.A1(\V1/V3/V3/A1/M1/c1 ),
    .A2(\V1/V3/V3/A1/M1/c2 ),
    .ZN(\V1/V3/V3/A1/c1 ));
 AND2_X1 \V1/V3/V3/A1/M2/M1/_0_  (.A1(\V1/V3/V3/v2 [1]),
    .A2(\V1/V3/V3/v3 [1]),
    .ZN(\V1/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M2/M1/_1_  (.A(\V1/V3/V3/v2 [1]),
    .B(\V1/V3/V3/v3 [1]),
    .Z(\V1/V3/V3/A1/M2/s1 ));
 AND2_X1 \V1/V3/V3/A1/M2/M2/_0_  (.A1(\V1/V3/V3/A1/M2/s1 ),
    .A2(\V1/V3/V3/A1/c1 ),
    .ZN(\V1/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M2/M2/_1_  (.A(\V1/V3/V3/A1/M2/s1 ),
    .B(\V1/V3/V3/A1/c1 ),
    .Z(\V1/V3/V3/s1 [1]));
 OR2_X1 \V1/V3/V3/A1/M2/_0_  (.A1(\V1/V3/V3/A1/M2/c1 ),
    .A2(\V1/V3/V3/A1/M2/c2 ),
    .ZN(\V1/V3/V3/A1/c2 ));
 AND2_X1 \V1/V3/V3/A1/M3/M1/_0_  (.A1(\V1/V3/V3/v2 [2]),
    .A2(\V1/V3/V3/v3 [2]),
    .ZN(\V1/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M3/M1/_1_  (.A(\V1/V3/V3/v2 [2]),
    .B(\V1/V3/V3/v3 [2]),
    .Z(\V1/V3/V3/A1/M3/s1 ));
 AND2_X1 \V1/V3/V3/A1/M3/M2/_0_  (.A1(\V1/V3/V3/A1/M3/s1 ),
    .A2(\V1/V3/V3/A1/c2 ),
    .ZN(\V1/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M3/M2/_1_  (.A(\V1/V3/V3/A1/M3/s1 ),
    .B(\V1/V3/V3/A1/c2 ),
    .Z(\V1/V3/V3/s1 [2]));
 OR2_X1 \V1/V3/V3/A1/M3/_0_  (.A1(\V1/V3/V3/A1/M3/c1 ),
    .A2(\V1/V3/V3/A1/M3/c2 ),
    .ZN(\V1/V3/V3/A1/c3 ));
 AND2_X1 \V1/V3/V3/A1/M4/M1/_0_  (.A1(\V1/V3/V3/v2 [3]),
    .A2(\V1/V3/V3/v3 [3]),
    .ZN(\V1/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A1/M4/M1/_1_  (.A(\V1/V3/V3/v2 [3]),
    .B(\V1/V3/V3/v3 [3]),
    .Z(\V1/V3/V3/A1/M4/s1 ));
 AND2_X1 \V1/V3/V3/A1/M4/M2/_0_  (.A1(\V1/V3/V3/A1/M4/s1 ),
    .A2(\V1/V3/V3/A1/c3 ),
    .ZN(\V1/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A1/M4/M2/_1_  (.A(\V1/V3/V3/A1/M4/s1 ),
    .B(\V1/V3/V3/A1/c3 ),
    .Z(\V1/V3/V3/s1 [3]));
 OR2_X1 \V1/V3/V3/A1/M4/_0_  (.A1(\V1/V3/V3/A1/M4/c1 ),
    .A2(\V1/V3/V3/A1/M4/c2 ),
    .ZN(\V1/V3/V3/c1 ));
 AND2_X1 \V1/V3/V3/A2/M1/M1/_0_  (.A1(\V1/V3/V3/s1 [0]),
    .A2(\V1/V3/V3/v1 [2]),
    .ZN(\V1/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M1/M1/_1_  (.A(\V1/V3/V3/s1 [0]),
    .B(\V1/V3/V3/v1 [2]),
    .Z(\V1/V3/V3/A2/M1/s1 ));
 AND2_X1 \V1/V3/V3/A2/M1/M2/_0_  (.A1(\V1/V3/V3/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M1/M2/_1_  (.A(\V1/V3/V3/A2/M1/s1 ),
    .B(net5),
    .Z(\V1/V3/v3 [2]));
 OR2_X1 \V1/V3/V3/A2/M1/_0_  (.A1(\V1/V3/V3/A2/M1/c1 ),
    .A2(\V1/V3/V3/A2/M1/c2 ),
    .ZN(\V1/V3/V3/A2/c1 ));
 AND2_X1 \V1/V3/V3/A2/M2/M1/_0_  (.A1(\V1/V3/V3/s1 [1]),
    .A2(\V1/V3/V3/v1 [3]),
    .ZN(\V1/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M2/M1/_1_  (.A(\V1/V3/V3/s1 [1]),
    .B(\V1/V3/V3/v1 [3]),
    .Z(\V1/V3/V3/A2/M2/s1 ));
 AND2_X1 \V1/V3/V3/A2/M2/M2/_0_  (.A1(\V1/V3/V3/A2/M2/s1 ),
    .A2(\V1/V3/V3/A2/c1 ),
    .ZN(\V1/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M2/M2/_1_  (.A(\V1/V3/V3/A2/M2/s1 ),
    .B(\V1/V3/V3/A2/c1 ),
    .Z(\V1/V3/v3 [3]));
 OR2_X1 \V1/V3/V3/A2/M2/_0_  (.A1(\V1/V3/V3/A2/M2/c1 ),
    .A2(\V1/V3/V3/A2/M2/c2 ),
    .ZN(\V1/V3/V3/A2/c2 ));
 AND2_X1 \V1/V3/V3/A2/M3/M1/_0_  (.A1(\V1/V3/V3/s1 [2]),
    .A2(net5),
    .ZN(\V1/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M3/M1/_1_  (.A(\V1/V3/V3/s1 [2]),
    .B(net5),
    .Z(\V1/V3/V3/A2/M3/s1 ));
 AND2_X1 \V1/V3/V3/A2/M3/M2/_0_  (.A1(\V1/V3/V3/A2/M3/s1 ),
    .A2(\V1/V3/V3/A2/c2 ),
    .ZN(\V1/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M3/M2/_1_  (.A(\V1/V3/V3/A2/M3/s1 ),
    .B(\V1/V3/V3/A2/c2 ),
    .Z(\V1/V3/V3/s2 [2]));
 OR2_X1 \V1/V3/V3/A2/M3/_0_  (.A1(\V1/V3/V3/A2/M3/c1 ),
    .A2(\V1/V3/V3/A2/M3/c2 ),
    .ZN(\V1/V3/V3/A2/c3 ));
 AND2_X1 \V1/V3/V3/A2/M4/M1/_0_  (.A1(\V1/V3/V3/s1 [3]),
    .A2(net5),
    .ZN(\V1/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A2/M4/M1/_1_  (.A(\V1/V3/V3/s1 [3]),
    .B(net5),
    .Z(\V1/V3/V3/A2/M4/s1 ));
 AND2_X1 \V1/V3/V3/A2/M4/M2/_0_  (.A1(\V1/V3/V3/A2/M4/s1 ),
    .A2(\V1/V3/V3/A2/c3 ),
    .ZN(\V1/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A2/M4/M2/_1_  (.A(\V1/V3/V3/A2/M4/s1 ),
    .B(\V1/V3/V3/A2/c3 ),
    .Z(\V1/V3/V3/s2 [3]));
 OR2_X1 \V1/V3/V3/A2/M4/_0_  (.A1(\V1/V3/V3/A2/M4/c1 ),
    .A2(\V1/V3/V3/A2/M4/c2 ),
    .ZN(\V1/V3/V3/c2 ));
 AND2_X1 \V1/V3/V3/A3/M1/M1/_0_  (.A1(\V1/V3/V3/v4 [0]),
    .A2(\V1/V3/V3/s2 [2]),
    .ZN(\V1/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M1/M1/_1_  (.A(\V1/V3/V3/v4 [0]),
    .B(\V1/V3/V3/s2 [2]),
    .Z(\V1/V3/V3/A3/M1/s1 ));
 AND2_X1 \V1/V3/V3/A3/M1/M2/_0_  (.A1(\V1/V3/V3/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M1/M2/_1_  (.A(\V1/V3/V3/A3/M1/s1 ),
    .B(net5),
    .Z(\V1/V3/v3 [4]));
 OR2_X1 \V1/V3/V3/A3/M1/_0_  (.A1(\V1/V3/V3/A3/M1/c1 ),
    .A2(\V1/V3/V3/A3/M1/c2 ),
    .ZN(\V1/V3/V3/A3/c1 ));
 AND2_X1 \V1/V3/V3/A3/M2/M1/_0_  (.A1(\V1/V3/V3/v4 [1]),
    .A2(\V1/V3/V3/s2 [3]),
    .ZN(\V1/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M2/M1/_1_  (.A(\V1/V3/V3/v4 [1]),
    .B(\V1/V3/V3/s2 [3]),
    .Z(\V1/V3/V3/A3/M2/s1 ));
 AND2_X1 \V1/V3/V3/A3/M2/M2/_0_  (.A1(\V1/V3/V3/A3/M2/s1 ),
    .A2(\V1/V3/V3/A3/c1 ),
    .ZN(\V1/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M2/M2/_1_  (.A(\V1/V3/V3/A3/M2/s1 ),
    .B(\V1/V3/V3/A3/c1 ),
    .Z(\V1/V3/v3 [5]));
 OR2_X1 \V1/V3/V3/A3/M2/_0_  (.A1(\V1/V3/V3/A3/M2/c1 ),
    .A2(\V1/V3/V3/A3/M2/c2 ),
    .ZN(\V1/V3/V3/A3/c2 ));
 AND2_X1 \V1/V3/V3/A3/M3/M1/_0_  (.A1(\V1/V3/V3/v4 [2]),
    .A2(\V1/V3/V3/c3 ),
    .ZN(\V1/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M3/M1/_1_  (.A(\V1/V3/V3/v4 [2]),
    .B(\V1/V3/V3/c3 ),
    .Z(\V1/V3/V3/A3/M3/s1 ));
 AND2_X1 \V1/V3/V3/A3/M3/M2/_0_  (.A1(\V1/V3/V3/A3/M3/s1 ),
    .A2(\V1/V3/V3/A3/c2 ),
    .ZN(\V1/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M3/M2/_1_  (.A(\V1/V3/V3/A3/M3/s1 ),
    .B(\V1/V3/V3/A3/c2 ),
    .Z(\V1/V3/v3 [6]));
 OR2_X1 \V1/V3/V3/A3/M3/_0_  (.A1(\V1/V3/V3/A3/M3/c1 ),
    .A2(\V1/V3/V3/A3/M3/c2 ),
    .ZN(\V1/V3/V3/A3/c3 ));
 AND2_X1 \V1/V3/V3/A3/M4/M1/_0_  (.A1(\V1/V3/V3/v4 [3]),
    .A2(net5),
    .ZN(\V1/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V3/A3/M4/M1/_1_  (.A(\V1/V3/V3/v4 [3]),
    .B(net5),
    .Z(\V1/V3/V3/A3/M4/s1 ));
 AND2_X1 \V1/V3/V3/A3/M4/M2/_0_  (.A1(\V1/V3/V3/A3/M4/s1 ),
    .A2(\V1/V3/V3/A3/c3 ),
    .ZN(\V1/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V3/A3/M4/M2/_1_  (.A(\V1/V3/V3/A3/M4/s1 ),
    .B(\V1/V3/V3/A3/c3 ),
    .Z(\V1/V3/v3 [7]));
 OR2_X1 \V1/V3/V3/A3/M4/_0_  (.A1(\V1/V3/V3/A3/M4/c1 ),
    .A2(\V1/V3/V3/A3/M4/c2 ),
    .ZN(\V1/V3/V3/overflow ));
 AND2_X1 \V1/V3/V3/V1/HA1/_0_  (.A1(\V1/V3/V3/V1/w2 ),
    .A2(\V1/V3/V3/V1/w1 ),
    .ZN(\V1/V3/V3/V1/w4 ));
 XOR2_X2 \V1/V3/V3/V1/HA1/_1_  (.A(\V1/V3/V3/V1/w2 ),
    .B(\V1/V3/V3/V1/w1 ),
    .Z(\V1/V3/v3 [1]));
 AND2_X1 \V1/V3/V3/V1/HA2/_0_  (.A1(\V1/V3/V3/V1/w4 ),
    .A2(\V1/V3/V3/V1/w3 ),
    .ZN(\V1/V3/V3/v1 [3]));
 XOR2_X2 \V1/V3/V3/V1/HA2/_1_  (.A(\V1/V3/V3/V1/w4 ),
    .B(\V1/V3/V3/V1/w3 ),
    .Z(\V1/V3/V3/v1 [2]));
 AND2_X1 \V1/V3/V3/V1/_0_  (.A1(net48),
    .A2(B[12]),
    .ZN(\V1/V3/v3 [0]));
 AND2_X1 \V1/V3/V3/V1/_1_  (.A1(net48),
    .A2(B[13]),
    .ZN(\V1/V3/V3/V1/w1 ));
 AND2_X1 \V1/V3/V3/V1/_2_  (.A1(B[12]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V1/w2 ));
 AND2_X1 \V1/V3/V3/V1/_3_  (.A1(B[13]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V1/w3 ));
 AND2_X1 \V1/V3/V3/V2/HA1/_0_  (.A1(\V1/V3/V3/V2/w2 ),
    .A2(\V1/V3/V3/V2/w1 ),
    .ZN(\V1/V3/V3/V2/w4 ));
 XOR2_X2 \V1/V3/V3/V2/HA1/_1_  (.A(\V1/V3/V3/V2/w2 ),
    .B(\V1/V3/V3/V2/w1 ),
    .Z(\V1/V3/V3/v2 [1]));
 AND2_X1 \V1/V3/V3/V2/HA2/_0_  (.A1(\V1/V3/V3/V2/w4 ),
    .A2(\V1/V3/V3/V2/w3 ),
    .ZN(\V1/V3/V3/v2 [3]));
 XOR2_X2 \V1/V3/V3/V2/HA2/_1_  (.A(\V1/V3/V3/V2/w4 ),
    .B(\V1/V3/V3/V2/w3 ),
    .Z(\V1/V3/V3/v2 [2]));
 AND2_X1 \V1/V3/V3/V2/_0_  (.A1(A[2]),
    .A2(B[12]),
    .ZN(\V1/V3/V3/v2 [0]));
 AND2_X1 \V1/V3/V3/V2/_1_  (.A1(A[2]),
    .A2(B[13]),
    .ZN(\V1/V3/V3/V2/w1 ));
 AND2_X1 \V1/V3/V3/V2/_2_  (.A1(B[12]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V2/w2 ));
 AND2_X1 \V1/V3/V3/V2/_3_  (.A1(B[13]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V2/w3 ));
 AND2_X1 \V1/V3/V3/V3/HA1/_0_  (.A1(\V1/V3/V3/V3/w2 ),
    .A2(\V1/V3/V3/V3/w1 ),
    .ZN(\V1/V3/V3/V3/w4 ));
 XOR2_X2 \V1/V3/V3/V3/HA1/_1_  (.A(\V1/V3/V3/V3/w2 ),
    .B(\V1/V3/V3/V3/w1 ),
    .Z(\V1/V3/V3/v3 [1]));
 AND2_X1 \V1/V3/V3/V3/HA2/_0_  (.A1(\V1/V3/V3/V3/w4 ),
    .A2(\V1/V3/V3/V3/w3 ),
    .ZN(\V1/V3/V3/v3 [3]));
 XOR2_X2 \V1/V3/V3/V3/HA2/_1_  (.A(\V1/V3/V3/V3/w4 ),
    .B(\V1/V3/V3/V3/w3 ),
    .Z(\V1/V3/V3/v3 [2]));
 AND2_X1 \V1/V3/V3/V3/_0_  (.A1(net48),
    .A2(B[14]),
    .ZN(\V1/V3/V3/v3 [0]));
 AND2_X1 \V1/V3/V3/V3/_1_  (.A1(net48),
    .A2(B[15]),
    .ZN(\V1/V3/V3/V3/w1 ));
 AND2_X1 \V1/V3/V3/V3/_2_  (.A1(B[14]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V3/w2 ));
 AND2_X1 \V1/V3/V3/V3/_3_  (.A1(B[15]),
    .A2(A[1]),
    .ZN(\V1/V3/V3/V3/w3 ));
 AND2_X1 \V1/V3/V3/V4/HA1/_0_  (.A1(\V1/V3/V3/V4/w2 ),
    .A2(\V1/V3/V3/V4/w1 ),
    .ZN(\V1/V3/V3/V4/w4 ));
 XOR2_X2 \V1/V3/V3/V4/HA1/_1_  (.A(\V1/V3/V3/V4/w2 ),
    .B(\V1/V3/V3/V4/w1 ),
    .Z(\V1/V3/V3/v4 [1]));
 AND2_X1 \V1/V3/V3/V4/HA2/_0_  (.A1(\V1/V3/V3/V4/w4 ),
    .A2(\V1/V3/V3/V4/w3 ),
    .ZN(\V1/V3/V3/v4 [3]));
 XOR2_X2 \V1/V3/V3/V4/HA2/_1_  (.A(\V1/V3/V3/V4/w4 ),
    .B(\V1/V3/V3/V4/w3 ),
    .Z(\V1/V3/V3/v4 [2]));
 AND2_X1 \V1/V3/V3/V4/_0_  (.A1(A[2]),
    .A2(B[14]),
    .ZN(\V1/V3/V3/v4 [0]));
 AND2_X1 \V1/V3/V3/V4/_1_  (.A1(A[2]),
    .A2(B[15]),
    .ZN(\V1/V3/V3/V4/w1 ));
 AND2_X1 \V1/V3/V3/V4/_2_  (.A1(B[14]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V4/w2 ));
 AND2_X1 \V1/V3/V3/V4/_3_  (.A1(B[15]),
    .A2(A[3]),
    .ZN(\V1/V3/V3/V4/w3 ));
 OR2_X1 \V1/V3/V3/_0_  (.A1(\V1/V3/V3/c1 ),
    .A2(\V1/V3/V3/c2 ),
    .ZN(\V1/V3/V3/c3 ));
 AND2_X1 \V1/V3/V4/A1/M1/M1/_0_  (.A1(\V1/V3/V4/v2 [0]),
    .A2(\V1/V3/V4/v3 [0]),
    .ZN(\V1/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M1/M1/_1_  (.A(\V1/V3/V4/v2 [0]),
    .B(\V1/V3/V4/v3 [0]),
    .Z(\V1/V3/V4/A1/M1/s1 ));
 AND2_X1 \V1/V3/V4/A1/M1/M2/_0_  (.A1(\V1/V3/V4/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M1/M2/_1_  (.A(\V1/V3/V4/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V3/V4/s1 [0]));
 OR2_X1 \V1/V3/V4/A1/M1/_0_  (.A1(\V1/V3/V4/A1/M1/c1 ),
    .A2(\V1/V3/V4/A1/M1/c2 ),
    .ZN(\V1/V3/V4/A1/c1 ));
 AND2_X1 \V1/V3/V4/A1/M2/M1/_0_  (.A1(\V1/V3/V4/v2 [1]),
    .A2(\V1/V3/V4/v3 [1]),
    .ZN(\V1/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M2/M1/_1_  (.A(\V1/V3/V4/v2 [1]),
    .B(\V1/V3/V4/v3 [1]),
    .Z(\V1/V3/V4/A1/M2/s1 ));
 AND2_X1 \V1/V3/V4/A1/M2/M2/_0_  (.A1(\V1/V3/V4/A1/M2/s1 ),
    .A2(\V1/V3/V4/A1/c1 ),
    .ZN(\V1/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M2/M2/_1_  (.A(\V1/V3/V4/A1/M2/s1 ),
    .B(\V1/V3/V4/A1/c1 ),
    .Z(\V1/V3/V4/s1 [1]));
 OR2_X1 \V1/V3/V4/A1/M2/_0_  (.A1(\V1/V3/V4/A1/M2/c1 ),
    .A2(\V1/V3/V4/A1/M2/c2 ),
    .ZN(\V1/V3/V4/A1/c2 ));
 AND2_X1 \V1/V3/V4/A1/M3/M1/_0_  (.A1(\V1/V3/V4/v2 [2]),
    .A2(\V1/V3/V4/v3 [2]),
    .ZN(\V1/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M3/M1/_1_  (.A(\V1/V3/V4/v2 [2]),
    .B(\V1/V3/V4/v3 [2]),
    .Z(\V1/V3/V4/A1/M3/s1 ));
 AND2_X1 \V1/V3/V4/A1/M3/M2/_0_  (.A1(\V1/V3/V4/A1/M3/s1 ),
    .A2(\V1/V3/V4/A1/c2 ),
    .ZN(\V1/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M3/M2/_1_  (.A(\V1/V3/V4/A1/M3/s1 ),
    .B(\V1/V3/V4/A1/c2 ),
    .Z(\V1/V3/V4/s1 [2]));
 OR2_X1 \V1/V3/V4/A1/M3/_0_  (.A1(\V1/V3/V4/A1/M3/c1 ),
    .A2(\V1/V3/V4/A1/M3/c2 ),
    .ZN(\V1/V3/V4/A1/c3 ));
 AND2_X1 \V1/V3/V4/A1/M4/M1/_0_  (.A1(\V1/V3/V4/v2 [3]),
    .A2(\V1/V3/V4/v3 [3]),
    .ZN(\V1/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A1/M4/M1/_1_  (.A(\V1/V3/V4/v2 [3]),
    .B(\V1/V3/V4/v3 [3]),
    .Z(\V1/V3/V4/A1/M4/s1 ));
 AND2_X1 \V1/V3/V4/A1/M4/M2/_0_  (.A1(\V1/V3/V4/A1/M4/s1 ),
    .A2(\V1/V3/V4/A1/c3 ),
    .ZN(\V1/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A1/M4/M2/_1_  (.A(\V1/V3/V4/A1/M4/s1 ),
    .B(\V1/V3/V4/A1/c3 ),
    .Z(\V1/V3/V4/s1 [3]));
 OR2_X1 \V1/V3/V4/A1/M4/_0_  (.A1(\V1/V3/V4/A1/M4/c1 ),
    .A2(\V1/V3/V4/A1/M4/c2 ),
    .ZN(\V1/V3/V4/c1 ));
 AND2_X1 \V1/V3/V4/A2/M1/M1/_0_  (.A1(\V1/V3/V4/s1 [0]),
    .A2(\V1/V3/V4/v1 [2]),
    .ZN(\V1/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M1/M1/_1_  (.A(\V1/V3/V4/s1 [0]),
    .B(\V1/V3/V4/v1 [2]),
    .Z(\V1/V3/V4/A2/M1/s1 ));
 AND2_X1 \V1/V3/V4/A2/M1/M2/_0_  (.A1(\V1/V3/V4/A2/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M1/M2/_1_  (.A(\V1/V3/V4/A2/M1/s1 ),
    .B(net3),
    .Z(\V1/V3/v4 [2]));
 OR2_X1 \V1/V3/V4/A2/M1/_0_  (.A1(\V1/V3/V4/A2/M1/c1 ),
    .A2(\V1/V3/V4/A2/M1/c2 ),
    .ZN(\V1/V3/V4/A2/c1 ));
 AND2_X1 \V1/V3/V4/A2/M2/M1/_0_  (.A1(\V1/V3/V4/s1 [1]),
    .A2(\V1/V3/V4/v1 [3]),
    .ZN(\V1/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M2/M1/_1_  (.A(\V1/V3/V4/s1 [1]),
    .B(\V1/V3/V4/v1 [3]),
    .Z(\V1/V3/V4/A2/M2/s1 ));
 AND2_X1 \V1/V3/V4/A2/M2/M2/_0_  (.A1(\V1/V3/V4/A2/M2/s1 ),
    .A2(\V1/V3/V4/A2/c1 ),
    .ZN(\V1/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M2/M2/_1_  (.A(\V1/V3/V4/A2/M2/s1 ),
    .B(\V1/V3/V4/A2/c1 ),
    .Z(\V1/V3/v4 [3]));
 OR2_X1 \V1/V3/V4/A2/M2/_0_  (.A1(\V1/V3/V4/A2/M2/c1 ),
    .A2(\V1/V3/V4/A2/M2/c2 ),
    .ZN(\V1/V3/V4/A2/c2 ));
 AND2_X1 \V1/V3/V4/A2/M3/M1/_0_  (.A1(\V1/V3/V4/s1 [2]),
    .A2(net3),
    .ZN(\V1/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M3/M1/_1_  (.A(\V1/V3/V4/s1 [2]),
    .B(net3),
    .Z(\V1/V3/V4/A2/M3/s1 ));
 AND2_X1 \V1/V3/V4/A2/M3/M2/_0_  (.A1(\V1/V3/V4/A2/M3/s1 ),
    .A2(\V1/V3/V4/A2/c2 ),
    .ZN(\V1/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M3/M2/_1_  (.A(\V1/V3/V4/A2/M3/s1 ),
    .B(\V1/V3/V4/A2/c2 ),
    .Z(\V1/V3/V4/s2 [2]));
 OR2_X1 \V1/V3/V4/A2/M3/_0_  (.A1(\V1/V3/V4/A2/M3/c1 ),
    .A2(\V1/V3/V4/A2/M3/c2 ),
    .ZN(\V1/V3/V4/A2/c3 ));
 AND2_X1 \V1/V3/V4/A2/M4/M1/_0_  (.A1(\V1/V3/V4/s1 [3]),
    .A2(net3),
    .ZN(\V1/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A2/M4/M1/_1_  (.A(\V1/V3/V4/s1 [3]),
    .B(net3),
    .Z(\V1/V3/V4/A2/M4/s1 ));
 AND2_X1 \V1/V3/V4/A2/M4/M2/_0_  (.A1(\V1/V3/V4/A2/M4/s1 ),
    .A2(\V1/V3/V4/A2/c3 ),
    .ZN(\V1/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A2/M4/M2/_1_  (.A(\V1/V3/V4/A2/M4/s1 ),
    .B(\V1/V3/V4/A2/c3 ),
    .Z(\V1/V3/V4/s2 [3]));
 OR2_X1 \V1/V3/V4/A2/M4/_0_  (.A1(\V1/V3/V4/A2/M4/c1 ),
    .A2(\V1/V3/V4/A2/M4/c2 ),
    .ZN(\V1/V3/V4/c2 ));
 AND2_X1 \V1/V3/V4/A3/M1/M1/_0_  (.A1(\V1/V3/V4/v4 [0]),
    .A2(\V1/V3/V4/s2 [2]),
    .ZN(\V1/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M1/M1/_1_  (.A(\V1/V3/V4/v4 [0]),
    .B(\V1/V3/V4/s2 [2]),
    .Z(\V1/V3/V4/A3/M1/s1 ));
 AND2_X1 \V1/V3/V4/A3/M1/M2/_0_  (.A1(\V1/V3/V4/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M1/M2/_1_  (.A(\V1/V3/V4/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V3/v4 [4]));
 OR2_X1 \V1/V3/V4/A3/M1/_0_  (.A1(\V1/V3/V4/A3/M1/c1 ),
    .A2(\V1/V3/V4/A3/M1/c2 ),
    .ZN(\V1/V3/V4/A3/c1 ));
 AND2_X1 \V1/V3/V4/A3/M2/M1/_0_  (.A1(\V1/V3/V4/v4 [1]),
    .A2(\V1/V3/V4/s2 [3]),
    .ZN(\V1/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M2/M1/_1_  (.A(\V1/V3/V4/v4 [1]),
    .B(\V1/V3/V4/s2 [3]),
    .Z(\V1/V3/V4/A3/M2/s1 ));
 AND2_X1 \V1/V3/V4/A3/M2/M2/_0_  (.A1(\V1/V3/V4/A3/M2/s1 ),
    .A2(\V1/V3/V4/A3/c1 ),
    .ZN(\V1/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M2/M2/_1_  (.A(\V1/V3/V4/A3/M2/s1 ),
    .B(\V1/V3/V4/A3/c1 ),
    .Z(\V1/V3/v4 [5]));
 OR2_X1 \V1/V3/V4/A3/M2/_0_  (.A1(\V1/V3/V4/A3/M2/c1 ),
    .A2(\V1/V3/V4/A3/M2/c2 ),
    .ZN(\V1/V3/V4/A3/c2 ));
 AND2_X1 \V1/V3/V4/A3/M3/M1/_0_  (.A1(\V1/V3/V4/v4 [2]),
    .A2(\V1/V3/V4/c3 ),
    .ZN(\V1/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M3/M1/_1_  (.A(\V1/V3/V4/v4 [2]),
    .B(\V1/V3/V4/c3 ),
    .Z(\V1/V3/V4/A3/M3/s1 ));
 AND2_X1 \V1/V3/V4/A3/M3/M2/_0_  (.A1(\V1/V3/V4/A3/M3/s1 ),
    .A2(\V1/V3/V4/A3/c2 ),
    .ZN(\V1/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M3/M2/_1_  (.A(\V1/V3/V4/A3/M3/s1 ),
    .B(\V1/V3/V4/A3/c2 ),
    .Z(\V1/V3/v4 [6]));
 OR2_X1 \V1/V3/V4/A3/M3/_0_  (.A1(\V1/V3/V4/A3/M3/c1 ),
    .A2(\V1/V3/V4/A3/M3/c2 ),
    .ZN(\V1/V3/V4/A3/c3 ));
 AND2_X1 \V1/V3/V4/A3/M4/M1/_0_  (.A1(\V1/V3/V4/v4 [3]),
    .A2(net3),
    .ZN(\V1/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V3/V4/A3/M4/M1/_1_  (.A(\V1/V3/V4/v4 [3]),
    .B(net3),
    .Z(\V1/V3/V4/A3/M4/s1 ));
 AND2_X1 \V1/V3/V4/A3/M4/M2/_0_  (.A1(\V1/V3/V4/A3/M4/s1 ),
    .A2(\V1/V3/V4/A3/c3 ),
    .ZN(\V1/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V3/V4/A3/M4/M2/_1_  (.A(\V1/V3/V4/A3/M4/s1 ),
    .B(\V1/V3/V4/A3/c3 ),
    .Z(\V1/V3/v4 [7]));
 OR2_X1 \V1/V3/V4/A3/M4/_0_  (.A1(\V1/V3/V4/A3/M4/c1 ),
    .A2(\V1/V3/V4/A3/M4/c2 ),
    .ZN(\V1/V3/V4/overflow ));
 AND2_X1 \V1/V3/V4/V1/HA1/_0_  (.A1(\V1/V3/V4/V1/w2 ),
    .A2(\V1/V3/V4/V1/w1 ),
    .ZN(\V1/V3/V4/V1/w4 ));
 XOR2_X2 \V1/V3/V4/V1/HA1/_1_  (.A(\V1/V3/V4/V1/w2 ),
    .B(\V1/V3/V4/V1/w1 ),
    .Z(\V1/V3/v4 [1]));
 AND2_X1 \V1/V3/V4/V1/HA2/_0_  (.A1(\V1/V3/V4/V1/w4 ),
    .A2(\V1/V3/V4/V1/w3 ),
    .ZN(\V1/V3/V4/v1 [3]));
 XOR2_X2 \V1/V3/V4/V1/HA2/_1_  (.A(\V1/V3/V4/V1/w4 ),
    .B(\V1/V3/V4/V1/w3 ),
    .Z(\V1/V3/V4/v1 [2]));
 AND2_X1 \V1/V3/V4/V1/_0_  (.A1(A[4]),
    .A2(B[12]),
    .ZN(\V1/V3/v4 [0]));
 AND2_X1 \V1/V3/V4/V1/_1_  (.A1(A[4]),
    .A2(B[13]),
    .ZN(\V1/V3/V4/V1/w1 ));
 AND2_X1 \V1/V3/V4/V1/_2_  (.A1(B[12]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V1/w2 ));
 AND2_X1 \V1/V3/V4/V1/_3_  (.A1(B[13]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V1/w3 ));
 AND2_X1 \V1/V3/V4/V2/HA1/_0_  (.A1(\V1/V3/V4/V2/w2 ),
    .A2(\V1/V3/V4/V2/w1 ),
    .ZN(\V1/V3/V4/V2/w4 ));
 XOR2_X2 \V1/V3/V4/V2/HA1/_1_  (.A(\V1/V3/V4/V2/w2 ),
    .B(\V1/V3/V4/V2/w1 ),
    .Z(\V1/V3/V4/v2 [1]));
 AND2_X1 \V1/V3/V4/V2/HA2/_0_  (.A1(\V1/V3/V4/V2/w4 ),
    .A2(\V1/V3/V4/V2/w3 ),
    .ZN(\V1/V3/V4/v2 [3]));
 XOR2_X2 \V1/V3/V4/V2/HA2/_1_  (.A(\V1/V3/V4/V2/w4 ),
    .B(\V1/V3/V4/V2/w3 ),
    .Z(\V1/V3/V4/v2 [2]));
 AND2_X1 \V1/V3/V4/V2/_0_  (.A1(A[6]),
    .A2(B[12]),
    .ZN(\V1/V3/V4/v2 [0]));
 AND2_X1 \V1/V3/V4/V2/_1_  (.A1(A[6]),
    .A2(B[13]),
    .ZN(\V1/V3/V4/V2/w1 ));
 AND2_X1 \V1/V3/V4/V2/_2_  (.A1(B[12]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V2/w2 ));
 AND2_X1 \V1/V3/V4/V2/_3_  (.A1(B[13]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V2/w3 ));
 AND2_X1 \V1/V3/V4/V3/HA1/_0_  (.A1(\V1/V3/V4/V3/w2 ),
    .A2(\V1/V3/V4/V3/w1 ),
    .ZN(\V1/V3/V4/V3/w4 ));
 XOR2_X2 \V1/V3/V4/V3/HA1/_1_  (.A(\V1/V3/V4/V3/w2 ),
    .B(\V1/V3/V4/V3/w1 ),
    .Z(\V1/V3/V4/v3 [1]));
 AND2_X1 \V1/V3/V4/V3/HA2/_0_  (.A1(\V1/V3/V4/V3/w4 ),
    .A2(\V1/V3/V4/V3/w3 ),
    .ZN(\V1/V3/V4/v3 [3]));
 XOR2_X2 \V1/V3/V4/V3/HA2/_1_  (.A(\V1/V3/V4/V3/w4 ),
    .B(\V1/V3/V4/V3/w3 ),
    .Z(\V1/V3/V4/v3 [2]));
 AND2_X1 \V1/V3/V4/V3/_0_  (.A1(A[4]),
    .A2(B[14]),
    .ZN(\V1/V3/V4/v3 [0]));
 AND2_X1 \V1/V3/V4/V3/_1_  (.A1(A[4]),
    .A2(B[15]),
    .ZN(\V1/V3/V4/V3/w1 ));
 AND2_X1 \V1/V3/V4/V3/_2_  (.A1(B[14]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V3/w2 ));
 AND2_X1 \V1/V3/V4/V3/_3_  (.A1(B[15]),
    .A2(A[5]),
    .ZN(\V1/V3/V4/V3/w3 ));
 AND2_X1 \V1/V3/V4/V4/HA1/_0_  (.A1(\V1/V3/V4/V4/w2 ),
    .A2(\V1/V3/V4/V4/w1 ),
    .ZN(\V1/V3/V4/V4/w4 ));
 XOR2_X2 \V1/V3/V4/V4/HA1/_1_  (.A(\V1/V3/V4/V4/w2 ),
    .B(\V1/V3/V4/V4/w1 ),
    .Z(\V1/V3/V4/v4 [1]));
 AND2_X1 \V1/V3/V4/V4/HA2/_0_  (.A1(\V1/V3/V4/V4/w4 ),
    .A2(\V1/V3/V4/V4/w3 ),
    .ZN(\V1/V3/V4/v4 [3]));
 XOR2_X2 \V1/V3/V4/V4/HA2/_1_  (.A(\V1/V3/V4/V4/w4 ),
    .B(\V1/V3/V4/V4/w3 ),
    .Z(\V1/V3/V4/v4 [2]));
 AND2_X1 \V1/V3/V4/V4/_0_  (.A1(A[6]),
    .A2(B[14]),
    .ZN(\V1/V3/V4/v4 [0]));
 AND2_X1 \V1/V3/V4/V4/_1_  (.A1(A[6]),
    .A2(B[15]),
    .ZN(\V1/V3/V4/V4/w1 ));
 AND2_X1 \V1/V3/V4/V4/_2_  (.A1(B[14]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V4/w2 ));
 AND2_X1 \V1/V3/V4/V4/_3_  (.A1(B[15]),
    .A2(A[7]),
    .ZN(\V1/V3/V4/V4/w3 ));
 OR2_X1 \V1/V3/V4/_0_  (.A1(\V1/V3/V4/c1 ),
    .A2(\V1/V3/V4/c2 ),
    .ZN(\V1/V3/V4/c3 ));
 OR2_X1 \V1/V3/_0_  (.A1(\V1/V3/c1 ),
    .A2(\V1/V3/c2 ),
    .ZN(\V1/V3/c3 ));
 AND2_X1 \V1/V4/A1/A1/M1/M1/_0_  (.A1(\V1/V4/v2 [0]),
    .A2(\V1/V4/v3 [0]),
    .ZN(\V1/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M1/M1/_1_  (.A(\V1/V4/v2 [0]),
    .B(\V1/V4/v3 [0]),
    .Z(\V1/V4/A1/A1/M1/s1 ));
 AND2_X1 \V1/V4/A1/A1/M1/M2/_0_  (.A1(\V1/V4/A1/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M1/M2/_1_  (.A(\V1/V4/A1/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/V4/s1 [0]));
 OR2_X1 \V1/V4/A1/A1/M1/_0_  (.A1(\V1/V4/A1/A1/M1/c1 ),
    .A2(\V1/V4/A1/A1/M1/c2 ),
    .ZN(\V1/V4/A1/A1/c1 ));
 AND2_X1 \V1/V4/A1/A1/M2/M1/_0_  (.A1(\V1/V4/v2 [1]),
    .A2(\V1/V4/v3 [1]),
    .ZN(\V1/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M2/M1/_1_  (.A(\V1/V4/v2 [1]),
    .B(\V1/V4/v3 [1]),
    .Z(\V1/V4/A1/A1/M2/s1 ));
 AND2_X1 \V1/V4/A1/A1/M2/M2/_0_  (.A1(\V1/V4/A1/A1/M2/s1 ),
    .A2(\V1/V4/A1/A1/c1 ),
    .ZN(\V1/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M2/M2/_1_  (.A(\V1/V4/A1/A1/M2/s1 ),
    .B(\V1/V4/A1/A1/c1 ),
    .Z(\V1/V4/s1 [1]));
 OR2_X1 \V1/V4/A1/A1/M2/_0_  (.A1(\V1/V4/A1/A1/M2/c1 ),
    .A2(\V1/V4/A1/A1/M2/c2 ),
    .ZN(\V1/V4/A1/A1/c2 ));
 AND2_X1 \V1/V4/A1/A1/M3/M1/_0_  (.A1(\V1/V4/v2 [2]),
    .A2(\V1/V4/v3 [2]),
    .ZN(\V1/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M3/M1/_1_  (.A(\V1/V4/v2 [2]),
    .B(\V1/V4/v3 [2]),
    .Z(\V1/V4/A1/A1/M3/s1 ));
 AND2_X1 \V1/V4/A1/A1/M3/M2/_0_  (.A1(\V1/V4/A1/A1/M3/s1 ),
    .A2(\V1/V4/A1/A1/c2 ),
    .ZN(\V1/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M3/M2/_1_  (.A(\V1/V4/A1/A1/M3/s1 ),
    .B(\V1/V4/A1/A1/c2 ),
    .Z(\V1/V4/s1 [2]));
 OR2_X1 \V1/V4/A1/A1/M3/_0_  (.A1(\V1/V4/A1/A1/M3/c1 ),
    .A2(\V1/V4/A1/A1/M3/c2 ),
    .ZN(\V1/V4/A1/A1/c3 ));
 AND2_X1 \V1/V4/A1/A1/M4/M1/_0_  (.A1(\V1/V4/v2 [3]),
    .A2(\V1/V4/v3 [3]),
    .ZN(\V1/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A1/A1/M4/M1/_1_  (.A(\V1/V4/v2 [3]),
    .B(\V1/V4/v3 [3]),
    .Z(\V1/V4/A1/A1/M4/s1 ));
 AND2_X1 \V1/V4/A1/A1/M4/M2/_0_  (.A1(\V1/V4/A1/A1/M4/s1 ),
    .A2(\V1/V4/A1/A1/c3 ),
    .ZN(\V1/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A1/A1/M4/M2/_1_  (.A(\V1/V4/A1/A1/M4/s1 ),
    .B(\V1/V4/A1/A1/c3 ),
    .Z(\V1/V4/s1 [3]));
 OR2_X1 \V1/V4/A1/A1/M4/_0_  (.A1(\V1/V4/A1/A1/M4/c1 ),
    .A2(\V1/V4/A1/A1/M4/c2 ),
    .ZN(\V1/V4/A1/c1 ));
 AND2_X1 \V1/V4/A1/A2/M1/M1/_0_  (.A1(\V1/V4/v2 [4]),
    .A2(\V1/V4/v3 [4]),
    .ZN(\V1/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M1/M1/_1_  (.A(\V1/V4/v2 [4]),
    .B(\V1/V4/v3 [4]),
    .Z(\V1/V4/A1/A2/M1/s1 ));
 AND2_X1 \V1/V4/A1/A2/M1/M2/_0_  (.A1(\V1/V4/A1/A2/M1/s1 ),
    .A2(\V1/V4/A1/c1 ),
    .ZN(\V1/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M1/M2/_1_  (.A(\V1/V4/A1/A2/M1/s1 ),
    .B(\V1/V4/A1/c1 ),
    .Z(\V1/V4/s1 [4]));
 OR2_X1 \V1/V4/A1/A2/M1/_0_  (.A1(\V1/V4/A1/A2/M1/c1 ),
    .A2(\V1/V4/A1/A2/M1/c2 ),
    .ZN(\V1/V4/A1/A2/c1 ));
 AND2_X1 \V1/V4/A1/A2/M2/M1/_0_  (.A1(\V1/V4/v2 [5]),
    .A2(\V1/V4/v3 [5]),
    .ZN(\V1/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M2/M1/_1_  (.A(\V1/V4/v2 [5]),
    .B(\V1/V4/v3 [5]),
    .Z(\V1/V4/A1/A2/M2/s1 ));
 AND2_X1 \V1/V4/A1/A2/M2/M2/_0_  (.A1(\V1/V4/A1/A2/M2/s1 ),
    .A2(\V1/V4/A1/A2/c1 ),
    .ZN(\V1/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M2/M2/_1_  (.A(\V1/V4/A1/A2/M2/s1 ),
    .B(\V1/V4/A1/A2/c1 ),
    .Z(\V1/V4/s1 [5]));
 OR2_X1 \V1/V4/A1/A2/M2/_0_  (.A1(\V1/V4/A1/A2/M2/c1 ),
    .A2(\V1/V4/A1/A2/M2/c2 ),
    .ZN(\V1/V4/A1/A2/c2 ));
 AND2_X1 \V1/V4/A1/A2/M3/M1/_0_  (.A1(\V1/V4/v2 [6]),
    .A2(\V1/V4/v3 [6]),
    .ZN(\V1/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M3/M1/_1_  (.A(\V1/V4/v2 [6]),
    .B(\V1/V4/v3 [6]),
    .Z(\V1/V4/A1/A2/M3/s1 ));
 AND2_X1 \V1/V4/A1/A2/M3/M2/_0_  (.A1(\V1/V4/A1/A2/M3/s1 ),
    .A2(\V1/V4/A1/A2/c2 ),
    .ZN(\V1/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M3/M2/_1_  (.A(\V1/V4/A1/A2/M3/s1 ),
    .B(\V1/V4/A1/A2/c2 ),
    .Z(\V1/V4/s1 [6]));
 OR2_X1 \V1/V4/A1/A2/M3/_0_  (.A1(\V1/V4/A1/A2/M3/c1 ),
    .A2(\V1/V4/A1/A2/M3/c2 ),
    .ZN(\V1/V4/A1/A2/c3 ));
 AND2_X1 \V1/V4/A1/A2/M4/M1/_0_  (.A1(\V1/V4/v2 [7]),
    .A2(\V1/V4/v3 [7]),
    .ZN(\V1/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A1/A2/M4/M1/_1_  (.A(\V1/V4/v2 [7]),
    .B(\V1/V4/v3 [7]),
    .Z(\V1/V4/A1/A2/M4/s1 ));
 AND2_X1 \V1/V4/A1/A2/M4/M2/_0_  (.A1(\V1/V4/A1/A2/M4/s1 ),
    .A2(\V1/V4/A1/A2/c3 ),
    .ZN(\V1/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A1/A2/M4/M2/_1_  (.A(\V1/V4/A1/A2/M4/s1 ),
    .B(\V1/V4/A1/A2/c3 ),
    .Z(\V1/V4/s1 [7]));
 OR2_X1 \V1/V4/A1/A2/M4/_0_  (.A1(\V1/V4/A1/A2/M4/c1 ),
    .A2(\V1/V4/A1/A2/M4/c2 ),
    .ZN(\V1/V4/c1 ));
 AND2_X1 \V1/V4/A2/A1/M1/M1/_0_  (.A1(\V1/V4/s1 [0]),
    .A2(\V1/V4/v1 [4]),
    .ZN(\V1/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M1/M1/_1_  (.A(\V1/V4/s1 [0]),
    .B(\V1/V4/v1 [4]),
    .Z(\V1/V4/A2/A1/M1/s1 ));
 AND2_X1 \V1/V4/A2/A1/M1/M2/_0_  (.A1(\V1/V4/A2/A1/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M1/M2/_1_  (.A(\V1/V4/A2/A1/M1/s1 ),
    .B(net3),
    .Z(\V1/v4 [4]));
 OR2_X1 \V1/V4/A2/A1/M1/_0_  (.A1(\V1/V4/A2/A1/M1/c1 ),
    .A2(\V1/V4/A2/A1/M1/c2 ),
    .ZN(\V1/V4/A2/A1/c1 ));
 AND2_X1 \V1/V4/A2/A1/M2/M1/_0_  (.A1(\V1/V4/s1 [1]),
    .A2(\V1/V4/v1 [5]),
    .ZN(\V1/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M2/M1/_1_  (.A(\V1/V4/s1 [1]),
    .B(\V1/V4/v1 [5]),
    .Z(\V1/V4/A2/A1/M2/s1 ));
 AND2_X1 \V1/V4/A2/A1/M2/M2/_0_  (.A1(\V1/V4/A2/A1/M2/s1 ),
    .A2(\V1/V4/A2/A1/c1 ),
    .ZN(\V1/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M2/M2/_1_  (.A(\V1/V4/A2/A1/M2/s1 ),
    .B(\V1/V4/A2/A1/c1 ),
    .Z(\V1/v4 [5]));
 OR2_X1 \V1/V4/A2/A1/M2/_0_  (.A1(\V1/V4/A2/A1/M2/c1 ),
    .A2(\V1/V4/A2/A1/M2/c2 ),
    .ZN(\V1/V4/A2/A1/c2 ));
 AND2_X1 \V1/V4/A2/A1/M3/M1/_0_  (.A1(\V1/V4/s1 [2]),
    .A2(\V1/V4/v1 [6]),
    .ZN(\V1/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M3/M1/_1_  (.A(\V1/V4/s1 [2]),
    .B(\V1/V4/v1 [6]),
    .Z(\V1/V4/A2/A1/M3/s1 ));
 AND2_X1 \V1/V4/A2/A1/M3/M2/_0_  (.A1(\V1/V4/A2/A1/M3/s1 ),
    .A2(\V1/V4/A2/A1/c2 ),
    .ZN(\V1/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M3/M2/_1_  (.A(\V1/V4/A2/A1/M3/s1 ),
    .B(\V1/V4/A2/A1/c2 ),
    .Z(\V1/v4 [6]));
 OR2_X1 \V1/V4/A2/A1/M3/_0_  (.A1(\V1/V4/A2/A1/M3/c1 ),
    .A2(\V1/V4/A2/A1/M3/c2 ),
    .ZN(\V1/V4/A2/A1/c3 ));
 AND2_X1 \V1/V4/A2/A1/M4/M1/_0_  (.A1(\V1/V4/s1 [3]),
    .A2(\V1/V4/v1 [7]),
    .ZN(\V1/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A2/A1/M4/M1/_1_  (.A(\V1/V4/s1 [3]),
    .B(\V1/V4/v1 [7]),
    .Z(\V1/V4/A2/A1/M4/s1 ));
 AND2_X1 \V1/V4/A2/A1/M4/M2/_0_  (.A1(\V1/V4/A2/A1/M4/s1 ),
    .A2(\V1/V4/A2/A1/c3 ),
    .ZN(\V1/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A2/A1/M4/M2/_1_  (.A(\V1/V4/A2/A1/M4/s1 ),
    .B(\V1/V4/A2/A1/c3 ),
    .Z(\V1/v4 [7]));
 OR2_X1 \V1/V4/A2/A1/M4/_0_  (.A1(\V1/V4/A2/A1/M4/c1 ),
    .A2(\V1/V4/A2/A1/M4/c2 ),
    .ZN(\V1/V4/A2/c1 ));
 AND2_X1 \V1/V4/A2/A2/M1/M1/_0_  (.A1(\V1/V4/s1 [4]),
    .A2(net4),
    .ZN(\V1/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M1/M1/_1_  (.A(\V1/V4/s1 [4]),
    .B(net4),
    .Z(\V1/V4/A2/A2/M1/s1 ));
 AND2_X1 \V1/V4/A2/A2/M1/M2/_0_  (.A1(\V1/V4/A2/A2/M1/s1 ),
    .A2(\V1/V4/A2/c1 ),
    .ZN(\V1/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M1/M2/_1_  (.A(\V1/V4/A2/A2/M1/s1 ),
    .B(\V1/V4/A2/c1 ),
    .Z(\V1/V4/s2 [4]));
 OR2_X1 \V1/V4/A2/A2/M1/_0_  (.A1(\V1/V4/A2/A2/M1/c1 ),
    .A2(\V1/V4/A2/A2/M1/c2 ),
    .ZN(\V1/V4/A2/A2/c1 ));
 AND2_X1 \V1/V4/A2/A2/M2/M1/_0_  (.A1(\V1/V4/s1 [5]),
    .A2(net4),
    .ZN(\V1/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M2/M1/_1_  (.A(\V1/V4/s1 [5]),
    .B(net4),
    .Z(\V1/V4/A2/A2/M2/s1 ));
 AND2_X1 \V1/V4/A2/A2/M2/M2/_0_  (.A1(\V1/V4/A2/A2/M2/s1 ),
    .A2(\V1/V4/A2/A2/c1 ),
    .ZN(\V1/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M2/M2/_1_  (.A(\V1/V4/A2/A2/M2/s1 ),
    .B(\V1/V4/A2/A2/c1 ),
    .Z(\V1/V4/s2 [5]));
 OR2_X1 \V1/V4/A2/A2/M2/_0_  (.A1(\V1/V4/A2/A2/M2/c1 ),
    .A2(\V1/V4/A2/A2/M2/c2 ),
    .ZN(\V1/V4/A2/A2/c2 ));
 AND2_X1 \V1/V4/A2/A2/M3/M1/_0_  (.A1(\V1/V4/s1 [6]),
    .A2(net4),
    .ZN(\V1/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M3/M1/_1_  (.A(\V1/V4/s1 [6]),
    .B(net4),
    .Z(\V1/V4/A2/A2/M3/s1 ));
 AND2_X1 \V1/V4/A2/A2/M3/M2/_0_  (.A1(\V1/V4/A2/A2/M3/s1 ),
    .A2(\V1/V4/A2/A2/c2 ),
    .ZN(\V1/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M3/M2/_1_  (.A(\V1/V4/A2/A2/M3/s1 ),
    .B(\V1/V4/A2/A2/c2 ),
    .Z(\V1/V4/s2 [6]));
 OR2_X1 \V1/V4/A2/A2/M3/_0_  (.A1(\V1/V4/A2/A2/M3/c1 ),
    .A2(\V1/V4/A2/A2/M3/c2 ),
    .ZN(\V1/V4/A2/A2/c3 ));
 AND2_X1 \V1/V4/A2/A2/M4/M1/_0_  (.A1(\V1/V4/s1 [7]),
    .A2(net4),
    .ZN(\V1/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A2/A2/M4/M1/_1_  (.A(\V1/V4/s1 [7]),
    .B(net4),
    .Z(\V1/V4/A2/A2/M4/s1 ));
 AND2_X1 \V1/V4/A2/A2/M4/M2/_0_  (.A1(\V1/V4/A2/A2/M4/s1 ),
    .A2(\V1/V4/A2/A2/c3 ),
    .ZN(\V1/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A2/A2/M4/M2/_1_  (.A(\V1/V4/A2/A2/M4/s1 ),
    .B(\V1/V4/A2/A2/c3 ),
    .Z(\V1/V4/s2 [7]));
 OR2_X1 \V1/V4/A2/A2/M4/_0_  (.A1(\V1/V4/A2/A2/M4/c1 ),
    .A2(\V1/V4/A2/A2/M4/c2 ),
    .ZN(\V1/V4/c2 ));
 AND2_X1 \V1/V4/A3/A1/M1/M1/_0_  (.A1(\V1/V4/v4 [0]),
    .A2(\V1/V4/s2 [4]),
    .ZN(\V1/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M1/M1/_1_  (.A(\V1/V4/v4 [0]),
    .B(\V1/V4/s2 [4]),
    .Z(\V1/V4/A3/A1/M1/s1 ));
 AND2_X1 \V1/V4/A3/A1/M1/M2/_0_  (.A1(\V1/V4/A3/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M1/M2/_1_  (.A(\V1/V4/A3/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/v4 [8]));
 OR2_X1 \V1/V4/A3/A1/M1/_0_  (.A1(\V1/V4/A3/A1/M1/c1 ),
    .A2(\V1/V4/A3/A1/M1/c2 ),
    .ZN(\V1/V4/A3/A1/c1 ));
 AND2_X1 \V1/V4/A3/A1/M2/M1/_0_  (.A1(\V1/V4/v4 [1]),
    .A2(\V1/V4/s2 [5]),
    .ZN(\V1/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M2/M1/_1_  (.A(\V1/V4/v4 [1]),
    .B(\V1/V4/s2 [5]),
    .Z(\V1/V4/A3/A1/M2/s1 ));
 AND2_X1 \V1/V4/A3/A1/M2/M2/_0_  (.A1(\V1/V4/A3/A1/M2/s1 ),
    .A2(\V1/V4/A3/A1/c1 ),
    .ZN(\V1/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M2/M2/_1_  (.A(\V1/V4/A3/A1/M2/s1 ),
    .B(\V1/V4/A3/A1/c1 ),
    .Z(\V1/v4 [9]));
 OR2_X1 \V1/V4/A3/A1/M2/_0_  (.A1(\V1/V4/A3/A1/M2/c1 ),
    .A2(\V1/V4/A3/A1/M2/c2 ),
    .ZN(\V1/V4/A3/A1/c2 ));
 AND2_X1 \V1/V4/A3/A1/M3/M1/_0_  (.A1(\V1/V4/v4 [2]),
    .A2(\V1/V4/s2 [6]),
    .ZN(\V1/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M3/M1/_1_  (.A(\V1/V4/v4 [2]),
    .B(\V1/V4/s2 [6]),
    .Z(\V1/V4/A3/A1/M3/s1 ));
 AND2_X1 \V1/V4/A3/A1/M3/M2/_0_  (.A1(\V1/V4/A3/A1/M3/s1 ),
    .A2(\V1/V4/A3/A1/c2 ),
    .ZN(\V1/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M3/M2/_1_  (.A(\V1/V4/A3/A1/M3/s1 ),
    .B(\V1/V4/A3/A1/c2 ),
    .Z(\V1/v4 [10]));
 OR2_X1 \V1/V4/A3/A1/M3/_0_  (.A1(\V1/V4/A3/A1/M3/c1 ),
    .A2(\V1/V4/A3/A1/M3/c2 ),
    .ZN(\V1/V4/A3/A1/c3 ));
 AND2_X1 \V1/V4/A3/A1/M4/M1/_0_  (.A1(\V1/V4/v4 [3]),
    .A2(\V1/V4/s2 [7]),
    .ZN(\V1/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V1/V4/A3/A1/M4/M1/_1_  (.A(\V1/V4/v4 [3]),
    .B(\V1/V4/s2 [7]),
    .Z(\V1/V4/A3/A1/M4/s1 ));
 AND2_X1 \V1/V4/A3/A1/M4/M2/_0_  (.A1(\V1/V4/A3/A1/M4/s1 ),
    .A2(\V1/V4/A3/A1/c3 ),
    .ZN(\V1/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V1/V4/A3/A1/M4/M2/_1_  (.A(\V1/V4/A3/A1/M4/s1 ),
    .B(\V1/V4/A3/A1/c3 ),
    .Z(\V1/v4 [11]));
 OR2_X1 \V1/V4/A3/A1/M4/_0_  (.A1(\V1/V4/A3/A1/M4/c1 ),
    .A2(\V1/V4/A3/A1/M4/c2 ),
    .ZN(\V1/V4/A3/c1 ));
 AND2_X1 \V1/V4/A3/A2/M1/M1/_0_  (.A1(\V1/V4/v4 [4]),
    .A2(\V1/V4/c3 ),
    .ZN(\V1/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M1/M1/_1_  (.A(\V1/V4/v4 [4]),
    .B(\V1/V4/c3 ),
    .Z(\V1/V4/A3/A2/M1/s1 ));
 AND2_X1 \V1/V4/A3/A2/M1/M2/_0_  (.A1(\V1/V4/A3/A2/M1/s1 ),
    .A2(\V1/V4/A3/c1 ),
    .ZN(\V1/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M1/M2/_1_  (.A(\V1/V4/A3/A2/M1/s1 ),
    .B(\V1/V4/A3/c1 ),
    .Z(\V1/v4 [12]));
 OR2_X1 \V1/V4/A3/A2/M1/_0_  (.A1(\V1/V4/A3/A2/M1/c1 ),
    .A2(\V1/V4/A3/A2/M1/c2 ),
    .ZN(\V1/V4/A3/A2/c1 ));
 AND2_X1 \V1/V4/A3/A2/M2/M1/_0_  (.A1(\V1/V4/v4 [5]),
    .A2(net6),
    .ZN(\V1/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M2/M1/_1_  (.A(\V1/V4/v4 [5]),
    .B(net6),
    .Z(\V1/V4/A3/A2/M2/s1 ));
 AND2_X1 \V1/V4/A3/A2/M2/M2/_0_  (.A1(\V1/V4/A3/A2/M2/s1 ),
    .A2(\V1/V4/A3/A2/c1 ),
    .ZN(\V1/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M2/M2/_1_  (.A(\V1/V4/A3/A2/M2/s1 ),
    .B(\V1/V4/A3/A2/c1 ),
    .Z(\V1/v4 [13]));
 OR2_X1 \V1/V4/A3/A2/M2/_0_  (.A1(\V1/V4/A3/A2/M2/c1 ),
    .A2(\V1/V4/A3/A2/M2/c2 ),
    .ZN(\V1/V4/A3/A2/c2 ));
 AND2_X1 \V1/V4/A3/A2/M3/M1/_0_  (.A1(\V1/V4/v4 [6]),
    .A2(net6),
    .ZN(\V1/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M3/M1/_1_  (.A(\V1/V4/v4 [6]),
    .B(net6),
    .Z(\V1/V4/A3/A2/M3/s1 ));
 AND2_X1 \V1/V4/A3/A2/M3/M2/_0_  (.A1(\V1/V4/A3/A2/M3/s1 ),
    .A2(\V1/V4/A3/A2/c2 ),
    .ZN(\V1/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M3/M2/_1_  (.A(\V1/V4/A3/A2/M3/s1 ),
    .B(\V1/V4/A3/A2/c2 ),
    .Z(\V1/v4 [14]));
 OR2_X1 \V1/V4/A3/A2/M3/_0_  (.A1(\V1/V4/A3/A2/M3/c1 ),
    .A2(\V1/V4/A3/A2/M3/c2 ),
    .ZN(\V1/V4/A3/A2/c3 ));
 AND2_X1 \V1/V4/A3/A2/M4/M1/_0_  (.A1(\V1/V4/v4 [7]),
    .A2(net6),
    .ZN(\V1/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V1/V4/A3/A2/M4/M1/_1_  (.A(\V1/V4/v4 [7]),
    .B(net6),
    .Z(\V1/V4/A3/A2/M4/s1 ));
 AND2_X1 \V1/V4/A3/A2/M4/M2/_0_  (.A1(\V1/V4/A3/A2/M4/s1 ),
    .A2(\V1/V4/A3/A2/c3 ),
    .ZN(\V1/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V1/V4/A3/A2/M4/M2/_1_  (.A(\V1/V4/A3/A2/M4/s1 ),
    .B(\V1/V4/A3/A2/c3 ),
    .Z(\V1/v4 [15]));
 OR2_X1 \V1/V4/A3/A2/M4/_0_  (.A1(\V1/V4/A3/A2/M4/c1 ),
    .A2(\V1/V4/A3/A2/M4/c2 ),
    .ZN(\V1/V4/overflow ));
 AND2_X1 \V1/V4/V1/A1/M1/M1/_0_  (.A1(\V1/V4/V1/v2 [0]),
    .A2(\V1/V4/V1/v3 [0]),
    .ZN(\V1/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M1/M1/_1_  (.A(\V1/V4/V1/v2 [0]),
    .B(\V1/V4/V1/v3 [0]),
    .Z(\V1/V4/V1/A1/M1/s1 ));
 AND2_X1 \V1/V4/V1/A1/M1/M2/_0_  (.A1(\V1/V4/V1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M1/M2/_1_  (.A(\V1/V4/V1/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/V1/s1 [0]));
 OR2_X1 \V1/V4/V1/A1/M1/_0_  (.A1(\V1/V4/V1/A1/M1/c1 ),
    .A2(\V1/V4/V1/A1/M1/c2 ),
    .ZN(\V1/V4/V1/A1/c1 ));
 AND2_X1 \V1/V4/V1/A1/M2/M1/_0_  (.A1(\V1/V4/V1/v2 [1]),
    .A2(\V1/V4/V1/v3 [1]),
    .ZN(\V1/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M2/M1/_1_  (.A(\V1/V4/V1/v2 [1]),
    .B(\V1/V4/V1/v3 [1]),
    .Z(\V1/V4/V1/A1/M2/s1 ));
 AND2_X1 \V1/V4/V1/A1/M2/M2/_0_  (.A1(\V1/V4/V1/A1/M2/s1 ),
    .A2(\V1/V4/V1/A1/c1 ),
    .ZN(\V1/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M2/M2/_1_  (.A(\V1/V4/V1/A1/M2/s1 ),
    .B(\V1/V4/V1/A1/c1 ),
    .Z(\V1/V4/V1/s1 [1]));
 OR2_X1 \V1/V4/V1/A1/M2/_0_  (.A1(\V1/V4/V1/A1/M2/c1 ),
    .A2(\V1/V4/V1/A1/M2/c2 ),
    .ZN(\V1/V4/V1/A1/c2 ));
 AND2_X1 \V1/V4/V1/A1/M3/M1/_0_  (.A1(\V1/V4/V1/v2 [2]),
    .A2(\V1/V4/V1/v3 [2]),
    .ZN(\V1/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M3/M1/_1_  (.A(\V1/V4/V1/v2 [2]),
    .B(\V1/V4/V1/v3 [2]),
    .Z(\V1/V4/V1/A1/M3/s1 ));
 AND2_X1 \V1/V4/V1/A1/M3/M2/_0_  (.A1(\V1/V4/V1/A1/M3/s1 ),
    .A2(\V1/V4/V1/A1/c2 ),
    .ZN(\V1/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M3/M2/_1_  (.A(\V1/V4/V1/A1/M3/s1 ),
    .B(\V1/V4/V1/A1/c2 ),
    .Z(\V1/V4/V1/s1 [2]));
 OR2_X1 \V1/V4/V1/A1/M3/_0_  (.A1(\V1/V4/V1/A1/M3/c1 ),
    .A2(\V1/V4/V1/A1/M3/c2 ),
    .ZN(\V1/V4/V1/A1/c3 ));
 AND2_X1 \V1/V4/V1/A1/M4/M1/_0_  (.A1(\V1/V4/V1/v2 [3]),
    .A2(\V1/V4/V1/v3 [3]),
    .ZN(\V1/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A1/M4/M1/_1_  (.A(\V1/V4/V1/v2 [3]),
    .B(\V1/V4/V1/v3 [3]),
    .Z(\V1/V4/V1/A1/M4/s1 ));
 AND2_X1 \V1/V4/V1/A1/M4/M2/_0_  (.A1(\V1/V4/V1/A1/M4/s1 ),
    .A2(\V1/V4/V1/A1/c3 ),
    .ZN(\V1/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A1/M4/M2/_1_  (.A(\V1/V4/V1/A1/M4/s1 ),
    .B(\V1/V4/V1/A1/c3 ),
    .Z(\V1/V4/V1/s1 [3]));
 OR2_X1 \V1/V4/V1/A1/M4/_0_  (.A1(\V1/V4/V1/A1/M4/c1 ),
    .A2(\V1/V4/V1/A1/M4/c2 ),
    .ZN(\V1/V4/V1/c1 ));
 AND2_X1 \V1/V4/V1/A2/M1/M1/_0_  (.A1(\V1/V4/V1/s1 [0]),
    .A2(\V1/V4/V1/v1 [2]),
    .ZN(\V1/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M1/M1/_1_  (.A(\V1/V4/V1/s1 [0]),
    .B(\V1/V4/V1/v1 [2]),
    .Z(\V1/V4/V1/A2/M1/s1 ));
 AND2_X1 \V1/V4/V1/A2/M1/M2/_0_  (.A1(\V1/V4/V1/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M1/M2/_1_  (.A(\V1/V4/V1/A2/M1/s1 ),
    .B(net5),
    .Z(\V1/v4 [2]));
 OR2_X1 \V1/V4/V1/A2/M1/_0_  (.A1(\V1/V4/V1/A2/M1/c1 ),
    .A2(\V1/V4/V1/A2/M1/c2 ),
    .ZN(\V1/V4/V1/A2/c1 ));
 AND2_X1 \V1/V4/V1/A2/M2/M1/_0_  (.A1(\V1/V4/V1/s1 [1]),
    .A2(\V1/V4/V1/v1 [3]),
    .ZN(\V1/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M2/M1/_1_  (.A(\V1/V4/V1/s1 [1]),
    .B(\V1/V4/V1/v1 [3]),
    .Z(\V1/V4/V1/A2/M2/s1 ));
 AND2_X1 \V1/V4/V1/A2/M2/M2/_0_  (.A1(\V1/V4/V1/A2/M2/s1 ),
    .A2(\V1/V4/V1/A2/c1 ),
    .ZN(\V1/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M2/M2/_1_  (.A(\V1/V4/V1/A2/M2/s1 ),
    .B(\V1/V4/V1/A2/c1 ),
    .Z(\V1/v4 [3]));
 OR2_X1 \V1/V4/V1/A2/M2/_0_  (.A1(\V1/V4/V1/A2/M2/c1 ),
    .A2(\V1/V4/V1/A2/M2/c2 ),
    .ZN(\V1/V4/V1/A2/c2 ));
 AND2_X1 \V1/V4/V1/A2/M3/M1/_0_  (.A1(\V1/V4/V1/s1 [2]),
    .A2(net5),
    .ZN(\V1/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M3/M1/_1_  (.A(\V1/V4/V1/s1 [2]),
    .B(net5),
    .Z(\V1/V4/V1/A2/M3/s1 ));
 AND2_X1 \V1/V4/V1/A2/M3/M2/_0_  (.A1(\V1/V4/V1/A2/M3/s1 ),
    .A2(\V1/V4/V1/A2/c2 ),
    .ZN(\V1/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M3/M2/_1_  (.A(\V1/V4/V1/A2/M3/s1 ),
    .B(\V1/V4/V1/A2/c2 ),
    .Z(\V1/V4/V1/s2 [2]));
 OR2_X1 \V1/V4/V1/A2/M3/_0_  (.A1(\V1/V4/V1/A2/M3/c1 ),
    .A2(\V1/V4/V1/A2/M3/c2 ),
    .ZN(\V1/V4/V1/A2/c3 ));
 AND2_X1 \V1/V4/V1/A2/M4/M1/_0_  (.A1(\V1/V4/V1/s1 [3]),
    .A2(net5),
    .ZN(\V1/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A2/M4/M1/_1_  (.A(\V1/V4/V1/s1 [3]),
    .B(net5),
    .Z(\V1/V4/V1/A2/M4/s1 ));
 AND2_X1 \V1/V4/V1/A2/M4/M2/_0_  (.A1(\V1/V4/V1/A2/M4/s1 ),
    .A2(\V1/V4/V1/A2/c3 ),
    .ZN(\V1/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A2/M4/M2/_1_  (.A(\V1/V4/V1/A2/M4/s1 ),
    .B(\V1/V4/V1/A2/c3 ),
    .Z(\V1/V4/V1/s2 [3]));
 OR2_X1 \V1/V4/V1/A2/M4/_0_  (.A1(\V1/V4/V1/A2/M4/c1 ),
    .A2(\V1/V4/V1/A2/M4/c2 ),
    .ZN(\V1/V4/V1/c2 ));
 AND2_X1 \V1/V4/V1/A3/M1/M1/_0_  (.A1(\V1/V4/V1/v4 [0]),
    .A2(\V1/V4/V1/s2 [2]),
    .ZN(\V1/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M1/M1/_1_  (.A(\V1/V4/V1/v4 [0]),
    .B(\V1/V4/V1/s2 [2]),
    .Z(\V1/V4/V1/A3/M1/s1 ));
 AND2_X1 \V1/V4/V1/A3/M1/M2/_0_  (.A1(\V1/V4/V1/A3/M1/s1 ),
    .A2(net3),
    .ZN(\V1/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M1/M2/_1_  (.A(\V1/V4/V1/A3/M1/s1 ),
    .B(net3),
    .Z(\V1/V4/v1 [4]));
 OR2_X1 \V1/V4/V1/A3/M1/_0_  (.A1(\V1/V4/V1/A3/M1/c1 ),
    .A2(\V1/V4/V1/A3/M1/c2 ),
    .ZN(\V1/V4/V1/A3/c1 ));
 AND2_X1 \V1/V4/V1/A3/M2/M1/_0_  (.A1(\V1/V4/V1/v4 [1]),
    .A2(\V1/V4/V1/s2 [3]),
    .ZN(\V1/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M2/M1/_1_  (.A(\V1/V4/V1/v4 [1]),
    .B(\V1/V4/V1/s2 [3]),
    .Z(\V1/V4/V1/A3/M2/s1 ));
 AND2_X1 \V1/V4/V1/A3/M2/M2/_0_  (.A1(\V1/V4/V1/A3/M2/s1 ),
    .A2(\V1/V4/V1/A3/c1 ),
    .ZN(\V1/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M2/M2/_1_  (.A(\V1/V4/V1/A3/M2/s1 ),
    .B(\V1/V4/V1/A3/c1 ),
    .Z(\V1/V4/v1 [5]));
 OR2_X1 \V1/V4/V1/A3/M2/_0_  (.A1(\V1/V4/V1/A3/M2/c1 ),
    .A2(\V1/V4/V1/A3/M2/c2 ),
    .ZN(\V1/V4/V1/A3/c2 ));
 AND2_X1 \V1/V4/V1/A3/M3/M1/_0_  (.A1(\V1/V4/V1/v4 [2]),
    .A2(\V1/V4/V1/c3 ),
    .ZN(\V1/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M3/M1/_1_  (.A(\V1/V4/V1/v4 [2]),
    .B(\V1/V4/V1/c3 ),
    .Z(\V1/V4/V1/A3/M3/s1 ));
 AND2_X1 \V1/V4/V1/A3/M3/M2/_0_  (.A1(\V1/V4/V1/A3/M3/s1 ),
    .A2(\V1/V4/V1/A3/c2 ),
    .ZN(\V1/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M3/M2/_1_  (.A(\V1/V4/V1/A3/M3/s1 ),
    .B(\V1/V4/V1/A3/c2 ),
    .Z(\V1/V4/v1 [6]));
 OR2_X1 \V1/V4/V1/A3/M3/_0_  (.A1(\V1/V4/V1/A3/M3/c1 ),
    .A2(\V1/V4/V1/A3/M3/c2 ),
    .ZN(\V1/V4/V1/A3/c3 ));
 AND2_X1 \V1/V4/V1/A3/M4/M1/_0_  (.A1(\V1/V4/V1/v4 [3]),
    .A2(net5),
    .ZN(\V1/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V1/A3/M4/M1/_1_  (.A(\V1/V4/V1/v4 [3]),
    .B(net5),
    .Z(\V1/V4/V1/A3/M4/s1 ));
 AND2_X1 \V1/V4/V1/A3/M4/M2/_0_  (.A1(\V1/V4/V1/A3/M4/s1 ),
    .A2(\V1/V4/V1/A3/c3 ),
    .ZN(\V1/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V1/A3/M4/M2/_1_  (.A(\V1/V4/V1/A3/M4/s1 ),
    .B(\V1/V4/V1/A3/c3 ),
    .Z(\V1/V4/v1 [7]));
 OR2_X1 \V1/V4/V1/A3/M4/_0_  (.A1(\V1/V4/V1/A3/M4/c1 ),
    .A2(\V1/V4/V1/A3/M4/c2 ),
    .ZN(\V1/V4/V1/overflow ));
 AND2_X1 \V1/V4/V1/V1/HA1/_0_  (.A1(\V1/V4/V1/V1/w2 ),
    .A2(\V1/V4/V1/V1/w1 ),
    .ZN(\V1/V4/V1/V1/w4 ));
 XOR2_X2 \V1/V4/V1/V1/HA1/_1_  (.A(\V1/V4/V1/V1/w2 ),
    .B(\V1/V4/V1/V1/w1 ),
    .Z(\V1/v4 [1]));
 AND2_X1 \V1/V4/V1/V1/HA2/_0_  (.A1(\V1/V4/V1/V1/w4 ),
    .A2(\V1/V4/V1/V1/w3 ),
    .ZN(\V1/V4/V1/v1 [3]));
 XOR2_X2 \V1/V4/V1/V1/HA2/_1_  (.A(\V1/V4/V1/V1/w4 ),
    .B(\V1/V4/V1/V1/w3 ),
    .Z(\V1/V4/V1/v1 [2]));
 AND2_X1 \V1/V4/V1/V1/_0_  (.A1(net25),
    .A2(net12),
    .ZN(\V1/v4 [0]));
 AND2_X1 \V1/V4/V1/V1/_1_  (.A1(net25),
    .A2(net11),
    .ZN(\V1/V4/V1/V1/w1 ));
 AND2_X1 \V1/V4/V1/V1/_2_  (.A1(net12),
    .A2(net24),
    .ZN(\V1/V4/V1/V1/w2 ));
 AND2_X1 \V1/V4/V1/V1/_3_  (.A1(net11),
    .A2(net24),
    .ZN(\V1/V4/V1/V1/w3 ));
 AND2_X1 \V1/V4/V1/V2/HA1/_0_  (.A1(\V1/V4/V1/V2/w2 ),
    .A2(\V1/V4/V1/V2/w1 ),
    .ZN(\V1/V4/V1/V2/w4 ));
 XOR2_X2 \V1/V4/V1/V2/HA1/_1_  (.A(\V1/V4/V1/V2/w2 ),
    .B(\V1/V4/V1/V2/w1 ),
    .Z(\V1/V4/V1/v2 [1]));
 AND2_X1 \V1/V4/V1/V2/HA2/_0_  (.A1(\V1/V4/V1/V2/w4 ),
    .A2(\V1/V4/V1/V2/w3 ),
    .ZN(\V1/V4/V1/v2 [3]));
 XOR2_X2 \V1/V4/V1/V2/HA2/_1_  (.A(\V1/V4/V1/V2/w4 ),
    .B(\V1/V4/V1/V2/w3 ),
    .Z(\V1/V4/V1/v2 [2]));
 AND2_X1 \V1/V4/V1/V2/_0_  (.A1(net47),
    .A2(net12),
    .ZN(\V1/V4/V1/v2 [0]));
 AND2_X1 \V1/V4/V1/V2/_1_  (.A1(net47),
    .A2(net11),
    .ZN(\V1/V4/V1/V2/w1 ));
 AND2_X1 \V1/V4/V1/V2/_2_  (.A1(net12),
    .A2(net46),
    .ZN(\V1/V4/V1/V2/w2 ));
 AND2_X1 \V1/V4/V1/V2/_3_  (.A1(net11),
    .A2(net46),
    .ZN(\V1/V4/V1/V2/w3 ));
 AND2_X1 \V1/V4/V1/V3/HA1/_0_  (.A1(\V1/V4/V1/V3/w2 ),
    .A2(\V1/V4/V1/V3/w1 ),
    .ZN(\V1/V4/V1/V3/w4 ));
 XOR2_X2 \V1/V4/V1/V3/HA1/_1_  (.A(\V1/V4/V1/V3/w2 ),
    .B(\V1/V4/V1/V3/w1 ),
    .Z(\V1/V4/V1/v3 [1]));
 AND2_X1 \V1/V4/V1/V3/HA2/_0_  (.A1(\V1/V4/V1/V3/w4 ),
    .A2(\V1/V4/V1/V3/w3 ),
    .ZN(\V1/V4/V1/v3 [3]));
 XOR2_X2 \V1/V4/V1/V3/HA2/_1_  (.A(\V1/V4/V1/V3/w4 ),
    .B(\V1/V4/V1/V3/w3 ),
    .Z(\V1/V4/V1/v3 [2]));
 AND2_X1 \V1/V4/V1/V3/_0_  (.A1(net25),
    .A2(B[10]),
    .ZN(\V1/V4/V1/v3 [0]));
 AND2_X1 \V1/V4/V1/V3/_1_  (.A1(net25),
    .A2(B[11]),
    .ZN(\V1/V4/V1/V3/w1 ));
 AND2_X1 \V1/V4/V1/V3/_2_  (.A1(B[10]),
    .A2(net24),
    .ZN(\V1/V4/V1/V3/w2 ));
 AND2_X1 \V1/V4/V1/V3/_3_  (.A1(B[11]),
    .A2(net24),
    .ZN(\V1/V4/V1/V3/w3 ));
 AND2_X1 \V1/V4/V1/V4/HA1/_0_  (.A1(\V1/V4/V1/V4/w2 ),
    .A2(\V1/V4/V1/V4/w1 ),
    .ZN(\V1/V4/V1/V4/w4 ));
 XOR2_X2 \V1/V4/V1/V4/HA1/_1_  (.A(\V1/V4/V1/V4/w2 ),
    .B(\V1/V4/V1/V4/w1 ),
    .Z(\V1/V4/V1/v4 [1]));
 AND2_X1 \V1/V4/V1/V4/HA2/_0_  (.A1(\V1/V4/V1/V4/w4 ),
    .A2(\V1/V4/V1/V4/w3 ),
    .ZN(\V1/V4/V1/v4 [3]));
 XOR2_X2 \V1/V4/V1/V4/HA2/_1_  (.A(\V1/V4/V1/V4/w4 ),
    .B(\V1/V4/V1/V4/w3 ),
    .Z(\V1/V4/V1/v4 [2]));
 AND2_X1 \V1/V4/V1/V4/_0_  (.A1(net47),
    .A2(B[10]),
    .ZN(\V1/V4/V1/v4 [0]));
 AND2_X1 \V1/V4/V1/V4/_1_  (.A1(net47),
    .A2(B[11]),
    .ZN(\V1/V4/V1/V4/w1 ));
 AND2_X1 \V1/V4/V1/V4/_2_  (.A1(B[10]),
    .A2(net46),
    .ZN(\V1/V4/V1/V4/w2 ));
 AND2_X1 \V1/V4/V1/V4/_3_  (.A1(B[11]),
    .A2(net46),
    .ZN(\V1/V4/V1/V4/w3 ));
 OR2_X1 \V1/V4/V1/_0_  (.A1(\V1/V4/V1/c1 ),
    .A2(\V1/V4/V1/c2 ),
    .ZN(\V1/V4/V1/c3 ));
 AND2_X1 \V1/V4/V2/A1/M1/M1/_0_  (.A1(\V1/V4/V2/v2 [0]),
    .A2(\V1/V4/V2/v3 [0]),
    .ZN(\V1/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M1/M1/_1_  (.A(\V1/V4/V2/v2 [0]),
    .B(\V1/V4/V2/v3 [0]),
    .Z(\V1/V4/V2/A1/M1/s1 ));
 AND2_X1 \V1/V4/V2/A1/M1/M2/_0_  (.A1(\V1/V4/V2/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M1/M2/_1_  (.A(\V1/V4/V2/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/V2/s1 [0]));
 OR2_X1 \V1/V4/V2/A1/M1/_0_  (.A1(\V1/V4/V2/A1/M1/c1 ),
    .A2(\V1/V4/V2/A1/M1/c2 ),
    .ZN(\V1/V4/V2/A1/c1 ));
 AND2_X1 \V1/V4/V2/A1/M2/M1/_0_  (.A1(\V1/V4/V2/v2 [1]),
    .A2(\V1/V4/V2/v3 [1]),
    .ZN(\V1/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M2/M1/_1_  (.A(\V1/V4/V2/v2 [1]),
    .B(\V1/V4/V2/v3 [1]),
    .Z(\V1/V4/V2/A1/M2/s1 ));
 AND2_X1 \V1/V4/V2/A1/M2/M2/_0_  (.A1(\V1/V4/V2/A1/M2/s1 ),
    .A2(\V1/V4/V2/A1/c1 ),
    .ZN(\V1/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M2/M2/_1_  (.A(\V1/V4/V2/A1/M2/s1 ),
    .B(\V1/V4/V2/A1/c1 ),
    .Z(\V1/V4/V2/s1 [1]));
 OR2_X1 \V1/V4/V2/A1/M2/_0_  (.A1(\V1/V4/V2/A1/M2/c1 ),
    .A2(\V1/V4/V2/A1/M2/c2 ),
    .ZN(\V1/V4/V2/A1/c2 ));
 AND2_X1 \V1/V4/V2/A1/M3/M1/_0_  (.A1(\V1/V4/V2/v2 [2]),
    .A2(\V1/V4/V2/v3 [2]),
    .ZN(\V1/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M3/M1/_1_  (.A(\V1/V4/V2/v2 [2]),
    .B(\V1/V4/V2/v3 [2]),
    .Z(\V1/V4/V2/A1/M3/s1 ));
 AND2_X1 \V1/V4/V2/A1/M3/M2/_0_  (.A1(\V1/V4/V2/A1/M3/s1 ),
    .A2(\V1/V4/V2/A1/c2 ),
    .ZN(\V1/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M3/M2/_1_  (.A(\V1/V4/V2/A1/M3/s1 ),
    .B(\V1/V4/V2/A1/c2 ),
    .Z(\V1/V4/V2/s1 [2]));
 OR2_X1 \V1/V4/V2/A1/M3/_0_  (.A1(\V1/V4/V2/A1/M3/c1 ),
    .A2(\V1/V4/V2/A1/M3/c2 ),
    .ZN(\V1/V4/V2/A1/c3 ));
 AND2_X1 \V1/V4/V2/A1/M4/M1/_0_  (.A1(\V1/V4/V2/v2 [3]),
    .A2(\V1/V4/V2/v3 [3]),
    .ZN(\V1/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A1/M4/M1/_1_  (.A(\V1/V4/V2/v2 [3]),
    .B(\V1/V4/V2/v3 [3]),
    .Z(\V1/V4/V2/A1/M4/s1 ));
 AND2_X1 \V1/V4/V2/A1/M4/M2/_0_  (.A1(\V1/V4/V2/A1/M4/s1 ),
    .A2(\V1/V4/V2/A1/c3 ),
    .ZN(\V1/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A1/M4/M2/_1_  (.A(\V1/V4/V2/A1/M4/s1 ),
    .B(\V1/V4/V2/A1/c3 ),
    .Z(\V1/V4/V2/s1 [3]));
 OR2_X1 \V1/V4/V2/A1/M4/_0_  (.A1(\V1/V4/V2/A1/M4/c1 ),
    .A2(\V1/V4/V2/A1/M4/c2 ),
    .ZN(\V1/V4/V2/c1 ));
 AND2_X1 \V1/V4/V2/A2/M1/M1/_0_  (.A1(\V1/V4/V2/s1 [0]),
    .A2(\V1/V4/V2/v1 [2]),
    .ZN(\V1/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M1/M1/_1_  (.A(\V1/V4/V2/s1 [0]),
    .B(\V1/V4/V2/v1 [2]),
    .Z(\V1/V4/V2/A2/M1/s1 ));
 AND2_X1 \V1/V4/V2/A2/M1/M2/_0_  (.A1(\V1/V4/V2/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M1/M2/_1_  (.A(\V1/V4/V2/A2/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/v2 [2]));
 OR2_X1 \V1/V4/V2/A2/M1/_0_  (.A1(\V1/V4/V2/A2/M1/c1 ),
    .A2(\V1/V4/V2/A2/M1/c2 ),
    .ZN(\V1/V4/V2/A2/c1 ));
 AND2_X1 \V1/V4/V2/A2/M2/M1/_0_  (.A1(\V1/V4/V2/s1 [1]),
    .A2(\V1/V4/V2/v1 [3]),
    .ZN(\V1/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M2/M1/_1_  (.A(\V1/V4/V2/s1 [1]),
    .B(\V1/V4/V2/v1 [3]),
    .Z(\V1/V4/V2/A2/M2/s1 ));
 AND2_X1 \V1/V4/V2/A2/M2/M2/_0_  (.A1(\V1/V4/V2/A2/M2/s1 ),
    .A2(\V1/V4/V2/A2/c1 ),
    .ZN(\V1/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M2/M2/_1_  (.A(\V1/V4/V2/A2/M2/s1 ),
    .B(\V1/V4/V2/A2/c1 ),
    .Z(\V1/V4/v2 [3]));
 OR2_X1 \V1/V4/V2/A2/M2/_0_  (.A1(\V1/V4/V2/A2/M2/c1 ),
    .A2(\V1/V4/V2/A2/M2/c2 ),
    .ZN(\V1/V4/V2/A2/c2 ));
 AND2_X1 \V1/V4/V2/A2/M3/M1/_0_  (.A1(\V1/V4/V2/s1 [2]),
    .A2(net5),
    .ZN(\V1/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M3/M1/_1_  (.A(\V1/V4/V2/s1 [2]),
    .B(net5),
    .Z(\V1/V4/V2/A2/M3/s1 ));
 AND2_X1 \V1/V4/V2/A2/M3/M2/_0_  (.A1(\V1/V4/V2/A2/M3/s1 ),
    .A2(\V1/V4/V2/A2/c2 ),
    .ZN(\V1/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M3/M2/_1_  (.A(\V1/V4/V2/A2/M3/s1 ),
    .B(\V1/V4/V2/A2/c2 ),
    .Z(\V1/V4/V2/s2 [2]));
 OR2_X1 \V1/V4/V2/A2/M3/_0_  (.A1(\V1/V4/V2/A2/M3/c1 ),
    .A2(\V1/V4/V2/A2/M3/c2 ),
    .ZN(\V1/V4/V2/A2/c3 ));
 AND2_X1 \V1/V4/V2/A2/M4/M1/_0_  (.A1(\V1/V4/V2/s1 [3]),
    .A2(net5),
    .ZN(\V1/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A2/M4/M1/_1_  (.A(\V1/V4/V2/s1 [3]),
    .B(net5),
    .Z(\V1/V4/V2/A2/M4/s1 ));
 AND2_X1 \V1/V4/V2/A2/M4/M2/_0_  (.A1(\V1/V4/V2/A2/M4/s1 ),
    .A2(\V1/V4/V2/A2/c3 ),
    .ZN(\V1/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A2/M4/M2/_1_  (.A(\V1/V4/V2/A2/M4/s1 ),
    .B(\V1/V4/V2/A2/c3 ),
    .Z(\V1/V4/V2/s2 [3]));
 OR2_X1 \V1/V4/V2/A2/M4/_0_  (.A1(\V1/V4/V2/A2/M4/c1 ),
    .A2(\V1/V4/V2/A2/M4/c2 ),
    .ZN(\V1/V4/V2/c2 ));
 AND2_X1 \V1/V4/V2/A3/M1/M1/_0_  (.A1(\V1/V4/V2/v4 [0]),
    .A2(\V1/V4/V2/s2 [2]),
    .ZN(\V1/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M1/M1/_1_  (.A(\V1/V4/V2/v4 [0]),
    .B(\V1/V4/V2/s2 [2]),
    .Z(\V1/V4/V2/A3/M1/s1 ));
 AND2_X1 \V1/V4/V2/A3/M1/M2/_0_  (.A1(\V1/V4/V2/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M1/M2/_1_  (.A(\V1/V4/V2/A3/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/v2 [4]));
 OR2_X1 \V1/V4/V2/A3/M1/_0_  (.A1(\V1/V4/V2/A3/M1/c1 ),
    .A2(\V1/V4/V2/A3/M1/c2 ),
    .ZN(\V1/V4/V2/A3/c1 ));
 AND2_X1 \V1/V4/V2/A3/M2/M1/_0_  (.A1(\V1/V4/V2/v4 [1]),
    .A2(\V1/V4/V2/s2 [3]),
    .ZN(\V1/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M2/M1/_1_  (.A(\V1/V4/V2/v4 [1]),
    .B(\V1/V4/V2/s2 [3]),
    .Z(\V1/V4/V2/A3/M2/s1 ));
 AND2_X1 \V1/V4/V2/A3/M2/M2/_0_  (.A1(\V1/V4/V2/A3/M2/s1 ),
    .A2(\V1/V4/V2/A3/c1 ),
    .ZN(\V1/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M2/M2/_1_  (.A(\V1/V4/V2/A3/M2/s1 ),
    .B(\V1/V4/V2/A3/c1 ),
    .Z(\V1/V4/v2 [5]));
 OR2_X1 \V1/V4/V2/A3/M2/_0_  (.A1(\V1/V4/V2/A3/M2/c1 ),
    .A2(\V1/V4/V2/A3/M2/c2 ),
    .ZN(\V1/V4/V2/A3/c2 ));
 AND2_X1 \V1/V4/V2/A3/M3/M1/_0_  (.A1(\V1/V4/V2/v4 [2]),
    .A2(\V1/V4/V2/c3 ),
    .ZN(\V1/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M3/M1/_1_  (.A(\V1/V4/V2/v4 [2]),
    .B(\V1/V4/V2/c3 ),
    .Z(\V1/V4/V2/A3/M3/s1 ));
 AND2_X1 \V1/V4/V2/A3/M3/M2/_0_  (.A1(\V1/V4/V2/A3/M3/s1 ),
    .A2(\V1/V4/V2/A3/c2 ),
    .ZN(\V1/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M3/M2/_1_  (.A(\V1/V4/V2/A3/M3/s1 ),
    .B(\V1/V4/V2/A3/c2 ),
    .Z(\V1/V4/v2 [6]));
 OR2_X1 \V1/V4/V2/A3/M3/_0_  (.A1(\V1/V4/V2/A3/M3/c1 ),
    .A2(\V1/V4/V2/A3/M3/c2 ),
    .ZN(\V1/V4/V2/A3/c3 ));
 AND2_X1 \V1/V4/V2/A3/M4/M1/_0_  (.A1(\V1/V4/V2/v4 [3]),
    .A2(net5),
    .ZN(\V1/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V2/A3/M4/M1/_1_  (.A(\V1/V4/V2/v4 [3]),
    .B(net5),
    .Z(\V1/V4/V2/A3/M4/s1 ));
 AND2_X1 \V1/V4/V2/A3/M4/M2/_0_  (.A1(\V1/V4/V2/A3/M4/s1 ),
    .A2(\V1/V4/V2/A3/c3 ),
    .ZN(\V1/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V2/A3/M4/M2/_1_  (.A(\V1/V4/V2/A3/M4/s1 ),
    .B(\V1/V4/V2/A3/c3 ),
    .Z(\V1/V4/v2 [7]));
 OR2_X1 \V1/V4/V2/A3/M4/_0_  (.A1(\V1/V4/V2/A3/M4/c1 ),
    .A2(\V1/V4/V2/A3/M4/c2 ),
    .ZN(\V1/V4/V2/overflow ));
 AND2_X1 \V1/V4/V2/V1/HA1/_0_  (.A1(\V1/V4/V2/V1/w2 ),
    .A2(\V1/V4/V2/V1/w1 ),
    .ZN(\V1/V4/V2/V1/w4 ));
 XOR2_X2 \V1/V4/V2/V1/HA1/_1_  (.A(\V1/V4/V2/V1/w2 ),
    .B(\V1/V4/V2/V1/w1 ),
    .Z(\V1/V4/v2 [1]));
 AND2_X1 \V1/V4/V2/V1/HA2/_0_  (.A1(\V1/V4/V2/V1/w4 ),
    .A2(\V1/V4/V2/V1/w3 ),
    .ZN(\V1/V4/V2/v1 [3]));
 XOR2_X2 \V1/V4/V2/V1/HA2/_1_  (.A(\V1/V4/V2/V1/w4 ),
    .B(\V1/V4/V2/V1/w3 ),
    .Z(\V1/V4/V2/v1 [2]));
 AND2_X1 \V1/V4/V2/V1/_0_  (.A1(net45),
    .A2(net12),
    .ZN(\V1/V4/v2 [0]));
 AND2_X1 \V1/V4/V2/V1/_1_  (.A1(net45),
    .A2(net11),
    .ZN(\V1/V4/V2/V1/w1 ));
 AND2_X1 \V1/V4/V2/V1/_2_  (.A1(net12),
    .A2(net44),
    .ZN(\V1/V4/V2/V1/w2 ));
 AND2_X1 \V1/V4/V2/V1/_3_  (.A1(net11),
    .A2(net44),
    .ZN(\V1/V4/V2/V1/w3 ));
 AND2_X1 \V1/V4/V2/V2/HA1/_0_  (.A1(\V1/V4/V2/V2/w2 ),
    .A2(\V1/V4/V2/V2/w1 ),
    .ZN(\V1/V4/V2/V2/w4 ));
 XOR2_X2 \V1/V4/V2/V2/HA1/_1_  (.A(\V1/V4/V2/V2/w2 ),
    .B(\V1/V4/V2/V2/w1 ),
    .Z(\V1/V4/V2/v2 [1]));
 AND2_X1 \V1/V4/V2/V2/HA2/_0_  (.A1(\V1/V4/V2/V2/w4 ),
    .A2(\V1/V4/V2/V2/w3 ),
    .ZN(\V1/V4/V2/v2 [3]));
 XOR2_X2 \V1/V4/V2/V2/HA2/_1_  (.A(\V1/V4/V2/V2/w4 ),
    .B(\V1/V4/V2/V2/w3 ),
    .Z(\V1/V4/V2/v2 [2]));
 AND2_X1 \V1/V4/V2/V2/_0_  (.A1(net43),
    .A2(net12),
    .ZN(\V1/V4/V2/v2 [0]));
 AND2_X1 \V1/V4/V2/V2/_1_  (.A1(net43),
    .A2(net11),
    .ZN(\V1/V4/V2/V2/w1 ));
 AND2_X1 \V1/V4/V2/V2/_2_  (.A1(net12),
    .A2(net42),
    .ZN(\V1/V4/V2/V2/w2 ));
 AND2_X1 \V1/V4/V2/V2/_3_  (.A1(net11),
    .A2(net42),
    .ZN(\V1/V4/V2/V2/w3 ));
 AND2_X1 \V1/V4/V2/V3/HA1/_0_  (.A1(\V1/V4/V2/V3/w2 ),
    .A2(\V1/V4/V2/V3/w1 ),
    .ZN(\V1/V4/V2/V3/w4 ));
 XOR2_X2 \V1/V4/V2/V3/HA1/_1_  (.A(\V1/V4/V2/V3/w2 ),
    .B(\V1/V4/V2/V3/w1 ),
    .Z(\V1/V4/V2/v3 [1]));
 AND2_X1 \V1/V4/V2/V3/HA2/_0_  (.A1(\V1/V4/V2/V3/w4 ),
    .A2(\V1/V4/V2/V3/w3 ),
    .ZN(\V1/V4/V2/v3 [3]));
 XOR2_X2 \V1/V4/V2/V3/HA2/_1_  (.A(\V1/V4/V2/V3/w4 ),
    .B(\V1/V4/V2/V3/w3 ),
    .Z(\V1/V4/V2/v3 [2]));
 AND2_X1 \V1/V4/V2/V3/_0_  (.A1(net45),
    .A2(B[10]),
    .ZN(\V1/V4/V2/v3 [0]));
 AND2_X1 \V1/V4/V2/V3/_1_  (.A1(net45),
    .A2(B[11]),
    .ZN(\V1/V4/V2/V3/w1 ));
 AND2_X1 \V1/V4/V2/V3/_2_  (.A1(B[10]),
    .A2(net44),
    .ZN(\V1/V4/V2/V3/w2 ));
 AND2_X1 \V1/V4/V2/V3/_3_  (.A1(B[11]),
    .A2(net44),
    .ZN(\V1/V4/V2/V3/w3 ));
 AND2_X1 \V1/V4/V2/V4/HA1/_0_  (.A1(\V1/V4/V2/V4/w2 ),
    .A2(\V1/V4/V2/V4/w1 ),
    .ZN(\V1/V4/V2/V4/w4 ));
 XOR2_X2 \V1/V4/V2/V4/HA1/_1_  (.A(\V1/V4/V2/V4/w2 ),
    .B(\V1/V4/V2/V4/w1 ),
    .Z(\V1/V4/V2/v4 [1]));
 AND2_X1 \V1/V4/V2/V4/HA2/_0_  (.A1(\V1/V4/V2/V4/w4 ),
    .A2(\V1/V4/V2/V4/w3 ),
    .ZN(\V1/V4/V2/v4 [3]));
 XOR2_X2 \V1/V4/V2/V4/HA2/_1_  (.A(\V1/V4/V2/V4/w4 ),
    .B(\V1/V4/V2/V4/w3 ),
    .Z(\V1/V4/V2/v4 [2]));
 AND2_X1 \V1/V4/V2/V4/_0_  (.A1(net43),
    .A2(B[10]),
    .ZN(\V1/V4/V2/v4 [0]));
 AND2_X1 \V1/V4/V2/V4/_1_  (.A1(net43),
    .A2(B[11]),
    .ZN(\V1/V4/V2/V4/w1 ));
 AND2_X1 \V1/V4/V2/V4/_2_  (.A1(B[10]),
    .A2(net42),
    .ZN(\V1/V4/V2/V4/w2 ));
 AND2_X1 \V1/V4/V2/V4/_3_  (.A1(B[11]),
    .A2(net42),
    .ZN(\V1/V4/V2/V4/w3 ));
 OR2_X1 \V1/V4/V2/_0_  (.A1(\V1/V4/V2/c1 ),
    .A2(\V1/V4/V2/c2 ),
    .ZN(\V1/V4/V2/c3 ));
 AND2_X1 \V1/V4/V3/A1/M1/M1/_0_  (.A1(\V1/V4/V3/v2 [0]),
    .A2(\V1/V4/V3/v3 [0]),
    .ZN(\V1/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M1/M1/_1_  (.A(\V1/V4/V3/v2 [0]),
    .B(\V1/V4/V3/v3 [0]),
    .Z(\V1/V4/V3/A1/M1/s1 ));
 AND2_X1 \V1/V4/V3/A1/M1/M2/_0_  (.A1(\V1/V4/V3/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M1/M2/_1_  (.A(\V1/V4/V3/A1/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/V3/s1 [0]));
 OR2_X1 \V1/V4/V3/A1/M1/_0_  (.A1(\V1/V4/V3/A1/M1/c1 ),
    .A2(\V1/V4/V3/A1/M1/c2 ),
    .ZN(\V1/V4/V3/A1/c1 ));
 AND2_X1 \V1/V4/V3/A1/M2/M1/_0_  (.A1(\V1/V4/V3/v2 [1]),
    .A2(\V1/V4/V3/v3 [1]),
    .ZN(\V1/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M2/M1/_1_  (.A(\V1/V4/V3/v2 [1]),
    .B(\V1/V4/V3/v3 [1]),
    .Z(\V1/V4/V3/A1/M2/s1 ));
 AND2_X1 \V1/V4/V3/A1/M2/M2/_0_  (.A1(\V1/V4/V3/A1/M2/s1 ),
    .A2(\V1/V4/V3/A1/c1 ),
    .ZN(\V1/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M2/M2/_1_  (.A(\V1/V4/V3/A1/M2/s1 ),
    .B(\V1/V4/V3/A1/c1 ),
    .Z(\V1/V4/V3/s1 [1]));
 OR2_X1 \V1/V4/V3/A1/M2/_0_  (.A1(\V1/V4/V3/A1/M2/c1 ),
    .A2(\V1/V4/V3/A1/M2/c2 ),
    .ZN(\V1/V4/V3/A1/c2 ));
 AND2_X1 \V1/V4/V3/A1/M3/M1/_0_  (.A1(\V1/V4/V3/v2 [2]),
    .A2(\V1/V4/V3/v3 [2]),
    .ZN(\V1/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M3/M1/_1_  (.A(\V1/V4/V3/v2 [2]),
    .B(\V1/V4/V3/v3 [2]),
    .Z(\V1/V4/V3/A1/M3/s1 ));
 AND2_X1 \V1/V4/V3/A1/M3/M2/_0_  (.A1(\V1/V4/V3/A1/M3/s1 ),
    .A2(\V1/V4/V3/A1/c2 ),
    .ZN(\V1/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M3/M2/_1_  (.A(\V1/V4/V3/A1/M3/s1 ),
    .B(\V1/V4/V3/A1/c2 ),
    .Z(\V1/V4/V3/s1 [2]));
 OR2_X1 \V1/V4/V3/A1/M3/_0_  (.A1(\V1/V4/V3/A1/M3/c1 ),
    .A2(\V1/V4/V3/A1/M3/c2 ),
    .ZN(\V1/V4/V3/A1/c3 ));
 AND2_X1 \V1/V4/V3/A1/M4/M1/_0_  (.A1(\V1/V4/V3/v2 [3]),
    .A2(\V1/V4/V3/v3 [3]),
    .ZN(\V1/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A1/M4/M1/_1_  (.A(\V1/V4/V3/v2 [3]),
    .B(\V1/V4/V3/v3 [3]),
    .Z(\V1/V4/V3/A1/M4/s1 ));
 AND2_X1 \V1/V4/V3/A1/M4/M2/_0_  (.A1(\V1/V4/V3/A1/M4/s1 ),
    .A2(\V1/V4/V3/A1/c3 ),
    .ZN(\V1/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A1/M4/M2/_1_  (.A(\V1/V4/V3/A1/M4/s1 ),
    .B(\V1/V4/V3/A1/c3 ),
    .Z(\V1/V4/V3/s1 [3]));
 OR2_X1 \V1/V4/V3/A1/M4/_0_  (.A1(\V1/V4/V3/A1/M4/c1 ),
    .A2(\V1/V4/V3/A1/M4/c2 ),
    .ZN(\V1/V4/V3/c1 ));
 AND2_X1 \V1/V4/V3/A2/M1/M1/_0_  (.A1(\V1/V4/V3/s1 [0]),
    .A2(\V1/V4/V3/v1 [2]),
    .ZN(\V1/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M1/M1/_1_  (.A(\V1/V4/V3/s1 [0]),
    .B(\V1/V4/V3/v1 [2]),
    .Z(\V1/V4/V3/A2/M1/s1 ));
 AND2_X1 \V1/V4/V3/A2/M1/M2/_0_  (.A1(\V1/V4/V3/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M1/M2/_1_  (.A(\V1/V4/V3/A2/M1/s1 ),
    .B(net5),
    .Z(\V1/V4/v3 [2]));
 OR2_X1 \V1/V4/V3/A2/M1/_0_  (.A1(\V1/V4/V3/A2/M1/c1 ),
    .A2(\V1/V4/V3/A2/M1/c2 ),
    .ZN(\V1/V4/V3/A2/c1 ));
 AND2_X1 \V1/V4/V3/A2/M2/M1/_0_  (.A1(\V1/V4/V3/s1 [1]),
    .A2(\V1/V4/V3/v1 [3]),
    .ZN(\V1/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M2/M1/_1_  (.A(\V1/V4/V3/s1 [1]),
    .B(\V1/V4/V3/v1 [3]),
    .Z(\V1/V4/V3/A2/M2/s1 ));
 AND2_X1 \V1/V4/V3/A2/M2/M2/_0_  (.A1(\V1/V4/V3/A2/M2/s1 ),
    .A2(\V1/V4/V3/A2/c1 ),
    .ZN(\V1/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M2/M2/_1_  (.A(\V1/V4/V3/A2/M2/s1 ),
    .B(\V1/V4/V3/A2/c1 ),
    .Z(\V1/V4/v3 [3]));
 OR2_X1 \V1/V4/V3/A2/M2/_0_  (.A1(\V1/V4/V3/A2/M2/c1 ),
    .A2(\V1/V4/V3/A2/M2/c2 ),
    .ZN(\V1/V4/V3/A2/c2 ));
 AND2_X1 \V1/V4/V3/A2/M3/M1/_0_  (.A1(\V1/V4/V3/s1 [2]),
    .A2(net5),
    .ZN(\V1/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M3/M1/_1_  (.A(\V1/V4/V3/s1 [2]),
    .B(net5),
    .Z(\V1/V4/V3/A2/M3/s1 ));
 AND2_X1 \V1/V4/V3/A2/M3/M2/_0_  (.A1(\V1/V4/V3/A2/M3/s1 ),
    .A2(\V1/V4/V3/A2/c2 ),
    .ZN(\V1/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M3/M2/_1_  (.A(\V1/V4/V3/A2/M3/s1 ),
    .B(\V1/V4/V3/A2/c2 ),
    .Z(\V1/V4/V3/s2 [2]));
 OR2_X1 \V1/V4/V3/A2/M3/_0_  (.A1(\V1/V4/V3/A2/M3/c1 ),
    .A2(\V1/V4/V3/A2/M3/c2 ),
    .ZN(\V1/V4/V3/A2/c3 ));
 AND2_X1 \V1/V4/V3/A2/M4/M1/_0_  (.A1(\V1/V4/V3/s1 [3]),
    .A2(net5),
    .ZN(\V1/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A2/M4/M1/_1_  (.A(\V1/V4/V3/s1 [3]),
    .B(net5),
    .Z(\V1/V4/V3/A2/M4/s1 ));
 AND2_X1 \V1/V4/V3/A2/M4/M2/_0_  (.A1(\V1/V4/V3/A2/M4/s1 ),
    .A2(\V1/V4/V3/A2/c3 ),
    .ZN(\V1/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A2/M4/M2/_1_  (.A(\V1/V4/V3/A2/M4/s1 ),
    .B(\V1/V4/V3/A2/c3 ),
    .Z(\V1/V4/V3/s2 [3]));
 OR2_X1 \V1/V4/V3/A2/M4/_0_  (.A1(\V1/V4/V3/A2/M4/c1 ),
    .A2(\V1/V4/V3/A2/M4/c2 ),
    .ZN(\V1/V4/V3/c2 ));
 AND2_X1 \V1/V4/V3/A3/M1/M1/_0_  (.A1(\V1/V4/V3/v4 [0]),
    .A2(\V1/V4/V3/s2 [2]),
    .ZN(\V1/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M1/M1/_1_  (.A(\V1/V4/V3/v4 [0]),
    .B(\V1/V4/V3/s2 [2]),
    .Z(\V1/V4/V3/A3/M1/s1 ));
 AND2_X1 \V1/V4/V3/A3/M1/M2/_0_  (.A1(\V1/V4/V3/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V1/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M1/M2/_1_  (.A(\V1/V4/V3/A3/M1/s1 ),
    .B(net4),
    .Z(\V1/V4/v3 [4]));
 OR2_X1 \V1/V4/V3/A3/M1/_0_  (.A1(\V1/V4/V3/A3/M1/c1 ),
    .A2(\V1/V4/V3/A3/M1/c2 ),
    .ZN(\V1/V4/V3/A3/c1 ));
 AND2_X1 \V1/V4/V3/A3/M2/M1/_0_  (.A1(\V1/V4/V3/v4 [1]),
    .A2(\V1/V4/V3/s2 [3]),
    .ZN(\V1/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M2/M1/_1_  (.A(\V1/V4/V3/v4 [1]),
    .B(\V1/V4/V3/s2 [3]),
    .Z(\V1/V4/V3/A3/M2/s1 ));
 AND2_X1 \V1/V4/V3/A3/M2/M2/_0_  (.A1(\V1/V4/V3/A3/M2/s1 ),
    .A2(\V1/V4/V3/A3/c1 ),
    .ZN(\V1/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M2/M2/_1_  (.A(\V1/V4/V3/A3/M2/s1 ),
    .B(\V1/V4/V3/A3/c1 ),
    .Z(\V1/V4/v3 [5]));
 OR2_X1 \V1/V4/V3/A3/M2/_0_  (.A1(\V1/V4/V3/A3/M2/c1 ),
    .A2(\V1/V4/V3/A3/M2/c2 ),
    .ZN(\V1/V4/V3/A3/c2 ));
 AND2_X1 \V1/V4/V3/A3/M3/M1/_0_  (.A1(\V1/V4/V3/v4 [2]),
    .A2(\V1/V4/V3/c3 ),
    .ZN(\V1/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M3/M1/_1_  (.A(\V1/V4/V3/v4 [2]),
    .B(\V1/V4/V3/c3 ),
    .Z(\V1/V4/V3/A3/M3/s1 ));
 AND2_X1 \V1/V4/V3/A3/M3/M2/_0_  (.A1(\V1/V4/V3/A3/M3/s1 ),
    .A2(\V1/V4/V3/A3/c2 ),
    .ZN(\V1/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M3/M2/_1_  (.A(\V1/V4/V3/A3/M3/s1 ),
    .B(\V1/V4/V3/A3/c2 ),
    .Z(\V1/V4/v3 [6]));
 OR2_X1 \V1/V4/V3/A3/M3/_0_  (.A1(\V1/V4/V3/A3/M3/c1 ),
    .A2(\V1/V4/V3/A3/M3/c2 ),
    .ZN(\V1/V4/V3/A3/c3 ));
 AND2_X1 \V1/V4/V3/A3/M4/M1/_0_  (.A1(\V1/V4/V3/v4 [3]),
    .A2(net5),
    .ZN(\V1/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V3/A3/M4/M1/_1_  (.A(\V1/V4/V3/v4 [3]),
    .B(net5),
    .Z(\V1/V4/V3/A3/M4/s1 ));
 AND2_X1 \V1/V4/V3/A3/M4/M2/_0_  (.A1(\V1/V4/V3/A3/M4/s1 ),
    .A2(\V1/V4/V3/A3/c3 ),
    .ZN(\V1/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V3/A3/M4/M2/_1_  (.A(\V1/V4/V3/A3/M4/s1 ),
    .B(\V1/V4/V3/A3/c3 ),
    .Z(\V1/V4/v3 [7]));
 OR2_X1 \V1/V4/V3/A3/M4/_0_  (.A1(\V1/V4/V3/A3/M4/c1 ),
    .A2(\V1/V4/V3/A3/M4/c2 ),
    .ZN(\V1/V4/V3/overflow ));
 AND2_X1 \V1/V4/V3/V1/HA1/_0_  (.A1(\V1/V4/V3/V1/w2 ),
    .A2(\V1/V4/V3/V1/w1 ),
    .ZN(\V1/V4/V3/V1/w4 ));
 XOR2_X2 \V1/V4/V3/V1/HA1/_1_  (.A(\V1/V4/V3/V1/w2 ),
    .B(\V1/V4/V3/V1/w1 ),
    .Z(\V1/V4/v3 [1]));
 AND2_X1 \V1/V4/V3/V1/HA2/_0_  (.A1(\V1/V4/V3/V1/w4 ),
    .A2(\V1/V4/V3/V1/w3 ),
    .ZN(\V1/V4/V3/v1 [3]));
 XOR2_X2 \V1/V4/V3/V1/HA2/_1_  (.A(\V1/V4/V3/V1/w4 ),
    .B(\V1/V4/V3/V1/w3 ),
    .Z(\V1/V4/V3/v1 [2]));
 AND2_X1 \V1/V4/V3/V1/_0_  (.A1(net25),
    .A2(B[12]),
    .ZN(\V1/V4/v3 [0]));
 AND2_X1 \V1/V4/V3/V1/_1_  (.A1(net25),
    .A2(B[13]),
    .ZN(\V1/V4/V3/V1/w1 ));
 AND2_X1 \V1/V4/V3/V1/_2_  (.A1(B[12]),
    .A2(net24),
    .ZN(\V1/V4/V3/V1/w2 ));
 AND2_X1 \V1/V4/V3/V1/_3_  (.A1(B[13]),
    .A2(net24),
    .ZN(\V1/V4/V3/V1/w3 ));
 AND2_X1 \V1/V4/V3/V2/HA1/_0_  (.A1(\V1/V4/V3/V2/w2 ),
    .A2(\V1/V4/V3/V2/w1 ),
    .ZN(\V1/V4/V3/V2/w4 ));
 XOR2_X2 \V1/V4/V3/V2/HA1/_1_  (.A(\V1/V4/V3/V2/w2 ),
    .B(\V1/V4/V3/V2/w1 ),
    .Z(\V1/V4/V3/v2 [1]));
 AND2_X1 \V1/V4/V3/V2/HA2/_0_  (.A1(\V1/V4/V3/V2/w4 ),
    .A2(\V1/V4/V3/V2/w3 ),
    .ZN(\V1/V4/V3/v2 [3]));
 XOR2_X2 \V1/V4/V3/V2/HA2/_1_  (.A(\V1/V4/V3/V2/w4 ),
    .B(\V1/V4/V3/V2/w3 ),
    .Z(\V1/V4/V3/v2 [2]));
 AND2_X1 \V1/V4/V3/V2/_0_  (.A1(net47),
    .A2(B[12]),
    .ZN(\V1/V4/V3/v2 [0]));
 AND2_X1 \V1/V4/V3/V2/_1_  (.A1(net47),
    .A2(B[13]),
    .ZN(\V1/V4/V3/V2/w1 ));
 AND2_X1 \V1/V4/V3/V2/_2_  (.A1(B[12]),
    .A2(net46),
    .ZN(\V1/V4/V3/V2/w2 ));
 AND2_X1 \V1/V4/V3/V2/_3_  (.A1(B[13]),
    .A2(net46),
    .ZN(\V1/V4/V3/V2/w3 ));
 AND2_X1 \V1/V4/V3/V3/HA1/_0_  (.A1(\V1/V4/V3/V3/w2 ),
    .A2(\V1/V4/V3/V3/w1 ),
    .ZN(\V1/V4/V3/V3/w4 ));
 XOR2_X2 \V1/V4/V3/V3/HA1/_1_  (.A(\V1/V4/V3/V3/w2 ),
    .B(\V1/V4/V3/V3/w1 ),
    .Z(\V1/V4/V3/v3 [1]));
 AND2_X1 \V1/V4/V3/V3/HA2/_0_  (.A1(\V1/V4/V3/V3/w4 ),
    .A2(\V1/V4/V3/V3/w3 ),
    .ZN(\V1/V4/V3/v3 [3]));
 XOR2_X2 \V1/V4/V3/V3/HA2/_1_  (.A(\V1/V4/V3/V3/w4 ),
    .B(\V1/V4/V3/V3/w3 ),
    .Z(\V1/V4/V3/v3 [2]));
 AND2_X1 \V1/V4/V3/V3/_0_  (.A1(net25),
    .A2(B[14]),
    .ZN(\V1/V4/V3/v3 [0]));
 AND2_X1 \V1/V4/V3/V3/_1_  (.A1(net25),
    .A2(B[15]),
    .ZN(\V1/V4/V3/V3/w1 ));
 AND2_X1 \V1/V4/V3/V3/_2_  (.A1(B[14]),
    .A2(net24),
    .ZN(\V1/V4/V3/V3/w2 ));
 AND2_X1 \V1/V4/V3/V3/_3_  (.A1(B[15]),
    .A2(net24),
    .ZN(\V1/V4/V3/V3/w3 ));
 AND2_X1 \V1/V4/V3/V4/HA1/_0_  (.A1(\V1/V4/V3/V4/w2 ),
    .A2(\V1/V4/V3/V4/w1 ),
    .ZN(\V1/V4/V3/V4/w4 ));
 XOR2_X2 \V1/V4/V3/V4/HA1/_1_  (.A(\V1/V4/V3/V4/w2 ),
    .B(\V1/V4/V3/V4/w1 ),
    .Z(\V1/V4/V3/v4 [1]));
 AND2_X1 \V1/V4/V3/V4/HA2/_0_  (.A1(\V1/V4/V3/V4/w4 ),
    .A2(\V1/V4/V3/V4/w3 ),
    .ZN(\V1/V4/V3/v4 [3]));
 XOR2_X2 \V1/V4/V3/V4/HA2/_1_  (.A(\V1/V4/V3/V4/w4 ),
    .B(\V1/V4/V3/V4/w3 ),
    .Z(\V1/V4/V3/v4 [2]));
 AND2_X1 \V1/V4/V3/V4/_0_  (.A1(net47),
    .A2(B[14]),
    .ZN(\V1/V4/V3/v4 [0]));
 AND2_X1 \V1/V4/V3/V4/_1_  (.A1(net47),
    .A2(B[15]),
    .ZN(\V1/V4/V3/V4/w1 ));
 AND2_X1 \V1/V4/V3/V4/_2_  (.A1(B[14]),
    .A2(net46),
    .ZN(\V1/V4/V3/V4/w2 ));
 AND2_X1 \V1/V4/V3/V4/_3_  (.A1(B[15]),
    .A2(net46),
    .ZN(\V1/V4/V3/V4/w3 ));
 OR2_X1 \V1/V4/V3/_0_  (.A1(\V1/V4/V3/c1 ),
    .A2(\V1/V4/V3/c2 ),
    .ZN(\V1/V4/V3/c3 ));
 AND2_X1 \V1/V4/V4/A1/M1/M1/_0_  (.A1(\V1/V4/V4/v2 [0]),
    .A2(\V1/V4/V4/v3 [0]),
    .ZN(\V1/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M1/M1/_1_  (.A(\V1/V4/V4/v2 [0]),
    .B(\V1/V4/V4/v3 [0]),
    .Z(\V1/V4/V4/A1/M1/s1 ));
 AND2_X1 \V1/V4/V4/A1/M1/M2/_0_  (.A1(\V1/V4/V4/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M1/M2/_1_  (.A(\V1/V4/V4/A1/M1/s1 ),
    .B(net4),
    .Z(\V1/V4/V4/s1 [0]));
 OR2_X1 \V1/V4/V4/A1/M1/_0_  (.A1(\V1/V4/V4/A1/M1/c1 ),
    .A2(\V1/V4/V4/A1/M1/c2 ),
    .ZN(\V1/V4/V4/A1/c1 ));
 AND2_X1 \V1/V4/V4/A1/M2/M1/_0_  (.A1(\V1/V4/V4/v2 [1]),
    .A2(\V1/V4/V4/v3 [1]),
    .ZN(\V1/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M2/M1/_1_  (.A(\V1/V4/V4/v2 [1]),
    .B(\V1/V4/V4/v3 [1]),
    .Z(\V1/V4/V4/A1/M2/s1 ));
 AND2_X1 \V1/V4/V4/A1/M2/M2/_0_  (.A1(\V1/V4/V4/A1/M2/s1 ),
    .A2(\V1/V4/V4/A1/c1 ),
    .ZN(\V1/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M2/M2/_1_  (.A(\V1/V4/V4/A1/M2/s1 ),
    .B(\V1/V4/V4/A1/c1 ),
    .Z(\V1/V4/V4/s1 [1]));
 OR2_X1 \V1/V4/V4/A1/M2/_0_  (.A1(\V1/V4/V4/A1/M2/c1 ),
    .A2(\V1/V4/V4/A1/M2/c2 ),
    .ZN(\V1/V4/V4/A1/c2 ));
 AND2_X1 \V1/V4/V4/A1/M3/M1/_0_  (.A1(\V1/V4/V4/v2 [2]),
    .A2(\V1/V4/V4/v3 [2]),
    .ZN(\V1/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M3/M1/_1_  (.A(\V1/V4/V4/v2 [2]),
    .B(\V1/V4/V4/v3 [2]),
    .Z(\V1/V4/V4/A1/M3/s1 ));
 AND2_X1 \V1/V4/V4/A1/M3/M2/_0_  (.A1(\V1/V4/V4/A1/M3/s1 ),
    .A2(\V1/V4/V4/A1/c2 ),
    .ZN(\V1/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M3/M2/_1_  (.A(\V1/V4/V4/A1/M3/s1 ),
    .B(\V1/V4/V4/A1/c2 ),
    .Z(\V1/V4/V4/s1 [2]));
 OR2_X1 \V1/V4/V4/A1/M3/_0_  (.A1(\V1/V4/V4/A1/M3/c1 ),
    .A2(\V1/V4/V4/A1/M3/c2 ),
    .ZN(\V1/V4/V4/A1/c3 ));
 AND2_X1 \V1/V4/V4/A1/M4/M1/_0_  (.A1(\V1/V4/V4/v2 [3]),
    .A2(\V1/V4/V4/v3 [3]),
    .ZN(\V1/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A1/M4/M1/_1_  (.A(\V1/V4/V4/v2 [3]),
    .B(\V1/V4/V4/v3 [3]),
    .Z(\V1/V4/V4/A1/M4/s1 ));
 AND2_X1 \V1/V4/V4/A1/M4/M2/_0_  (.A1(\V1/V4/V4/A1/M4/s1 ),
    .A2(\V1/V4/V4/A1/c3 ),
    .ZN(\V1/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A1/M4/M2/_1_  (.A(\V1/V4/V4/A1/M4/s1 ),
    .B(\V1/V4/V4/A1/c3 ),
    .Z(\V1/V4/V4/s1 [3]));
 OR2_X1 \V1/V4/V4/A1/M4/_0_  (.A1(\V1/V4/V4/A1/M4/c1 ),
    .A2(\V1/V4/V4/A1/M4/c2 ),
    .ZN(\V1/V4/V4/c1 ));
 AND2_X1 \V1/V4/V4/A2/M1/M1/_0_  (.A1(\V1/V4/V4/s1 [0]),
    .A2(\V1/V4/V4/v1 [2]),
    .ZN(\V1/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M1/M1/_1_  (.A(\V1/V4/V4/s1 [0]),
    .B(\V1/V4/V4/v1 [2]),
    .Z(\V1/V4/V4/A2/M1/s1 ));
 AND2_X1 \V1/V4/V4/A2/M1/M2/_0_  (.A1(\V1/V4/V4/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V1/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M1/M2/_1_  (.A(\V1/V4/V4/A2/M1/s1 ),
    .B(net4),
    .Z(\V1/V4/v4 [2]));
 OR2_X1 \V1/V4/V4/A2/M1/_0_  (.A1(\V1/V4/V4/A2/M1/c1 ),
    .A2(\V1/V4/V4/A2/M1/c2 ),
    .ZN(\V1/V4/V4/A2/c1 ));
 AND2_X1 \V1/V4/V4/A2/M2/M1/_0_  (.A1(\V1/V4/V4/s1 [1]),
    .A2(\V1/V4/V4/v1 [3]),
    .ZN(\V1/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M2/M1/_1_  (.A(\V1/V4/V4/s1 [1]),
    .B(\V1/V4/V4/v1 [3]),
    .Z(\V1/V4/V4/A2/M2/s1 ));
 AND2_X1 \V1/V4/V4/A2/M2/M2/_0_  (.A1(\V1/V4/V4/A2/M2/s1 ),
    .A2(\V1/V4/V4/A2/c1 ),
    .ZN(\V1/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M2/M2/_1_  (.A(\V1/V4/V4/A2/M2/s1 ),
    .B(\V1/V4/V4/A2/c1 ),
    .Z(\V1/V4/v4 [3]));
 OR2_X1 \V1/V4/V4/A2/M2/_0_  (.A1(\V1/V4/V4/A2/M2/c1 ),
    .A2(\V1/V4/V4/A2/M2/c2 ),
    .ZN(\V1/V4/V4/A2/c2 ));
 AND2_X1 \V1/V4/V4/A2/M3/M1/_0_  (.A1(\V1/V4/V4/s1 [2]),
    .A2(net4),
    .ZN(\V1/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M3/M1/_1_  (.A(\V1/V4/V4/s1 [2]),
    .B(net4),
    .Z(\V1/V4/V4/A2/M3/s1 ));
 AND2_X1 \V1/V4/V4/A2/M3/M2/_0_  (.A1(\V1/V4/V4/A2/M3/s1 ),
    .A2(\V1/V4/V4/A2/c2 ),
    .ZN(\V1/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M3/M2/_1_  (.A(\V1/V4/V4/A2/M3/s1 ),
    .B(\V1/V4/V4/A2/c2 ),
    .Z(\V1/V4/V4/s2 [2]));
 OR2_X1 \V1/V4/V4/A2/M3/_0_  (.A1(\V1/V4/V4/A2/M3/c1 ),
    .A2(\V1/V4/V4/A2/M3/c2 ),
    .ZN(\V1/V4/V4/A2/c3 ));
 AND2_X1 \V1/V4/V4/A2/M4/M1/_0_  (.A1(\V1/V4/V4/s1 [3]),
    .A2(net4),
    .ZN(\V1/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A2/M4/M1/_1_  (.A(\V1/V4/V4/s1 [3]),
    .B(net4),
    .Z(\V1/V4/V4/A2/M4/s1 ));
 AND2_X1 \V1/V4/V4/A2/M4/M2/_0_  (.A1(\V1/V4/V4/A2/M4/s1 ),
    .A2(\V1/V4/V4/A2/c3 ),
    .ZN(\V1/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A2/M4/M2/_1_  (.A(\V1/V4/V4/A2/M4/s1 ),
    .B(\V1/V4/V4/A2/c3 ),
    .Z(\V1/V4/V4/s2 [3]));
 OR2_X1 \V1/V4/V4/A2/M4/_0_  (.A1(\V1/V4/V4/A2/M4/c1 ),
    .A2(\V1/V4/V4/A2/M4/c2 ),
    .ZN(\V1/V4/V4/c2 ));
 AND2_X1 \V1/V4/V4/A3/M1/M1/_0_  (.A1(\V1/V4/V4/v4 [0]),
    .A2(\V1/V4/V4/s2 [2]),
    .ZN(\V1/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M1/M1/_1_  (.A(\V1/V4/V4/v4 [0]),
    .B(\V1/V4/V4/s2 [2]),
    .Z(\V1/V4/V4/A3/M1/s1 ));
 AND2_X1 \V1/V4/V4/A3/M1/M2/_0_  (.A1(\V1/V4/V4/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V1/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M1/M2/_1_  (.A(\V1/V4/V4/A3/M1/s1 ),
    .B(net6),
    .Z(\V1/V4/v4 [4]));
 OR2_X1 \V1/V4/V4/A3/M1/_0_  (.A1(\V1/V4/V4/A3/M1/c1 ),
    .A2(\V1/V4/V4/A3/M1/c2 ),
    .ZN(\V1/V4/V4/A3/c1 ));
 AND2_X1 \V1/V4/V4/A3/M2/M1/_0_  (.A1(\V1/V4/V4/v4 [1]),
    .A2(\V1/V4/V4/s2 [3]),
    .ZN(\V1/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M2/M1/_1_  (.A(\V1/V4/V4/v4 [1]),
    .B(\V1/V4/V4/s2 [3]),
    .Z(\V1/V4/V4/A3/M2/s1 ));
 AND2_X1 \V1/V4/V4/A3/M2/M2/_0_  (.A1(\V1/V4/V4/A3/M2/s1 ),
    .A2(\V1/V4/V4/A3/c1 ),
    .ZN(\V1/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M2/M2/_1_  (.A(\V1/V4/V4/A3/M2/s1 ),
    .B(\V1/V4/V4/A3/c1 ),
    .Z(\V1/V4/v4 [5]));
 OR2_X1 \V1/V4/V4/A3/M2/_0_  (.A1(\V1/V4/V4/A3/M2/c1 ),
    .A2(\V1/V4/V4/A3/M2/c2 ),
    .ZN(\V1/V4/V4/A3/c2 ));
 AND2_X1 \V1/V4/V4/A3/M3/M1/_0_  (.A1(\V1/V4/V4/v4 [2]),
    .A2(\V1/V4/V4/c3 ),
    .ZN(\V1/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M3/M1/_1_  (.A(\V1/V4/V4/v4 [2]),
    .B(\V1/V4/V4/c3 ),
    .Z(\V1/V4/V4/A3/M3/s1 ));
 AND2_X1 \V1/V4/V4/A3/M3/M2/_0_  (.A1(\V1/V4/V4/A3/M3/s1 ),
    .A2(\V1/V4/V4/A3/c2 ),
    .ZN(\V1/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M3/M2/_1_  (.A(\V1/V4/V4/A3/M3/s1 ),
    .B(\V1/V4/V4/A3/c2 ),
    .Z(\V1/V4/v4 [6]));
 OR2_X1 \V1/V4/V4/A3/M3/_0_  (.A1(\V1/V4/V4/A3/M3/c1 ),
    .A2(\V1/V4/V4/A3/M3/c2 ),
    .ZN(\V1/V4/V4/A3/c3 ));
 AND2_X1 \V1/V4/V4/A3/M4/M1/_0_  (.A1(\V1/V4/V4/v4 [3]),
    .A2(net6),
    .ZN(\V1/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V1/V4/V4/A3/M4/M1/_1_  (.A(\V1/V4/V4/v4 [3]),
    .B(net6),
    .Z(\V1/V4/V4/A3/M4/s1 ));
 AND2_X1 \V1/V4/V4/A3/M4/M2/_0_  (.A1(\V1/V4/V4/A3/M4/s1 ),
    .A2(\V1/V4/V4/A3/c3 ),
    .ZN(\V1/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V1/V4/V4/A3/M4/M2/_1_  (.A(\V1/V4/V4/A3/M4/s1 ),
    .B(\V1/V4/V4/A3/c3 ),
    .Z(\V1/V4/v4 [7]));
 OR2_X1 \V1/V4/V4/A3/M4/_0_  (.A1(\V1/V4/V4/A3/M4/c1 ),
    .A2(\V1/V4/V4/A3/M4/c2 ),
    .ZN(\V1/V4/V4/overflow ));
 AND2_X1 \V1/V4/V4/V1/HA1/_0_  (.A1(\V1/V4/V4/V1/w2 ),
    .A2(\V1/V4/V4/V1/w1 ),
    .ZN(\V1/V4/V4/V1/w4 ));
 XOR2_X2 \V1/V4/V4/V1/HA1/_1_  (.A(\V1/V4/V4/V1/w2 ),
    .B(\V1/V4/V4/V1/w1 ),
    .Z(\V1/V4/v4 [1]));
 AND2_X1 \V1/V4/V4/V1/HA2/_0_  (.A1(\V1/V4/V4/V1/w4 ),
    .A2(\V1/V4/V4/V1/w3 ),
    .ZN(\V1/V4/V4/v1 [3]));
 XOR2_X2 \V1/V4/V4/V1/HA2/_1_  (.A(\V1/V4/V4/V1/w4 ),
    .B(\V1/V4/V4/V1/w3 ),
    .Z(\V1/V4/V4/v1 [2]));
 AND2_X1 \V1/V4/V4/V1/_0_  (.A1(net45),
    .A2(B[12]),
    .ZN(\V1/V4/v4 [0]));
 AND2_X1 \V1/V4/V4/V1/_1_  (.A1(net45),
    .A2(B[13]),
    .ZN(\V1/V4/V4/V1/w1 ));
 AND2_X1 \V1/V4/V4/V1/_2_  (.A1(B[12]),
    .A2(net44),
    .ZN(\V1/V4/V4/V1/w2 ));
 AND2_X1 \V1/V4/V4/V1/_3_  (.A1(B[13]),
    .A2(net44),
    .ZN(\V1/V4/V4/V1/w3 ));
 AND2_X1 \V1/V4/V4/V2/HA1/_0_  (.A1(\V1/V4/V4/V2/w2 ),
    .A2(\V1/V4/V4/V2/w1 ),
    .ZN(\V1/V4/V4/V2/w4 ));
 XOR2_X2 \V1/V4/V4/V2/HA1/_1_  (.A(\V1/V4/V4/V2/w2 ),
    .B(\V1/V4/V4/V2/w1 ),
    .Z(\V1/V4/V4/v2 [1]));
 AND2_X1 \V1/V4/V4/V2/HA2/_0_  (.A1(\V1/V4/V4/V2/w4 ),
    .A2(\V1/V4/V4/V2/w3 ),
    .ZN(\V1/V4/V4/v2 [3]));
 XOR2_X2 \V1/V4/V4/V2/HA2/_1_  (.A(\V1/V4/V4/V2/w4 ),
    .B(\V1/V4/V4/V2/w3 ),
    .Z(\V1/V4/V4/v2 [2]));
 AND2_X1 \V1/V4/V4/V2/_0_  (.A1(net43),
    .A2(B[12]),
    .ZN(\V1/V4/V4/v2 [0]));
 AND2_X1 \V1/V4/V4/V2/_1_  (.A1(net43),
    .A2(B[13]),
    .ZN(\V1/V4/V4/V2/w1 ));
 AND2_X1 \V1/V4/V4/V2/_2_  (.A1(B[12]),
    .A2(net42),
    .ZN(\V1/V4/V4/V2/w2 ));
 AND2_X1 \V1/V4/V4/V2/_3_  (.A1(B[13]),
    .A2(net42),
    .ZN(\V1/V4/V4/V2/w3 ));
 AND2_X1 \V1/V4/V4/V3/HA1/_0_  (.A1(\V1/V4/V4/V3/w2 ),
    .A2(\V1/V4/V4/V3/w1 ),
    .ZN(\V1/V4/V4/V3/w4 ));
 XOR2_X2 \V1/V4/V4/V3/HA1/_1_  (.A(\V1/V4/V4/V3/w2 ),
    .B(\V1/V4/V4/V3/w1 ),
    .Z(\V1/V4/V4/v3 [1]));
 AND2_X1 \V1/V4/V4/V3/HA2/_0_  (.A1(\V1/V4/V4/V3/w4 ),
    .A2(\V1/V4/V4/V3/w3 ),
    .ZN(\V1/V4/V4/v3 [3]));
 XOR2_X2 \V1/V4/V4/V3/HA2/_1_  (.A(\V1/V4/V4/V3/w4 ),
    .B(\V1/V4/V4/V3/w3 ),
    .Z(\V1/V4/V4/v3 [2]));
 AND2_X1 \V1/V4/V4/V3/_0_  (.A1(net45),
    .A2(B[14]),
    .ZN(\V1/V4/V4/v3 [0]));
 AND2_X1 \V1/V4/V4/V3/_1_  (.A1(net45),
    .A2(B[15]),
    .ZN(\V1/V4/V4/V3/w1 ));
 AND2_X1 \V1/V4/V4/V3/_2_  (.A1(B[14]),
    .A2(net44),
    .ZN(\V1/V4/V4/V3/w2 ));
 AND2_X1 \V1/V4/V4/V3/_3_  (.A1(B[15]),
    .A2(net44),
    .ZN(\V1/V4/V4/V3/w3 ));
 AND2_X1 \V1/V4/V4/V4/HA1/_0_  (.A1(\V1/V4/V4/V4/w2 ),
    .A2(\V1/V4/V4/V4/w1 ),
    .ZN(\V1/V4/V4/V4/w4 ));
 XOR2_X2 \V1/V4/V4/V4/HA1/_1_  (.A(\V1/V4/V4/V4/w2 ),
    .B(\V1/V4/V4/V4/w1 ),
    .Z(\V1/V4/V4/v4 [1]));
 AND2_X1 \V1/V4/V4/V4/HA2/_0_  (.A1(\V1/V4/V4/V4/w4 ),
    .A2(\V1/V4/V4/V4/w3 ),
    .ZN(\V1/V4/V4/v4 [3]));
 XOR2_X2 \V1/V4/V4/V4/HA2/_1_  (.A(\V1/V4/V4/V4/w4 ),
    .B(\V1/V4/V4/V4/w3 ),
    .Z(\V1/V4/V4/v4 [2]));
 AND2_X1 \V1/V4/V4/V4/_0_  (.A1(net43),
    .A2(B[14]),
    .ZN(\V1/V4/V4/v4 [0]));
 AND2_X1 \V1/V4/V4/V4/_1_  (.A1(net43),
    .A2(B[15]),
    .ZN(\V1/V4/V4/V4/w1 ));
 AND2_X1 \V1/V4/V4/V4/_2_  (.A1(B[14]),
    .A2(net42),
    .ZN(\V1/V4/V4/V4/w2 ));
 AND2_X1 \V1/V4/V4/V4/_3_  (.A1(B[15]),
    .A2(net42),
    .ZN(\V1/V4/V4/V4/w3 ));
 OR2_X1 \V1/V4/V4/_0_  (.A1(\V1/V4/V4/c1 ),
    .A2(\V1/V4/V4/c2 ),
    .ZN(\V1/V4/V4/c3 ));
 OR2_X1 \V1/V4/_0_  (.A1(\V1/V4/c1 ),
    .A2(\V1/V4/c2 ),
    .ZN(\V1/V4/c3 ));
 OR2_X2 \V1/_0_  (.A1(\V1/c1 ),
    .A2(\V1/c2 ),
    .ZN(\V1/c3 ));
 AND2_X1 \V2/A1/A1/A1/M1/M1/_0_  (.A1(\V2/v2 [0]),
    .A2(\V2/v3 [0]),
    .ZN(\V2/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M1/M1/_1_  (.A(\V2/v2 [0]),
    .B(\V2/v3 [0]),
    .Z(\V2/A1/A1/A1/M1/s1 ));
 AND2_X1 \V2/A1/A1/A1/M1/M2/_0_  (.A1(\V2/A1/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V2/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M1/M2/_1_  (.A(\V2/A1/A1/A1/M1/s1 ),
    .B(net6),
    .Z(\V2/s1 [0]));
 OR2_X1 \V2/A1/A1/A1/M1/_0_  (.A1(\V2/A1/A1/A1/M1/c1 ),
    .A2(\V2/A1/A1/A1/M1/c2 ),
    .ZN(\V2/A1/A1/A1/c1 ));
 AND2_X1 \V2/A1/A1/A1/M2/M1/_0_  (.A1(\V2/v2 [1]),
    .A2(\V2/v3 [1]),
    .ZN(\V2/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M2/M1/_1_  (.A(\V2/v2 [1]),
    .B(\V2/v3 [1]),
    .Z(\V2/A1/A1/A1/M2/s1 ));
 AND2_X1 \V2/A1/A1/A1/M2/M2/_0_  (.A1(\V2/A1/A1/A1/M2/s1 ),
    .A2(\V2/A1/A1/A1/c1 ),
    .ZN(\V2/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M2/M2/_1_  (.A(\V2/A1/A1/A1/M2/s1 ),
    .B(\V2/A1/A1/A1/c1 ),
    .Z(\V2/s1 [1]));
 OR2_X1 \V2/A1/A1/A1/M2/_0_  (.A1(\V2/A1/A1/A1/M2/c1 ),
    .A2(\V2/A1/A1/A1/M2/c2 ),
    .ZN(\V2/A1/A1/A1/c2 ));
 AND2_X1 \V2/A1/A1/A1/M3/M1/_0_  (.A1(\V2/v2 [2]),
    .A2(\V2/v3 [2]),
    .ZN(\V2/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M3/M1/_1_  (.A(\V2/v2 [2]),
    .B(\V2/v3 [2]),
    .Z(\V2/A1/A1/A1/M3/s1 ));
 AND2_X1 \V2/A1/A1/A1/M3/M2/_0_  (.A1(\V2/A1/A1/A1/M3/s1 ),
    .A2(\V2/A1/A1/A1/c2 ),
    .ZN(\V2/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M3/M2/_1_  (.A(\V2/A1/A1/A1/M3/s1 ),
    .B(\V2/A1/A1/A1/c2 ),
    .Z(\V2/s1 [2]));
 OR2_X1 \V2/A1/A1/A1/M3/_0_  (.A1(\V2/A1/A1/A1/M3/c1 ),
    .A2(\V2/A1/A1/A1/M3/c2 ),
    .ZN(\V2/A1/A1/A1/c3 ));
 AND2_X1 \V2/A1/A1/A1/M4/M1/_0_  (.A1(\V2/v2 [3]),
    .A2(\V2/v3 [3]),
    .ZN(\V2/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A1/A1/A1/M4/M1/_1_  (.A(\V2/v2 [3]),
    .B(\V2/v3 [3]),
    .Z(\V2/A1/A1/A1/M4/s1 ));
 AND2_X1 \V2/A1/A1/A1/M4/M2/_0_  (.A1(\V2/A1/A1/A1/M4/s1 ),
    .A2(\V2/A1/A1/A1/c3 ),
    .ZN(\V2/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A1/A1/A1/M4/M2/_1_  (.A(\V2/A1/A1/A1/M4/s1 ),
    .B(\V2/A1/A1/A1/c3 ),
    .Z(\V2/s1 [3]));
 OR2_X1 \V2/A1/A1/A1/M4/_0_  (.A1(\V2/A1/A1/A1/M4/c1 ),
    .A2(\V2/A1/A1/A1/M4/c2 ),
    .ZN(\V2/A1/A1/c1 ));
 AND2_X1 \V2/A1/A1/A2/M1/M1/_0_  (.A1(\V2/v2 [4]),
    .A2(\V2/v3 [4]),
    .ZN(\V2/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M1/M1/_1_  (.A(\V2/v2 [4]),
    .B(\V2/v3 [4]),
    .Z(\V2/A1/A1/A2/M1/s1 ));
 AND2_X1 \V2/A1/A1/A2/M1/M2/_0_  (.A1(\V2/A1/A1/A2/M1/s1 ),
    .A2(\V2/A1/A1/c1 ),
    .ZN(\V2/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M1/M2/_1_  (.A(\V2/A1/A1/A2/M1/s1 ),
    .B(\V2/A1/A1/c1 ),
    .Z(\V2/s1 [4]));
 OR2_X1 \V2/A1/A1/A2/M1/_0_  (.A1(\V2/A1/A1/A2/M1/c1 ),
    .A2(\V2/A1/A1/A2/M1/c2 ),
    .ZN(\V2/A1/A1/A2/c1 ));
 AND2_X1 \V2/A1/A1/A2/M2/M1/_0_  (.A1(\V2/v2 [5]),
    .A2(\V2/v3 [5]),
    .ZN(\V2/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M2/M1/_1_  (.A(\V2/v2 [5]),
    .B(\V2/v3 [5]),
    .Z(\V2/A1/A1/A2/M2/s1 ));
 AND2_X1 \V2/A1/A1/A2/M2/M2/_0_  (.A1(\V2/A1/A1/A2/M2/s1 ),
    .A2(\V2/A1/A1/A2/c1 ),
    .ZN(\V2/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M2/M2/_1_  (.A(\V2/A1/A1/A2/M2/s1 ),
    .B(\V2/A1/A1/A2/c1 ),
    .Z(\V2/s1 [5]));
 OR2_X1 \V2/A1/A1/A2/M2/_0_  (.A1(\V2/A1/A1/A2/M2/c1 ),
    .A2(\V2/A1/A1/A2/M2/c2 ),
    .ZN(\V2/A1/A1/A2/c2 ));
 AND2_X1 \V2/A1/A1/A2/M3/M1/_0_  (.A1(\V2/v2 [6]),
    .A2(\V2/v3 [6]),
    .ZN(\V2/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M3/M1/_1_  (.A(\V2/v2 [6]),
    .B(\V2/v3 [6]),
    .Z(\V2/A1/A1/A2/M3/s1 ));
 AND2_X1 \V2/A1/A1/A2/M3/M2/_0_  (.A1(\V2/A1/A1/A2/M3/s1 ),
    .A2(\V2/A1/A1/A2/c2 ),
    .ZN(\V2/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M3/M2/_1_  (.A(\V2/A1/A1/A2/M3/s1 ),
    .B(\V2/A1/A1/A2/c2 ),
    .Z(\V2/s1 [6]));
 OR2_X1 \V2/A1/A1/A2/M3/_0_  (.A1(\V2/A1/A1/A2/M3/c1 ),
    .A2(\V2/A1/A1/A2/M3/c2 ),
    .ZN(\V2/A1/A1/A2/c3 ));
 AND2_X1 \V2/A1/A1/A2/M4/M1/_0_  (.A1(\V2/v2 [7]),
    .A2(\V2/v3 [7]),
    .ZN(\V2/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A1/A1/A2/M4/M1/_1_  (.A(\V2/v2 [7]),
    .B(\V2/v3 [7]),
    .Z(\V2/A1/A1/A2/M4/s1 ));
 AND2_X1 \V2/A1/A1/A2/M4/M2/_0_  (.A1(\V2/A1/A1/A2/M4/s1 ),
    .A2(\V2/A1/A1/A2/c3 ),
    .ZN(\V2/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A1/A1/A2/M4/M2/_1_  (.A(\V2/A1/A1/A2/M4/s1 ),
    .B(\V2/A1/A1/A2/c3 ),
    .Z(\V2/s1 [7]));
 OR2_X1 \V2/A1/A1/A2/M4/_0_  (.A1(\V2/A1/A1/A2/M4/c1 ),
    .A2(\V2/A1/A1/A2/M4/c2 ),
    .ZN(\V2/A1/c1 ));
 AND2_X1 \V2/A1/A2/A1/M1/M1/_0_  (.A1(\V2/v2 [8]),
    .A2(\V2/v3 [8]),
    .ZN(\V2/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M1/M1/_1_  (.A(\V2/v2 [8]),
    .B(\V2/v3 [8]),
    .Z(\V2/A1/A2/A1/M1/s1 ));
 AND2_X1 \V2/A1/A2/A1/M1/M2/_0_  (.A1(\V2/A1/A2/A1/M1/s1 ),
    .A2(\V2/A1/c1 ),
    .ZN(\V2/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M1/M2/_1_  (.A(\V2/A1/A2/A1/M1/s1 ),
    .B(\V2/A1/c1 ),
    .Z(\V2/s1 [8]));
 OR2_X1 \V2/A1/A2/A1/M1/_0_  (.A1(\V2/A1/A2/A1/M1/c1 ),
    .A2(\V2/A1/A2/A1/M1/c2 ),
    .ZN(\V2/A1/A2/A1/c1 ));
 AND2_X1 \V2/A1/A2/A1/M2/M1/_0_  (.A1(\V2/v2 [9]),
    .A2(\V2/v3 [9]),
    .ZN(\V2/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M2/M1/_1_  (.A(\V2/v2 [9]),
    .B(\V2/v3 [9]),
    .Z(\V2/A1/A2/A1/M2/s1 ));
 AND2_X1 \V2/A1/A2/A1/M2/M2/_0_  (.A1(\V2/A1/A2/A1/M2/s1 ),
    .A2(\V2/A1/A2/A1/c1 ),
    .ZN(\V2/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M2/M2/_1_  (.A(\V2/A1/A2/A1/M2/s1 ),
    .B(\V2/A1/A2/A1/c1 ),
    .Z(\V2/s1 [9]));
 OR2_X1 \V2/A1/A2/A1/M2/_0_  (.A1(\V2/A1/A2/A1/M2/c1 ),
    .A2(\V2/A1/A2/A1/M2/c2 ),
    .ZN(\V2/A1/A2/A1/c2 ));
 AND2_X1 \V2/A1/A2/A1/M3/M1/_0_  (.A1(\V2/v2 [10]),
    .A2(\V2/v3 [10]),
    .ZN(\V2/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M3/M1/_1_  (.A(\V2/v2 [10]),
    .B(\V2/v3 [10]),
    .Z(\V2/A1/A2/A1/M3/s1 ));
 AND2_X1 \V2/A1/A2/A1/M3/M2/_0_  (.A1(\V2/A1/A2/A1/M3/s1 ),
    .A2(\V2/A1/A2/A1/c2 ),
    .ZN(\V2/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M3/M2/_1_  (.A(\V2/A1/A2/A1/M3/s1 ),
    .B(\V2/A1/A2/A1/c2 ),
    .Z(\V2/s1 [10]));
 OR2_X1 \V2/A1/A2/A1/M3/_0_  (.A1(\V2/A1/A2/A1/M3/c1 ),
    .A2(\V2/A1/A2/A1/M3/c2 ),
    .ZN(\V2/A1/A2/A1/c3 ));
 AND2_X1 \V2/A1/A2/A1/M4/M1/_0_  (.A1(\V2/v2 [11]),
    .A2(\V2/v3 [11]),
    .ZN(\V2/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A1/A2/A1/M4/M1/_1_  (.A(\V2/v2 [11]),
    .B(\V2/v3 [11]),
    .Z(\V2/A1/A2/A1/M4/s1 ));
 AND2_X1 \V2/A1/A2/A1/M4/M2/_0_  (.A1(\V2/A1/A2/A1/M4/s1 ),
    .A2(\V2/A1/A2/A1/c3 ),
    .ZN(\V2/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A1/A2/A1/M4/M2/_1_  (.A(\V2/A1/A2/A1/M4/s1 ),
    .B(\V2/A1/A2/A1/c3 ),
    .Z(\V2/s1 [11]));
 OR2_X1 \V2/A1/A2/A1/M4/_0_  (.A1(\V2/A1/A2/A1/M4/c1 ),
    .A2(\V2/A1/A2/A1/M4/c2 ),
    .ZN(\V2/A1/A2/c1 ));
 AND2_X1 \V2/A1/A2/A2/M1/M1/_0_  (.A1(\V2/v2 [12]),
    .A2(\V2/v3 [12]),
    .ZN(\V2/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M1/M1/_1_  (.A(\V2/v2 [12]),
    .B(\V2/v3 [12]),
    .Z(\V2/A1/A2/A2/M1/s1 ));
 AND2_X1 \V2/A1/A2/A2/M1/M2/_0_  (.A1(\V2/A1/A2/A2/M1/s1 ),
    .A2(\V2/A1/A2/c1 ),
    .ZN(\V2/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M1/M2/_1_  (.A(\V2/A1/A2/A2/M1/s1 ),
    .B(\V2/A1/A2/c1 ),
    .Z(\V2/s1 [12]));
 OR2_X1 \V2/A1/A2/A2/M1/_0_  (.A1(\V2/A1/A2/A2/M1/c1 ),
    .A2(\V2/A1/A2/A2/M1/c2 ),
    .ZN(\V2/A1/A2/A2/c1 ));
 AND2_X1 \V2/A1/A2/A2/M2/M1/_0_  (.A1(\V2/v2 [13]),
    .A2(\V2/v3 [13]),
    .ZN(\V2/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M2/M1/_1_  (.A(\V2/v2 [13]),
    .B(\V2/v3 [13]),
    .Z(\V2/A1/A2/A2/M2/s1 ));
 AND2_X1 \V2/A1/A2/A2/M2/M2/_0_  (.A1(\V2/A1/A2/A2/M2/s1 ),
    .A2(\V2/A1/A2/A2/c1 ),
    .ZN(\V2/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M2/M2/_1_  (.A(\V2/A1/A2/A2/M2/s1 ),
    .B(\V2/A1/A2/A2/c1 ),
    .Z(\V2/s1 [13]));
 OR2_X1 \V2/A1/A2/A2/M2/_0_  (.A1(\V2/A1/A2/A2/M2/c1 ),
    .A2(\V2/A1/A2/A2/M2/c2 ),
    .ZN(\V2/A1/A2/A2/c2 ));
 AND2_X1 \V2/A1/A2/A2/M3/M1/_0_  (.A1(\V2/v2 [14]),
    .A2(\V2/v3 [14]),
    .ZN(\V2/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M3/M1/_1_  (.A(\V2/v2 [14]),
    .B(\V2/v3 [14]),
    .Z(\V2/A1/A2/A2/M3/s1 ));
 AND2_X1 \V2/A1/A2/A2/M3/M2/_0_  (.A1(\V2/A1/A2/A2/M3/s1 ),
    .A2(\V2/A1/A2/A2/c2 ),
    .ZN(\V2/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M3/M2/_1_  (.A(\V2/A1/A2/A2/M3/s1 ),
    .B(\V2/A1/A2/A2/c2 ),
    .Z(\V2/s1 [14]));
 OR2_X1 \V2/A1/A2/A2/M3/_0_  (.A1(\V2/A1/A2/A2/M3/c1 ),
    .A2(\V2/A1/A2/A2/M3/c2 ),
    .ZN(\V2/A1/A2/A2/c3 ));
 AND2_X1 \V2/A1/A2/A2/M4/M1/_0_  (.A1(\V2/v2 [15]),
    .A2(\V2/v3 [15]),
    .ZN(\V2/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A1/A2/A2/M4/M1/_1_  (.A(\V2/v2 [15]),
    .B(\V2/v3 [15]),
    .Z(\V2/A1/A2/A2/M4/s1 ));
 AND2_X1 \V2/A1/A2/A2/M4/M2/_0_  (.A1(\V2/A1/A2/A2/M4/s1 ),
    .A2(\V2/A1/A2/A2/c3 ),
    .ZN(\V2/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A1/A2/A2/M4/M2/_1_  (.A(\V2/A1/A2/A2/M4/s1 ),
    .B(\V2/A1/A2/A2/c3 ),
    .Z(\V2/s1 [15]));
 OR2_X1 \V2/A1/A2/A2/M4/_0_  (.A1(\V2/A1/A2/A2/M4/c1 ),
    .A2(\V2/A1/A2/A2/M4/c2 ),
    .ZN(\V2/c1 ));
 AND2_X1 \V2/A2/A1/A1/M1/M1/_0_  (.A1(\V2/s1 [0]),
    .A2(\V2/v1 [8]),
    .ZN(\V2/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M1/M1/_1_  (.A(\V2/s1 [0]),
    .B(\V2/v1 [8]),
    .Z(\V2/A2/A1/A1/M1/s1 ));
 AND2_X1 \V2/A2/A1/A1/M1/M2/_0_  (.A1(\V2/A2/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V2/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M1/M2/_1_  (.A(\V2/A2/A1/A1/M1/s1 ),
    .B(net6),
    .Z(v2[8]));
 OR2_X1 \V2/A2/A1/A1/M1/_0_  (.A1(\V2/A2/A1/A1/M1/c1 ),
    .A2(\V2/A2/A1/A1/M1/c2 ),
    .ZN(\V2/A2/A1/A1/c1 ));
 AND2_X1 \V2/A2/A1/A1/M2/M1/_0_  (.A1(\V2/s1 [1]),
    .A2(\V2/v1 [9]),
    .ZN(\V2/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M2/M1/_1_  (.A(\V2/s1 [1]),
    .B(\V2/v1 [9]),
    .Z(\V2/A2/A1/A1/M2/s1 ));
 AND2_X1 \V2/A2/A1/A1/M2/M2/_0_  (.A1(\V2/A2/A1/A1/M2/s1 ),
    .A2(\V2/A2/A1/A1/c1 ),
    .ZN(\V2/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M2/M2/_1_  (.A(\V2/A2/A1/A1/M2/s1 ),
    .B(\V2/A2/A1/A1/c1 ),
    .Z(v2[9]));
 OR2_X1 \V2/A2/A1/A1/M2/_0_  (.A1(\V2/A2/A1/A1/M2/c1 ),
    .A2(\V2/A2/A1/A1/M2/c2 ),
    .ZN(\V2/A2/A1/A1/c2 ));
 AND2_X1 \V2/A2/A1/A1/M3/M1/_0_  (.A1(\V2/s1 [2]),
    .A2(\V2/v1 [10]),
    .ZN(\V2/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M3/M1/_1_  (.A(\V2/s1 [2]),
    .B(\V2/v1 [10]),
    .Z(\V2/A2/A1/A1/M3/s1 ));
 AND2_X1 \V2/A2/A1/A1/M3/M2/_0_  (.A1(\V2/A2/A1/A1/M3/s1 ),
    .A2(\V2/A2/A1/A1/c2 ),
    .ZN(\V2/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M3/M2/_1_  (.A(\V2/A2/A1/A1/M3/s1 ),
    .B(\V2/A2/A1/A1/c2 ),
    .Z(v2[10]));
 OR2_X1 \V2/A2/A1/A1/M3/_0_  (.A1(\V2/A2/A1/A1/M3/c1 ),
    .A2(\V2/A2/A1/A1/M3/c2 ),
    .ZN(\V2/A2/A1/A1/c3 ));
 AND2_X1 \V2/A2/A1/A1/M4/M1/_0_  (.A1(\V2/s1 [3]),
    .A2(\V2/v1 [11]),
    .ZN(\V2/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A2/A1/A1/M4/M1/_1_  (.A(\V2/s1 [3]),
    .B(\V2/v1 [11]),
    .Z(\V2/A2/A1/A1/M4/s1 ));
 AND2_X1 \V2/A2/A1/A1/M4/M2/_0_  (.A1(\V2/A2/A1/A1/M4/s1 ),
    .A2(\V2/A2/A1/A1/c3 ),
    .ZN(\V2/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A2/A1/A1/M4/M2/_1_  (.A(\V2/A2/A1/A1/M4/s1 ),
    .B(\V2/A2/A1/A1/c3 ),
    .Z(v2[11]));
 OR2_X1 \V2/A2/A1/A1/M4/_0_  (.A1(\V2/A2/A1/A1/M4/c1 ),
    .A2(\V2/A2/A1/A1/M4/c2 ),
    .ZN(\V2/A2/A1/c1 ));
 AND2_X1 \V2/A2/A1/A2/M1/M1/_0_  (.A1(\V2/s1 [4]),
    .A2(\V2/v1 [12]),
    .ZN(\V2/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M1/M1/_1_  (.A(\V2/s1 [4]),
    .B(\V2/v1 [12]),
    .Z(\V2/A2/A1/A2/M1/s1 ));
 AND2_X1 \V2/A2/A1/A2/M1/M2/_0_  (.A1(\V2/A2/A1/A2/M1/s1 ),
    .A2(\V2/A2/A1/c1 ),
    .ZN(\V2/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M1/M2/_1_  (.A(\V2/A2/A1/A2/M1/s1 ),
    .B(\V2/A2/A1/c1 ),
    .Z(v2[12]));
 OR2_X1 \V2/A2/A1/A2/M1/_0_  (.A1(\V2/A2/A1/A2/M1/c1 ),
    .A2(\V2/A2/A1/A2/M1/c2 ),
    .ZN(\V2/A2/A1/A2/c1 ));
 AND2_X1 \V2/A2/A1/A2/M2/M1/_0_  (.A1(\V2/s1 [5]),
    .A2(\V2/v1 [13]),
    .ZN(\V2/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M2/M1/_1_  (.A(\V2/s1 [5]),
    .B(\V2/v1 [13]),
    .Z(\V2/A2/A1/A2/M2/s1 ));
 AND2_X1 \V2/A2/A1/A2/M2/M2/_0_  (.A1(\V2/A2/A1/A2/M2/s1 ),
    .A2(\V2/A2/A1/A2/c1 ),
    .ZN(\V2/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M2/M2/_1_  (.A(\V2/A2/A1/A2/M2/s1 ),
    .B(\V2/A2/A1/A2/c1 ),
    .Z(v2[13]));
 OR2_X1 \V2/A2/A1/A2/M2/_0_  (.A1(\V2/A2/A1/A2/M2/c1 ),
    .A2(\V2/A2/A1/A2/M2/c2 ),
    .ZN(\V2/A2/A1/A2/c2 ));
 AND2_X1 \V2/A2/A1/A2/M3/M1/_0_  (.A1(\V2/s1 [6]),
    .A2(\V2/v1 [14]),
    .ZN(\V2/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M3/M1/_1_  (.A(\V2/s1 [6]),
    .B(\V2/v1 [14]),
    .Z(\V2/A2/A1/A2/M3/s1 ));
 AND2_X1 \V2/A2/A1/A2/M3/M2/_0_  (.A1(\V2/A2/A1/A2/M3/s1 ),
    .A2(\V2/A2/A1/A2/c2 ),
    .ZN(\V2/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M3/M2/_1_  (.A(\V2/A2/A1/A2/M3/s1 ),
    .B(\V2/A2/A1/A2/c2 ),
    .Z(v2[14]));
 OR2_X1 \V2/A2/A1/A2/M3/_0_  (.A1(\V2/A2/A1/A2/M3/c1 ),
    .A2(\V2/A2/A1/A2/M3/c2 ),
    .ZN(\V2/A2/A1/A2/c3 ));
 AND2_X1 \V2/A2/A1/A2/M4/M1/_0_  (.A1(\V2/s1 [7]),
    .A2(\V2/v1 [15]),
    .ZN(\V2/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A2/A1/A2/M4/M1/_1_  (.A(\V2/s1 [7]),
    .B(\V2/v1 [15]),
    .Z(\V2/A2/A1/A2/M4/s1 ));
 AND2_X1 \V2/A2/A1/A2/M4/M2/_0_  (.A1(\V2/A2/A1/A2/M4/s1 ),
    .A2(\V2/A2/A1/A2/c3 ),
    .ZN(\V2/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A2/A1/A2/M4/M2/_1_  (.A(\V2/A2/A1/A2/M4/s1 ),
    .B(\V2/A2/A1/A2/c3 ),
    .Z(v2[15]));
 OR2_X1 \V2/A2/A1/A2/M4/_0_  (.A1(\V2/A2/A1/A2/M4/c1 ),
    .A2(\V2/A2/A1/A2/M4/c2 ),
    .ZN(\V2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A1/M1/M1/_0_  (.A1(\V2/s1 [8]),
    .A2(net7),
    .ZN(\V2/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M1/M1/_1_  (.A(\V2/s1 [8]),
    .B(net7),
    .Z(\V2/A2/A2/A1/M1/s1 ));
 AND2_X1 \V2/A2/A2/A1/M1/M2/_0_  (.A1(\V2/A2/A2/A1/M1/s1 ),
    .A2(\V2/A2/c1 ),
    .ZN(\V2/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M1/M2/_1_  (.A(\V2/A2/A2/A1/M1/s1 ),
    .B(\V2/A2/c1 ),
    .Z(\V2/s2 [8]));
 OR2_X1 \V2/A2/A2/A1/M1/_0_  (.A1(\V2/A2/A2/A1/M1/c1 ),
    .A2(\V2/A2/A2/A1/M1/c2 ),
    .ZN(\V2/A2/A2/A1/c1 ));
 AND2_X1 \V2/A2/A2/A1/M2/M1/_0_  (.A1(\V2/s1 [9]),
    .A2(net7),
    .ZN(\V2/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M2/M1/_1_  (.A(\V2/s1 [9]),
    .B(net7),
    .Z(\V2/A2/A2/A1/M2/s1 ));
 AND2_X1 \V2/A2/A2/A1/M2/M2/_0_  (.A1(\V2/A2/A2/A1/M2/s1 ),
    .A2(\V2/A2/A2/A1/c1 ),
    .ZN(\V2/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M2/M2/_1_  (.A(\V2/A2/A2/A1/M2/s1 ),
    .B(\V2/A2/A2/A1/c1 ),
    .Z(\V2/s2 [9]));
 OR2_X1 \V2/A2/A2/A1/M2/_0_  (.A1(\V2/A2/A2/A1/M2/c1 ),
    .A2(\V2/A2/A2/A1/M2/c2 ),
    .ZN(\V2/A2/A2/A1/c2 ));
 AND2_X1 \V2/A2/A2/A1/M3/M1/_0_  (.A1(\V2/s1 [10]),
    .A2(net7),
    .ZN(\V2/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M3/M1/_1_  (.A(\V2/s1 [10]),
    .B(net7),
    .Z(\V2/A2/A2/A1/M3/s1 ));
 AND2_X1 \V2/A2/A2/A1/M3/M2/_0_  (.A1(\V2/A2/A2/A1/M3/s1 ),
    .A2(\V2/A2/A2/A1/c2 ),
    .ZN(\V2/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M3/M2/_1_  (.A(\V2/A2/A2/A1/M3/s1 ),
    .B(\V2/A2/A2/A1/c2 ),
    .Z(\V2/s2 [10]));
 OR2_X1 \V2/A2/A2/A1/M3/_0_  (.A1(\V2/A2/A2/A1/M3/c1 ),
    .A2(\V2/A2/A2/A1/M3/c2 ),
    .ZN(\V2/A2/A2/A1/c3 ));
 AND2_X1 \V2/A2/A2/A1/M4/M1/_0_  (.A1(\V2/s1 [11]),
    .A2(net7),
    .ZN(\V2/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A2/A2/A1/M4/M1/_1_  (.A(\V2/s1 [11]),
    .B(net7),
    .Z(\V2/A2/A2/A1/M4/s1 ));
 AND2_X1 \V2/A2/A2/A1/M4/M2/_0_  (.A1(\V2/A2/A2/A1/M4/s1 ),
    .A2(\V2/A2/A2/A1/c3 ),
    .ZN(\V2/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A2/A2/A1/M4/M2/_1_  (.A(\V2/A2/A2/A1/M4/s1 ),
    .B(\V2/A2/A2/A1/c3 ),
    .Z(\V2/s2 [11]));
 OR2_X1 \V2/A2/A2/A1/M4/_0_  (.A1(\V2/A2/A2/A1/M4/c1 ),
    .A2(\V2/A2/A2/A1/M4/c2 ),
    .ZN(\V2/A2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A2/M1/M1/_0_  (.A1(\V2/s1 [12]),
    .A2(net7),
    .ZN(\V2/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M1/M1/_1_  (.A(\V2/s1 [12]),
    .B(net7),
    .Z(\V2/A2/A2/A2/M1/s1 ));
 AND2_X1 \V2/A2/A2/A2/M1/M2/_0_  (.A1(\V2/A2/A2/A2/M1/s1 ),
    .A2(\V2/A2/A2/c1 ),
    .ZN(\V2/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M1/M2/_1_  (.A(\V2/A2/A2/A2/M1/s1 ),
    .B(\V2/A2/A2/c1 ),
    .Z(\V2/s2 [12]));
 OR2_X1 \V2/A2/A2/A2/M1/_0_  (.A1(\V2/A2/A2/A2/M1/c1 ),
    .A2(\V2/A2/A2/A2/M1/c2 ),
    .ZN(\V2/A2/A2/A2/c1 ));
 AND2_X1 \V2/A2/A2/A2/M2/M1/_0_  (.A1(\V2/s1 [13]),
    .A2(net7),
    .ZN(\V2/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M2/M1/_1_  (.A(\V2/s1 [13]),
    .B(net7),
    .Z(\V2/A2/A2/A2/M2/s1 ));
 AND2_X1 \V2/A2/A2/A2/M2/M2/_0_  (.A1(\V2/A2/A2/A2/M2/s1 ),
    .A2(\V2/A2/A2/A2/c1 ),
    .ZN(\V2/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M2/M2/_1_  (.A(\V2/A2/A2/A2/M2/s1 ),
    .B(\V2/A2/A2/A2/c1 ),
    .Z(\V2/s2 [13]));
 OR2_X1 \V2/A2/A2/A2/M2/_0_  (.A1(\V2/A2/A2/A2/M2/c1 ),
    .A2(\V2/A2/A2/A2/M2/c2 ),
    .ZN(\V2/A2/A2/A2/c2 ));
 AND2_X1 \V2/A2/A2/A2/M3/M1/_0_  (.A1(\V2/s1 [14]),
    .A2(net7),
    .ZN(\V2/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M3/M1/_1_  (.A(\V2/s1 [14]),
    .B(net7),
    .Z(\V2/A2/A2/A2/M3/s1 ));
 AND2_X1 \V2/A2/A2/A2/M3/M2/_0_  (.A1(\V2/A2/A2/A2/M3/s1 ),
    .A2(\V2/A2/A2/A2/c2 ),
    .ZN(\V2/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M3/M2/_1_  (.A(\V2/A2/A2/A2/M3/s1 ),
    .B(\V2/A2/A2/A2/c2 ),
    .Z(\V2/s2 [14]));
 OR2_X1 \V2/A2/A2/A2/M3/_0_  (.A1(\V2/A2/A2/A2/M3/c1 ),
    .A2(\V2/A2/A2/A2/M3/c2 ),
    .ZN(\V2/A2/A2/A2/c3 ));
 AND2_X1 \V2/A2/A2/A2/M4/M1/_0_  (.A1(\V2/s1 [15]),
    .A2(net7),
    .ZN(\V2/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A2/A2/A2/M4/M1/_1_  (.A(\V2/s1 [15]),
    .B(net7),
    .Z(\V2/A2/A2/A2/M4/s1 ));
 AND2_X1 \V2/A2/A2/A2/M4/M2/_0_  (.A1(\V2/A2/A2/A2/M4/s1 ),
    .A2(\V2/A2/A2/A2/c3 ),
    .ZN(\V2/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A2/A2/A2/M4/M2/_1_  (.A(\V2/A2/A2/A2/M4/s1 ),
    .B(\V2/A2/A2/A2/c3 ),
    .Z(\V2/s2 [15]));
 OR2_X1 \V2/A2/A2/A2/M4/_0_  (.A1(\V2/A2/A2/A2/M4/c1 ),
    .A2(\V2/A2/A2/A2/M4/c2 ),
    .ZN(\V2/c2 ));
 AND2_X1 \V2/A3/A1/A1/M1/M1/_0_  (.A1(\V2/v4 [0]),
    .A2(\V2/s2 [8]),
    .ZN(\V2/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M1/M1/_1_  (.A(\V2/v4 [0]),
    .B(\V2/s2 [8]),
    .Z(\V2/A3/A1/A1/M1/s1 ));
 AND2_X1 \V2/A3/A1/A1/M1/M2/_0_  (.A1(\V2/A3/A1/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M1/M2/_1_  (.A(\V2/A3/A1/A1/M1/s1 ),
    .B(net7),
    .Z(v2[16]));
 OR2_X1 \V2/A3/A1/A1/M1/_0_  (.A1(\V2/A3/A1/A1/M1/c1 ),
    .A2(\V2/A3/A1/A1/M1/c2 ),
    .ZN(\V2/A3/A1/A1/c1 ));
 AND2_X1 \V2/A3/A1/A1/M2/M1/_0_  (.A1(\V2/v4 [1]),
    .A2(\V2/s2 [9]),
    .ZN(\V2/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M2/M1/_1_  (.A(\V2/v4 [1]),
    .B(\V2/s2 [9]),
    .Z(\V2/A3/A1/A1/M2/s1 ));
 AND2_X1 \V2/A3/A1/A1/M2/M2/_0_  (.A1(\V2/A3/A1/A1/M2/s1 ),
    .A2(\V2/A3/A1/A1/c1 ),
    .ZN(\V2/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M2/M2/_1_  (.A(\V2/A3/A1/A1/M2/s1 ),
    .B(\V2/A3/A1/A1/c1 ),
    .Z(v2[17]));
 OR2_X1 \V2/A3/A1/A1/M2/_0_  (.A1(\V2/A3/A1/A1/M2/c1 ),
    .A2(\V2/A3/A1/A1/M2/c2 ),
    .ZN(\V2/A3/A1/A1/c2 ));
 AND2_X1 \V2/A3/A1/A1/M3/M1/_0_  (.A1(\V2/v4 [2]),
    .A2(\V2/s2 [10]),
    .ZN(\V2/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M3/M1/_1_  (.A(\V2/v4 [2]),
    .B(\V2/s2 [10]),
    .Z(\V2/A3/A1/A1/M3/s1 ));
 AND2_X1 \V2/A3/A1/A1/M3/M2/_0_  (.A1(\V2/A3/A1/A1/M3/s1 ),
    .A2(\V2/A3/A1/A1/c2 ),
    .ZN(\V2/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M3/M2/_1_  (.A(\V2/A3/A1/A1/M3/s1 ),
    .B(\V2/A3/A1/A1/c2 ),
    .Z(v2[18]));
 OR2_X1 \V2/A3/A1/A1/M3/_0_  (.A1(\V2/A3/A1/A1/M3/c1 ),
    .A2(\V2/A3/A1/A1/M3/c2 ),
    .ZN(\V2/A3/A1/A1/c3 ));
 AND2_X1 \V2/A3/A1/A1/M4/M1/_0_  (.A1(\V2/v4 [3]),
    .A2(\V2/s2 [11]),
    .ZN(\V2/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V2/A3/A1/A1/M4/M1/_1_  (.A(\V2/v4 [3]),
    .B(\V2/s2 [11]),
    .Z(\V2/A3/A1/A1/M4/s1 ));
 AND2_X1 \V2/A3/A1/A1/M4/M2/_0_  (.A1(\V2/A3/A1/A1/M4/s1 ),
    .A2(\V2/A3/A1/A1/c3 ),
    .ZN(\V2/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V2/A3/A1/A1/M4/M2/_1_  (.A(\V2/A3/A1/A1/M4/s1 ),
    .B(\V2/A3/A1/A1/c3 ),
    .Z(v2[19]));
 OR2_X1 \V2/A3/A1/A1/M4/_0_  (.A1(\V2/A3/A1/A1/M4/c1 ),
    .A2(\V2/A3/A1/A1/M4/c2 ),
    .ZN(\V2/A3/A1/c1 ));
 AND2_X1 \V2/A3/A1/A2/M1/M1/_0_  (.A1(\V2/v4 [4]),
    .A2(\V2/s2 [12]),
    .ZN(\V2/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M1/M1/_1_  (.A(\V2/v4 [4]),
    .B(\V2/s2 [12]),
    .Z(\V2/A3/A1/A2/M1/s1 ));
 AND2_X1 \V2/A3/A1/A2/M1/M2/_0_  (.A1(\V2/A3/A1/A2/M1/s1 ),
    .A2(\V2/A3/A1/c1 ),
    .ZN(\V2/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M1/M2/_1_  (.A(\V2/A3/A1/A2/M1/s1 ),
    .B(\V2/A3/A1/c1 ),
    .Z(v2[20]));
 OR2_X1 \V2/A3/A1/A2/M1/_0_  (.A1(\V2/A3/A1/A2/M1/c1 ),
    .A2(\V2/A3/A1/A2/M1/c2 ),
    .ZN(\V2/A3/A1/A2/c1 ));
 AND2_X1 \V2/A3/A1/A2/M2/M1/_0_  (.A1(\V2/v4 [5]),
    .A2(\V2/s2 [13]),
    .ZN(\V2/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M2/M1/_1_  (.A(\V2/v4 [5]),
    .B(\V2/s2 [13]),
    .Z(\V2/A3/A1/A2/M2/s1 ));
 AND2_X1 \V2/A3/A1/A2/M2/M2/_0_  (.A1(\V2/A3/A1/A2/M2/s1 ),
    .A2(\V2/A3/A1/A2/c1 ),
    .ZN(\V2/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M2/M2/_1_  (.A(\V2/A3/A1/A2/M2/s1 ),
    .B(\V2/A3/A1/A2/c1 ),
    .Z(v2[21]));
 OR2_X1 \V2/A3/A1/A2/M2/_0_  (.A1(\V2/A3/A1/A2/M2/c1 ),
    .A2(\V2/A3/A1/A2/M2/c2 ),
    .ZN(\V2/A3/A1/A2/c2 ));
 AND2_X1 \V2/A3/A1/A2/M3/M1/_0_  (.A1(\V2/v4 [6]),
    .A2(\V2/s2 [14]),
    .ZN(\V2/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M3/M1/_1_  (.A(\V2/v4 [6]),
    .B(\V2/s2 [14]),
    .Z(\V2/A3/A1/A2/M3/s1 ));
 AND2_X1 \V2/A3/A1/A2/M3/M2/_0_  (.A1(\V2/A3/A1/A2/M3/s1 ),
    .A2(\V2/A3/A1/A2/c2 ),
    .ZN(\V2/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M3/M2/_1_  (.A(\V2/A3/A1/A2/M3/s1 ),
    .B(\V2/A3/A1/A2/c2 ),
    .Z(v2[22]));
 OR2_X1 \V2/A3/A1/A2/M3/_0_  (.A1(\V2/A3/A1/A2/M3/c1 ),
    .A2(\V2/A3/A1/A2/M3/c2 ),
    .ZN(\V2/A3/A1/A2/c3 ));
 AND2_X1 \V2/A3/A1/A2/M4/M1/_0_  (.A1(\V2/v4 [7]),
    .A2(\V2/s2 [15]),
    .ZN(\V2/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V2/A3/A1/A2/M4/M1/_1_  (.A(\V2/v4 [7]),
    .B(\V2/s2 [15]),
    .Z(\V2/A3/A1/A2/M4/s1 ));
 AND2_X1 \V2/A3/A1/A2/M4/M2/_0_  (.A1(\V2/A3/A1/A2/M4/s1 ),
    .A2(\V2/A3/A1/A2/c3 ),
    .ZN(\V2/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V2/A3/A1/A2/M4/M2/_1_  (.A(\V2/A3/A1/A2/M4/s1 ),
    .B(\V2/A3/A1/A2/c3 ),
    .Z(v2[23]));
 OR2_X1 \V2/A3/A1/A2/M4/_0_  (.A1(\V2/A3/A1/A2/M4/c1 ),
    .A2(\V2/A3/A1/A2/M4/c2 ),
    .ZN(\V2/A3/c1 ));
 AND2_X1 \V2/A3/A2/A1/M1/M1/_0_  (.A1(\V2/v4 [8]),
    .A2(\V2/c3 ),
    .ZN(\V2/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M1/M1/_1_  (.A(\V2/v4 [8]),
    .B(\V2/c3 ),
    .Z(\V2/A3/A2/A1/M1/s1 ));
 AND2_X1 \V2/A3/A2/A1/M1/M2/_0_  (.A1(\V2/A3/A2/A1/M1/s1 ),
    .A2(\V2/A3/c1 ),
    .ZN(\V2/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M1/M2/_1_  (.A(\V2/A3/A2/A1/M1/s1 ),
    .B(\V2/A3/c1 ),
    .Z(v2[24]));
 OR2_X1 \V2/A3/A2/A1/M1/_0_  (.A1(\V2/A3/A2/A1/M1/c1 ),
    .A2(\V2/A3/A2/A1/M1/c2 ),
    .ZN(\V2/A3/A2/A1/c1 ));
 AND2_X1 \V2/A3/A2/A1/M2/M1/_0_  (.A1(\V2/v4 [9]),
    .A2(net7),
    .ZN(\V2/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M2/M1/_1_  (.A(\V2/v4 [9]),
    .B(net7),
    .Z(\V2/A3/A2/A1/M2/s1 ));
 AND2_X1 \V2/A3/A2/A1/M2/M2/_0_  (.A1(\V2/A3/A2/A1/M2/s1 ),
    .A2(\V2/A3/A2/A1/c1 ),
    .ZN(\V2/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M2/M2/_1_  (.A(\V2/A3/A2/A1/M2/s1 ),
    .B(\V2/A3/A2/A1/c1 ),
    .Z(v2[25]));
 OR2_X1 \V2/A3/A2/A1/M2/_0_  (.A1(\V2/A3/A2/A1/M2/c1 ),
    .A2(\V2/A3/A2/A1/M2/c2 ),
    .ZN(\V2/A3/A2/A1/c2 ));
 AND2_X1 \V2/A3/A2/A1/M3/M1/_0_  (.A1(\V2/v4 [10]),
    .A2(net7),
    .ZN(\V2/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M3/M1/_1_  (.A(\V2/v4 [10]),
    .B(net7),
    .Z(\V2/A3/A2/A1/M3/s1 ));
 AND2_X1 \V2/A3/A2/A1/M3/M2/_0_  (.A1(\V2/A3/A2/A1/M3/s1 ),
    .A2(\V2/A3/A2/A1/c2 ),
    .ZN(\V2/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M3/M2/_1_  (.A(\V2/A3/A2/A1/M3/s1 ),
    .B(\V2/A3/A2/A1/c2 ),
    .Z(v2[26]));
 OR2_X1 \V2/A3/A2/A1/M3/_0_  (.A1(\V2/A3/A2/A1/M3/c1 ),
    .A2(\V2/A3/A2/A1/M3/c2 ),
    .ZN(\V2/A3/A2/A1/c3 ));
 AND2_X1 \V2/A3/A2/A1/M4/M1/_0_  (.A1(\V2/v4 [11]),
    .A2(net7),
    .ZN(\V2/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V2/A3/A2/A1/M4/M1/_1_  (.A(\V2/v4 [11]),
    .B(net7),
    .Z(\V2/A3/A2/A1/M4/s1 ));
 AND2_X1 \V2/A3/A2/A1/M4/M2/_0_  (.A1(\V2/A3/A2/A1/M4/s1 ),
    .A2(\V2/A3/A2/A1/c3 ),
    .ZN(\V2/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V2/A3/A2/A1/M4/M2/_1_  (.A(\V2/A3/A2/A1/M4/s1 ),
    .B(\V2/A3/A2/A1/c3 ),
    .Z(v2[27]));
 OR2_X1 \V2/A3/A2/A1/M4/_0_  (.A1(\V2/A3/A2/A1/M4/c1 ),
    .A2(\V2/A3/A2/A1/M4/c2 ),
    .ZN(\V2/A3/A2/c1 ));
 AND2_X1 \V2/A3/A2/A2/M1/M1/_0_  (.A1(\V2/v4 [12]),
    .A2(net7),
    .ZN(\V2/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M1/M1/_1_  (.A(\V2/v4 [12]),
    .B(net7),
    .Z(\V2/A3/A2/A2/M1/s1 ));
 AND2_X1 \V2/A3/A2/A2/M1/M2/_0_  (.A1(\V2/A3/A2/A2/M1/s1 ),
    .A2(\V2/A3/A2/c1 ),
    .ZN(\V2/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M1/M2/_1_  (.A(\V2/A3/A2/A2/M1/s1 ),
    .B(\V2/A3/A2/c1 ),
    .Z(v2[28]));
 OR2_X1 \V2/A3/A2/A2/M1/_0_  (.A1(\V2/A3/A2/A2/M1/c1 ),
    .A2(\V2/A3/A2/A2/M1/c2 ),
    .ZN(\V2/A3/A2/A2/c1 ));
 AND2_X1 \V2/A3/A2/A2/M2/M1/_0_  (.A1(\V2/v4 [13]),
    .A2(net7),
    .ZN(\V2/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M2/M1/_1_  (.A(\V2/v4 [13]),
    .B(net7),
    .Z(\V2/A3/A2/A2/M2/s1 ));
 AND2_X1 \V2/A3/A2/A2/M2/M2/_0_  (.A1(\V2/A3/A2/A2/M2/s1 ),
    .A2(\V2/A3/A2/A2/c1 ),
    .ZN(\V2/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M2/M2/_1_  (.A(\V2/A3/A2/A2/M2/s1 ),
    .B(\V2/A3/A2/A2/c1 ),
    .Z(v2[29]));
 OR2_X1 \V2/A3/A2/A2/M2/_0_  (.A1(\V2/A3/A2/A2/M2/c1 ),
    .A2(\V2/A3/A2/A2/M2/c2 ),
    .ZN(\V2/A3/A2/A2/c2 ));
 AND2_X1 \V2/A3/A2/A2/M3/M1/_0_  (.A1(\V2/v4 [14]),
    .A2(net7),
    .ZN(\V2/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M3/M1/_1_  (.A(\V2/v4 [14]),
    .B(net7),
    .Z(\V2/A3/A2/A2/M3/s1 ));
 AND2_X1 \V2/A3/A2/A2/M3/M2/_0_  (.A1(\V2/A3/A2/A2/M3/s1 ),
    .A2(\V2/A3/A2/A2/c2 ),
    .ZN(\V2/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M3/M2/_1_  (.A(\V2/A3/A2/A2/M3/s1 ),
    .B(\V2/A3/A2/A2/c2 ),
    .Z(v2[30]));
 OR2_X1 \V2/A3/A2/A2/M3/_0_  (.A1(\V2/A3/A2/A2/M3/c1 ),
    .A2(\V2/A3/A2/A2/M3/c2 ),
    .ZN(\V2/A3/A2/A2/c3 ));
 AND2_X1 \V2/A3/A2/A2/M4/M1/_0_  (.A1(\V2/v4 [15]),
    .A2(net7),
    .ZN(\V2/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V2/A3/A2/A2/M4/M1/_1_  (.A(\V2/v4 [15]),
    .B(net7),
    .Z(\V2/A3/A2/A2/M4/s1 ));
 AND2_X1 \V2/A3/A2/A2/M4/M2/_0_  (.A1(\V2/A3/A2/A2/M4/s1 ),
    .A2(\V2/A3/A2/A2/c3 ),
    .ZN(\V2/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V2/A3/A2/A2/M4/M2/_1_  (.A(\V2/A3/A2/A2/M4/s1 ),
    .B(\V2/A3/A2/A2/c3 ),
    .Z(v2[31]));
 OR2_X1 \V2/A3/A2/A2/M4/_0_  (.A1(\V2/A3/A2/A2/M4/c1 ),
    .A2(\V2/A3/A2/A2/M4/c2 ),
    .ZN(\V2/overflow ));
 AND2_X1 \V2/V1/A1/A1/M1/M1/_0_  (.A1(\V2/V1/v2 [0]),
    .A2(\V2/V1/v3 [0]),
    .ZN(\V2/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M1/M1/_1_  (.A(\V2/V1/v2 [0]),
    .B(\V2/V1/v3 [0]),
    .Z(\V2/V1/A1/A1/M1/s1 ));
 AND2_X1 \V2/V1/A1/A1/M1/M2/_0_  (.A1(\V2/V1/A1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M1/M2/_1_  (.A(\V2/V1/A1/A1/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/s1 [0]));
 OR2_X1 \V2/V1/A1/A1/M1/_0_  (.A1(\V2/V1/A1/A1/M1/c1 ),
    .A2(\V2/V1/A1/A1/M1/c2 ),
    .ZN(\V2/V1/A1/A1/c1 ));
 AND2_X1 \V2/V1/A1/A1/M2/M1/_0_  (.A1(\V2/V1/v2 [1]),
    .A2(\V2/V1/v3 [1]),
    .ZN(\V2/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M2/M1/_1_  (.A(\V2/V1/v2 [1]),
    .B(\V2/V1/v3 [1]),
    .Z(\V2/V1/A1/A1/M2/s1 ));
 AND2_X1 \V2/V1/A1/A1/M2/M2/_0_  (.A1(\V2/V1/A1/A1/M2/s1 ),
    .A2(\V2/V1/A1/A1/c1 ),
    .ZN(\V2/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M2/M2/_1_  (.A(\V2/V1/A1/A1/M2/s1 ),
    .B(\V2/V1/A1/A1/c1 ),
    .Z(\V2/V1/s1 [1]));
 OR2_X1 \V2/V1/A1/A1/M2/_0_  (.A1(\V2/V1/A1/A1/M2/c1 ),
    .A2(\V2/V1/A1/A1/M2/c2 ),
    .ZN(\V2/V1/A1/A1/c2 ));
 AND2_X1 \V2/V1/A1/A1/M3/M1/_0_  (.A1(\V2/V1/v2 [2]),
    .A2(\V2/V1/v3 [2]),
    .ZN(\V2/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M3/M1/_1_  (.A(\V2/V1/v2 [2]),
    .B(\V2/V1/v3 [2]),
    .Z(\V2/V1/A1/A1/M3/s1 ));
 AND2_X1 \V2/V1/A1/A1/M3/M2/_0_  (.A1(\V2/V1/A1/A1/M3/s1 ),
    .A2(\V2/V1/A1/A1/c2 ),
    .ZN(\V2/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M3/M2/_1_  (.A(\V2/V1/A1/A1/M3/s1 ),
    .B(\V2/V1/A1/A1/c2 ),
    .Z(\V2/V1/s1 [2]));
 OR2_X1 \V2/V1/A1/A1/M3/_0_  (.A1(\V2/V1/A1/A1/M3/c1 ),
    .A2(\V2/V1/A1/A1/M3/c2 ),
    .ZN(\V2/V1/A1/A1/c3 ));
 AND2_X1 \V2/V1/A1/A1/M4/M1/_0_  (.A1(\V2/V1/v2 [3]),
    .A2(\V2/V1/v3 [3]),
    .ZN(\V2/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A1/A1/M4/M1/_1_  (.A(\V2/V1/v2 [3]),
    .B(\V2/V1/v3 [3]),
    .Z(\V2/V1/A1/A1/M4/s1 ));
 AND2_X1 \V2/V1/A1/A1/M4/M2/_0_  (.A1(\V2/V1/A1/A1/M4/s1 ),
    .A2(\V2/V1/A1/A1/c3 ),
    .ZN(\V2/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A1/A1/M4/M2/_1_  (.A(\V2/V1/A1/A1/M4/s1 ),
    .B(\V2/V1/A1/A1/c3 ),
    .Z(\V2/V1/s1 [3]));
 OR2_X1 \V2/V1/A1/A1/M4/_0_  (.A1(\V2/V1/A1/A1/M4/c1 ),
    .A2(\V2/V1/A1/A1/M4/c2 ),
    .ZN(\V2/V1/A1/c1 ));
 AND2_X1 \V2/V1/A1/A2/M1/M1/_0_  (.A1(\V2/V1/v2 [4]),
    .A2(\V2/V1/v3 [4]),
    .ZN(\V2/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M1/M1/_1_  (.A(\V2/V1/v2 [4]),
    .B(\V2/V1/v3 [4]),
    .Z(\V2/V1/A1/A2/M1/s1 ));
 AND2_X1 \V2/V1/A1/A2/M1/M2/_0_  (.A1(\V2/V1/A1/A2/M1/s1 ),
    .A2(\V2/V1/A1/c1 ),
    .ZN(\V2/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M1/M2/_1_  (.A(\V2/V1/A1/A2/M1/s1 ),
    .B(\V2/V1/A1/c1 ),
    .Z(\V2/V1/s1 [4]));
 OR2_X1 \V2/V1/A1/A2/M1/_0_  (.A1(\V2/V1/A1/A2/M1/c1 ),
    .A2(\V2/V1/A1/A2/M1/c2 ),
    .ZN(\V2/V1/A1/A2/c1 ));
 AND2_X1 \V2/V1/A1/A2/M2/M1/_0_  (.A1(\V2/V1/v2 [5]),
    .A2(\V2/V1/v3 [5]),
    .ZN(\V2/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M2/M1/_1_  (.A(\V2/V1/v2 [5]),
    .B(\V2/V1/v3 [5]),
    .Z(\V2/V1/A1/A2/M2/s1 ));
 AND2_X1 \V2/V1/A1/A2/M2/M2/_0_  (.A1(\V2/V1/A1/A2/M2/s1 ),
    .A2(\V2/V1/A1/A2/c1 ),
    .ZN(\V2/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M2/M2/_1_  (.A(\V2/V1/A1/A2/M2/s1 ),
    .B(\V2/V1/A1/A2/c1 ),
    .Z(\V2/V1/s1 [5]));
 OR2_X1 \V2/V1/A1/A2/M2/_0_  (.A1(\V2/V1/A1/A2/M2/c1 ),
    .A2(\V2/V1/A1/A2/M2/c2 ),
    .ZN(\V2/V1/A1/A2/c2 ));
 AND2_X1 \V2/V1/A1/A2/M3/M1/_0_  (.A1(\V2/V1/v2 [6]),
    .A2(\V2/V1/v3 [6]),
    .ZN(\V2/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M3/M1/_1_  (.A(\V2/V1/v2 [6]),
    .B(\V2/V1/v3 [6]),
    .Z(\V2/V1/A1/A2/M3/s1 ));
 AND2_X1 \V2/V1/A1/A2/M3/M2/_0_  (.A1(\V2/V1/A1/A2/M3/s1 ),
    .A2(\V2/V1/A1/A2/c2 ),
    .ZN(\V2/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M3/M2/_1_  (.A(\V2/V1/A1/A2/M3/s1 ),
    .B(\V2/V1/A1/A2/c2 ),
    .Z(\V2/V1/s1 [6]));
 OR2_X1 \V2/V1/A1/A2/M3/_0_  (.A1(\V2/V1/A1/A2/M3/c1 ),
    .A2(\V2/V1/A1/A2/M3/c2 ),
    .ZN(\V2/V1/A1/A2/c3 ));
 AND2_X1 \V2/V1/A1/A2/M4/M1/_0_  (.A1(\V2/V1/v2 [7]),
    .A2(\V2/V1/v3 [7]),
    .ZN(\V2/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A1/A2/M4/M1/_1_  (.A(\V2/V1/v2 [7]),
    .B(\V2/V1/v3 [7]),
    .Z(\V2/V1/A1/A2/M4/s1 ));
 AND2_X1 \V2/V1/A1/A2/M4/M2/_0_  (.A1(\V2/V1/A1/A2/M4/s1 ),
    .A2(\V2/V1/A1/A2/c3 ),
    .ZN(\V2/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A1/A2/M4/M2/_1_  (.A(\V2/V1/A1/A2/M4/s1 ),
    .B(\V2/V1/A1/A2/c3 ),
    .Z(\V2/V1/s1 [7]));
 OR2_X1 \V2/V1/A1/A2/M4/_0_  (.A1(\V2/V1/A1/A2/M4/c1 ),
    .A2(\V2/V1/A1/A2/M4/c2 ),
    .ZN(\V2/V1/c1 ));
 AND2_X1 \V2/V1/A2/A1/M1/M1/_0_  (.A1(\V2/V1/s1 [0]),
    .A2(\V2/V1/v1 [4]),
    .ZN(\V2/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M1/M1/_1_  (.A(\V2/V1/s1 [0]),
    .B(\V2/V1/v1 [4]),
    .Z(\V2/V1/A2/A1/M1/s1 ));
 AND2_X1 \V2/V1/A2/A1/M1/M2/_0_  (.A1(\V2/V1/A2/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M1/M2/_1_  (.A(\V2/V1/A2/A1/M1/s1 ),
    .B(net4),
    .Z(v2[4]));
 OR2_X1 \V2/V1/A2/A1/M1/_0_  (.A1(\V2/V1/A2/A1/M1/c1 ),
    .A2(\V2/V1/A2/A1/M1/c2 ),
    .ZN(\V2/V1/A2/A1/c1 ));
 AND2_X1 \V2/V1/A2/A1/M2/M1/_0_  (.A1(\V2/V1/s1 [1]),
    .A2(\V2/V1/v1 [5]),
    .ZN(\V2/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M2/M1/_1_  (.A(\V2/V1/s1 [1]),
    .B(\V2/V1/v1 [5]),
    .Z(\V2/V1/A2/A1/M2/s1 ));
 AND2_X1 \V2/V1/A2/A1/M2/M2/_0_  (.A1(\V2/V1/A2/A1/M2/s1 ),
    .A2(\V2/V1/A2/A1/c1 ),
    .ZN(\V2/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M2/M2/_1_  (.A(\V2/V1/A2/A1/M2/s1 ),
    .B(\V2/V1/A2/A1/c1 ),
    .Z(v2[5]));
 OR2_X1 \V2/V1/A2/A1/M2/_0_  (.A1(\V2/V1/A2/A1/M2/c1 ),
    .A2(\V2/V1/A2/A1/M2/c2 ),
    .ZN(\V2/V1/A2/A1/c2 ));
 AND2_X1 \V2/V1/A2/A1/M3/M1/_0_  (.A1(\V2/V1/s1 [2]),
    .A2(\V2/V1/v1 [6]),
    .ZN(\V2/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M3/M1/_1_  (.A(\V2/V1/s1 [2]),
    .B(\V2/V1/v1 [6]),
    .Z(\V2/V1/A2/A1/M3/s1 ));
 AND2_X1 \V2/V1/A2/A1/M3/M2/_0_  (.A1(\V2/V1/A2/A1/M3/s1 ),
    .A2(\V2/V1/A2/A1/c2 ),
    .ZN(\V2/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M3/M2/_1_  (.A(\V2/V1/A2/A1/M3/s1 ),
    .B(\V2/V1/A2/A1/c2 ),
    .Z(v2[6]));
 OR2_X1 \V2/V1/A2/A1/M3/_0_  (.A1(\V2/V1/A2/A1/M3/c1 ),
    .A2(\V2/V1/A2/A1/M3/c2 ),
    .ZN(\V2/V1/A2/A1/c3 ));
 AND2_X1 \V2/V1/A2/A1/M4/M1/_0_  (.A1(\V2/V1/s1 [3]),
    .A2(\V2/V1/v1 [7]),
    .ZN(\V2/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A2/A1/M4/M1/_1_  (.A(\V2/V1/s1 [3]),
    .B(\V2/V1/v1 [7]),
    .Z(\V2/V1/A2/A1/M4/s1 ));
 AND2_X1 \V2/V1/A2/A1/M4/M2/_0_  (.A1(\V2/V1/A2/A1/M4/s1 ),
    .A2(\V2/V1/A2/A1/c3 ),
    .ZN(\V2/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A2/A1/M4/M2/_1_  (.A(\V2/V1/A2/A1/M4/s1 ),
    .B(\V2/V1/A2/A1/c3 ),
    .Z(v2[7]));
 OR2_X1 \V2/V1/A2/A1/M4/_0_  (.A1(\V2/V1/A2/A1/M4/c1 ),
    .A2(\V2/V1/A2/A1/M4/c2 ),
    .ZN(\V2/V1/A2/c1 ));
 AND2_X1 \V2/V1/A2/A2/M1/M1/_0_  (.A1(\V2/V1/s1 [4]),
    .A2(net4),
    .ZN(\V2/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M1/M1/_1_  (.A(\V2/V1/s1 [4]),
    .B(net4),
    .Z(\V2/V1/A2/A2/M1/s1 ));
 AND2_X1 \V2/V1/A2/A2/M1/M2/_0_  (.A1(\V2/V1/A2/A2/M1/s1 ),
    .A2(\V2/V1/A2/c1 ),
    .ZN(\V2/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M1/M2/_1_  (.A(\V2/V1/A2/A2/M1/s1 ),
    .B(\V2/V1/A2/c1 ),
    .Z(\V2/V1/s2 [4]));
 OR2_X1 \V2/V1/A2/A2/M1/_0_  (.A1(\V2/V1/A2/A2/M1/c1 ),
    .A2(\V2/V1/A2/A2/M1/c2 ),
    .ZN(\V2/V1/A2/A2/c1 ));
 AND2_X1 \V2/V1/A2/A2/M2/M1/_0_  (.A1(\V2/V1/s1 [5]),
    .A2(net4),
    .ZN(\V2/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M2/M1/_1_  (.A(\V2/V1/s1 [5]),
    .B(net4),
    .Z(\V2/V1/A2/A2/M2/s1 ));
 AND2_X1 \V2/V1/A2/A2/M2/M2/_0_  (.A1(\V2/V1/A2/A2/M2/s1 ),
    .A2(\V2/V1/A2/A2/c1 ),
    .ZN(\V2/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M2/M2/_1_  (.A(\V2/V1/A2/A2/M2/s1 ),
    .B(\V2/V1/A2/A2/c1 ),
    .Z(\V2/V1/s2 [5]));
 OR2_X1 \V2/V1/A2/A2/M2/_0_  (.A1(\V2/V1/A2/A2/M2/c1 ),
    .A2(\V2/V1/A2/A2/M2/c2 ),
    .ZN(\V2/V1/A2/A2/c2 ));
 AND2_X1 \V2/V1/A2/A2/M3/M1/_0_  (.A1(\V2/V1/s1 [6]),
    .A2(net4),
    .ZN(\V2/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M3/M1/_1_  (.A(\V2/V1/s1 [6]),
    .B(net4),
    .Z(\V2/V1/A2/A2/M3/s1 ));
 AND2_X1 \V2/V1/A2/A2/M3/M2/_0_  (.A1(\V2/V1/A2/A2/M3/s1 ),
    .A2(\V2/V1/A2/A2/c2 ),
    .ZN(\V2/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M3/M2/_1_  (.A(\V2/V1/A2/A2/M3/s1 ),
    .B(\V2/V1/A2/A2/c2 ),
    .Z(\V2/V1/s2 [6]));
 OR2_X1 \V2/V1/A2/A2/M3/_0_  (.A1(\V2/V1/A2/A2/M3/c1 ),
    .A2(\V2/V1/A2/A2/M3/c2 ),
    .ZN(\V2/V1/A2/A2/c3 ));
 AND2_X1 \V2/V1/A2/A2/M4/M1/_0_  (.A1(\V2/V1/s1 [7]),
    .A2(net4),
    .ZN(\V2/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A2/A2/M4/M1/_1_  (.A(\V2/V1/s1 [7]),
    .B(net4),
    .Z(\V2/V1/A2/A2/M4/s1 ));
 AND2_X1 \V2/V1/A2/A2/M4/M2/_0_  (.A1(\V2/V1/A2/A2/M4/s1 ),
    .A2(\V2/V1/A2/A2/c3 ),
    .ZN(\V2/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A2/A2/M4/M2/_1_  (.A(\V2/V1/A2/A2/M4/s1 ),
    .B(\V2/V1/A2/A2/c3 ),
    .Z(\V2/V1/s2 [7]));
 OR2_X1 \V2/V1/A2/A2/M4/_0_  (.A1(\V2/V1/A2/A2/M4/c1 ),
    .A2(\V2/V1/A2/A2/M4/c2 ),
    .ZN(\V2/V1/c2 ));
 AND2_X1 \V2/V1/A3/A1/M1/M1/_0_  (.A1(\V2/V1/v4 [0]),
    .A2(\V2/V1/s2 [4]),
    .ZN(\V2/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M1/M1/_1_  (.A(\V2/V1/v4 [0]),
    .B(\V2/V1/s2 [4]),
    .Z(\V2/V1/A3/A1/M1/s1 ));
 AND2_X1 \V2/V1/A3/A1/M1/M2/_0_  (.A1(\V2/V1/A3/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V2/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M1/M2/_1_  (.A(\V2/V1/A3/A1/M1/s1 ),
    .B(net6),
    .Z(\V2/v1 [8]));
 OR2_X1 \V2/V1/A3/A1/M1/_0_  (.A1(\V2/V1/A3/A1/M1/c1 ),
    .A2(\V2/V1/A3/A1/M1/c2 ),
    .ZN(\V2/V1/A3/A1/c1 ));
 AND2_X1 \V2/V1/A3/A1/M2/M1/_0_  (.A1(\V2/V1/v4 [1]),
    .A2(\V2/V1/s2 [5]),
    .ZN(\V2/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M2/M1/_1_  (.A(\V2/V1/v4 [1]),
    .B(\V2/V1/s2 [5]),
    .Z(\V2/V1/A3/A1/M2/s1 ));
 AND2_X1 \V2/V1/A3/A1/M2/M2/_0_  (.A1(\V2/V1/A3/A1/M2/s1 ),
    .A2(\V2/V1/A3/A1/c1 ),
    .ZN(\V2/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M2/M2/_1_  (.A(\V2/V1/A3/A1/M2/s1 ),
    .B(\V2/V1/A3/A1/c1 ),
    .Z(\V2/v1 [9]));
 OR2_X1 \V2/V1/A3/A1/M2/_0_  (.A1(\V2/V1/A3/A1/M2/c1 ),
    .A2(\V2/V1/A3/A1/M2/c2 ),
    .ZN(\V2/V1/A3/A1/c2 ));
 AND2_X1 \V2/V1/A3/A1/M3/M1/_0_  (.A1(\V2/V1/v4 [2]),
    .A2(\V2/V1/s2 [6]),
    .ZN(\V2/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M3/M1/_1_  (.A(\V2/V1/v4 [2]),
    .B(\V2/V1/s2 [6]),
    .Z(\V2/V1/A3/A1/M3/s1 ));
 AND2_X1 \V2/V1/A3/A1/M3/M2/_0_  (.A1(\V2/V1/A3/A1/M3/s1 ),
    .A2(\V2/V1/A3/A1/c2 ),
    .ZN(\V2/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M3/M2/_1_  (.A(\V2/V1/A3/A1/M3/s1 ),
    .B(\V2/V1/A3/A1/c2 ),
    .Z(\V2/v1 [10]));
 OR2_X1 \V2/V1/A3/A1/M3/_0_  (.A1(\V2/V1/A3/A1/M3/c1 ),
    .A2(\V2/V1/A3/A1/M3/c2 ),
    .ZN(\V2/V1/A3/A1/c3 ));
 AND2_X1 \V2/V1/A3/A1/M4/M1/_0_  (.A1(\V2/V1/v4 [3]),
    .A2(\V2/V1/s2 [7]),
    .ZN(\V2/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V1/A3/A1/M4/M1/_1_  (.A(\V2/V1/v4 [3]),
    .B(\V2/V1/s2 [7]),
    .Z(\V2/V1/A3/A1/M4/s1 ));
 AND2_X1 \V2/V1/A3/A1/M4/M2/_0_  (.A1(\V2/V1/A3/A1/M4/s1 ),
    .A2(\V2/V1/A3/A1/c3 ),
    .ZN(\V2/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V1/A3/A1/M4/M2/_1_  (.A(\V2/V1/A3/A1/M4/s1 ),
    .B(\V2/V1/A3/A1/c3 ),
    .Z(\V2/v1 [11]));
 OR2_X1 \V2/V1/A3/A1/M4/_0_  (.A1(\V2/V1/A3/A1/M4/c1 ),
    .A2(\V2/V1/A3/A1/M4/c2 ),
    .ZN(\V2/V1/A3/c1 ));
 AND2_X1 \V2/V1/A3/A2/M1/M1/_0_  (.A1(\V2/V1/v4 [4]),
    .A2(\V2/V1/c3 ),
    .ZN(\V2/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M1/M1/_1_  (.A(\V2/V1/v4 [4]),
    .B(\V2/V1/c3 ),
    .Z(\V2/V1/A3/A2/M1/s1 ));
 AND2_X1 \V2/V1/A3/A2/M1/M2/_0_  (.A1(\V2/V1/A3/A2/M1/s1 ),
    .A2(\V2/V1/A3/c1 ),
    .ZN(\V2/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M1/M2/_1_  (.A(\V2/V1/A3/A2/M1/s1 ),
    .B(\V2/V1/A3/c1 ),
    .Z(\V2/v1 [12]));
 OR2_X1 \V2/V1/A3/A2/M1/_0_  (.A1(\V2/V1/A3/A2/M1/c1 ),
    .A2(\V2/V1/A3/A2/M1/c2 ),
    .ZN(\V2/V1/A3/A2/c1 ));
 AND2_X1 \V2/V1/A3/A2/M2/M1/_0_  (.A1(\V2/V1/v4 [5]),
    .A2(net2),
    .ZN(\V2/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M2/M1/_1_  (.A(\V2/V1/v4 [5]),
    .B(net2),
    .Z(\V2/V1/A3/A2/M2/s1 ));
 AND2_X1 \V2/V1/A3/A2/M2/M2/_0_  (.A1(\V2/V1/A3/A2/M2/s1 ),
    .A2(\V2/V1/A3/A2/c1 ),
    .ZN(\V2/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M2/M2/_1_  (.A(\V2/V1/A3/A2/M2/s1 ),
    .B(\V2/V1/A3/A2/c1 ),
    .Z(\V2/v1 [13]));
 OR2_X1 \V2/V1/A3/A2/M2/_0_  (.A1(\V2/V1/A3/A2/M2/c1 ),
    .A2(\V2/V1/A3/A2/M2/c2 ),
    .ZN(\V2/V1/A3/A2/c2 ));
 AND2_X1 \V2/V1/A3/A2/M3/M1/_0_  (.A1(\V2/V1/v4 [6]),
    .A2(net2),
    .ZN(\V2/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M3/M1/_1_  (.A(\V2/V1/v4 [6]),
    .B(net2),
    .Z(\V2/V1/A3/A2/M3/s1 ));
 AND2_X1 \V2/V1/A3/A2/M3/M2/_0_  (.A1(\V2/V1/A3/A2/M3/s1 ),
    .A2(\V2/V1/A3/A2/c2 ),
    .ZN(\V2/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M3/M2/_1_  (.A(\V2/V1/A3/A2/M3/s1 ),
    .B(\V2/V1/A3/A2/c2 ),
    .Z(\V2/v1 [14]));
 OR2_X1 \V2/V1/A3/A2/M3/_0_  (.A1(\V2/V1/A3/A2/M3/c1 ),
    .A2(\V2/V1/A3/A2/M3/c2 ),
    .ZN(\V2/V1/A3/A2/c3 ));
 AND2_X1 \V2/V1/A3/A2/M4/M1/_0_  (.A1(\V2/V1/v4 [7]),
    .A2(net2),
    .ZN(\V2/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V1/A3/A2/M4/M1/_1_  (.A(\V2/V1/v4 [7]),
    .B(net2),
    .Z(\V2/V1/A3/A2/M4/s1 ));
 AND2_X1 \V2/V1/A3/A2/M4/M2/_0_  (.A1(\V2/V1/A3/A2/M4/s1 ),
    .A2(\V2/V1/A3/A2/c3 ),
    .ZN(\V2/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V1/A3/A2/M4/M2/_1_  (.A(\V2/V1/A3/A2/M4/s1 ),
    .B(\V2/V1/A3/A2/c3 ),
    .Z(\V2/v1 [15]));
 OR2_X1 \V2/V1/A3/A2/M4/_0_  (.A1(\V2/V1/A3/A2/M4/c1 ),
    .A2(\V2/V1/A3/A2/M4/c2 ),
    .ZN(\V2/V1/overflow ));
 AND2_X1 \V2/V1/V1/A1/M1/M1/_0_  (.A1(\V2/V1/V1/v2 [0]),
    .A2(\V2/V1/V1/v3 [0]),
    .ZN(\V2/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M1/M1/_1_  (.A(\V2/V1/V1/v2 [0]),
    .B(\V2/V1/V1/v3 [0]),
    .Z(\V2/V1/V1/A1/M1/s1 ));
 AND2_X1 \V2/V1/V1/A1/M1/M2/_0_  (.A1(\V2/V1/V1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M1/M2/_1_  (.A(\V2/V1/V1/A1/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/V1/s1 [0]));
 OR2_X1 \V2/V1/V1/A1/M1/_0_  (.A1(\V2/V1/V1/A1/M1/c1 ),
    .A2(\V2/V1/V1/A1/M1/c2 ),
    .ZN(\V2/V1/V1/A1/c1 ));
 AND2_X1 \V2/V1/V1/A1/M2/M1/_0_  (.A1(\V2/V1/V1/v2 [1]),
    .A2(\V2/V1/V1/v3 [1]),
    .ZN(\V2/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M2/M1/_1_  (.A(\V2/V1/V1/v2 [1]),
    .B(\V2/V1/V1/v3 [1]),
    .Z(\V2/V1/V1/A1/M2/s1 ));
 AND2_X1 \V2/V1/V1/A1/M2/M2/_0_  (.A1(\V2/V1/V1/A1/M2/s1 ),
    .A2(\V2/V1/V1/A1/c1 ),
    .ZN(\V2/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M2/M2/_1_  (.A(\V2/V1/V1/A1/M2/s1 ),
    .B(\V2/V1/V1/A1/c1 ),
    .Z(\V2/V1/V1/s1 [1]));
 OR2_X1 \V2/V1/V1/A1/M2/_0_  (.A1(\V2/V1/V1/A1/M2/c1 ),
    .A2(\V2/V1/V1/A1/M2/c2 ),
    .ZN(\V2/V1/V1/A1/c2 ));
 AND2_X1 \V2/V1/V1/A1/M3/M1/_0_  (.A1(\V2/V1/V1/v2 [2]),
    .A2(\V2/V1/V1/v3 [2]),
    .ZN(\V2/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M3/M1/_1_  (.A(\V2/V1/V1/v2 [2]),
    .B(\V2/V1/V1/v3 [2]),
    .Z(\V2/V1/V1/A1/M3/s1 ));
 AND2_X1 \V2/V1/V1/A1/M3/M2/_0_  (.A1(\V2/V1/V1/A1/M3/s1 ),
    .A2(\V2/V1/V1/A1/c2 ),
    .ZN(\V2/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M3/M2/_1_  (.A(\V2/V1/V1/A1/M3/s1 ),
    .B(\V2/V1/V1/A1/c2 ),
    .Z(\V2/V1/V1/s1 [2]));
 OR2_X1 \V2/V1/V1/A1/M3/_0_  (.A1(\V2/V1/V1/A1/M3/c1 ),
    .A2(\V2/V1/V1/A1/M3/c2 ),
    .ZN(\V2/V1/V1/A1/c3 ));
 AND2_X1 \V2/V1/V1/A1/M4/M1/_0_  (.A1(\V2/V1/V1/v2 [3]),
    .A2(\V2/V1/V1/v3 [3]),
    .ZN(\V2/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A1/M4/M1/_1_  (.A(\V2/V1/V1/v2 [3]),
    .B(\V2/V1/V1/v3 [3]),
    .Z(\V2/V1/V1/A1/M4/s1 ));
 AND2_X1 \V2/V1/V1/A1/M4/M2/_0_  (.A1(\V2/V1/V1/A1/M4/s1 ),
    .A2(\V2/V1/V1/A1/c3 ),
    .ZN(\V2/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A1/M4/M2/_1_  (.A(\V2/V1/V1/A1/M4/s1 ),
    .B(\V2/V1/V1/A1/c3 ),
    .Z(\V2/V1/V1/s1 [3]));
 OR2_X1 \V2/V1/V1/A1/M4/_0_  (.A1(\V2/V1/V1/A1/M4/c1 ),
    .A2(\V2/V1/V1/A1/M4/c2 ),
    .ZN(\V2/V1/V1/c1 ));
 AND2_X1 \V2/V1/V1/A2/M1/M1/_0_  (.A1(\V2/V1/V1/s1 [0]),
    .A2(\V2/V1/V1/v1 [2]),
    .ZN(\V2/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M1/M1/_1_  (.A(\V2/V1/V1/s1 [0]),
    .B(\V2/V1/V1/v1 [2]),
    .Z(\V2/V1/V1/A2/M1/s1 ));
 AND2_X1 \V2/V1/V1/A2/M1/M2/_0_  (.A1(\V2/V1/V1/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M1/M2/_1_  (.A(\V2/V1/V1/A2/M1/s1 ),
    .B(net4),
    .Z(v2[2]));
 OR2_X1 \V2/V1/V1/A2/M1/_0_  (.A1(\V2/V1/V1/A2/M1/c1 ),
    .A2(\V2/V1/V1/A2/M1/c2 ),
    .ZN(\V2/V1/V1/A2/c1 ));
 AND2_X1 \V2/V1/V1/A2/M2/M1/_0_  (.A1(\V2/V1/V1/s1 [1]),
    .A2(\V2/V1/V1/v1 [3]),
    .ZN(\V2/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M2/M1/_1_  (.A(\V2/V1/V1/s1 [1]),
    .B(\V2/V1/V1/v1 [3]),
    .Z(\V2/V1/V1/A2/M2/s1 ));
 AND2_X1 \V2/V1/V1/A2/M2/M2/_0_  (.A1(\V2/V1/V1/A2/M2/s1 ),
    .A2(\V2/V1/V1/A2/c1 ),
    .ZN(\V2/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M2/M2/_1_  (.A(\V2/V1/V1/A2/M2/s1 ),
    .B(\V2/V1/V1/A2/c1 ),
    .Z(v2[3]));
 OR2_X1 \V2/V1/V1/A2/M2/_0_  (.A1(\V2/V1/V1/A2/M2/c1 ),
    .A2(\V2/V1/V1/A2/M2/c2 ),
    .ZN(\V2/V1/V1/A2/c2 ));
 AND2_X1 \V2/V1/V1/A2/M3/M1/_0_  (.A1(\V2/V1/V1/s1 [2]),
    .A2(net4),
    .ZN(\V2/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M3/M1/_1_  (.A(\V2/V1/V1/s1 [2]),
    .B(net4),
    .Z(\V2/V1/V1/A2/M3/s1 ));
 AND2_X1 \V2/V1/V1/A2/M3/M2/_0_  (.A1(\V2/V1/V1/A2/M3/s1 ),
    .A2(\V2/V1/V1/A2/c2 ),
    .ZN(\V2/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M3/M2/_1_  (.A(\V2/V1/V1/A2/M3/s1 ),
    .B(\V2/V1/V1/A2/c2 ),
    .Z(\V2/V1/V1/s2 [2]));
 OR2_X1 \V2/V1/V1/A2/M3/_0_  (.A1(\V2/V1/V1/A2/M3/c1 ),
    .A2(\V2/V1/V1/A2/M3/c2 ),
    .ZN(\V2/V1/V1/A2/c3 ));
 AND2_X1 \V2/V1/V1/A2/M4/M1/_0_  (.A1(\V2/V1/V1/s1 [3]),
    .A2(net4),
    .ZN(\V2/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A2/M4/M1/_1_  (.A(\V2/V1/V1/s1 [3]),
    .B(net4),
    .Z(\V2/V1/V1/A2/M4/s1 ));
 AND2_X1 \V2/V1/V1/A2/M4/M2/_0_  (.A1(\V2/V1/V1/A2/M4/s1 ),
    .A2(\V2/V1/V1/A2/c3 ),
    .ZN(\V2/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A2/M4/M2/_1_  (.A(\V2/V1/V1/A2/M4/s1 ),
    .B(\V2/V1/V1/A2/c3 ),
    .Z(\V2/V1/V1/s2 [3]));
 OR2_X1 \V2/V1/V1/A2/M4/_0_  (.A1(\V2/V1/V1/A2/M4/c1 ),
    .A2(\V2/V1/V1/A2/M4/c2 ),
    .ZN(\V2/V1/V1/c2 ));
 AND2_X1 \V2/V1/V1/A3/M1/M1/_0_  (.A1(\V2/V1/V1/v4 [0]),
    .A2(\V2/V1/V1/s2 [2]),
    .ZN(\V2/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M1/M1/_1_  (.A(\V2/V1/V1/v4 [0]),
    .B(\V2/V1/V1/s2 [2]),
    .Z(\V2/V1/V1/A3/M1/s1 ));
 AND2_X1 \V2/V1/V1/A3/M1/M2/_0_  (.A1(\V2/V1/V1/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M1/M2/_1_  (.A(\V2/V1/V1/A3/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/v1 [4]));
 OR2_X1 \V2/V1/V1/A3/M1/_0_  (.A1(\V2/V1/V1/A3/M1/c1 ),
    .A2(\V2/V1/V1/A3/M1/c2 ),
    .ZN(\V2/V1/V1/A3/c1 ));
 AND2_X1 \V2/V1/V1/A3/M2/M1/_0_  (.A1(\V2/V1/V1/v4 [1]),
    .A2(\V2/V1/V1/s2 [3]),
    .ZN(\V2/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M2/M1/_1_  (.A(\V2/V1/V1/v4 [1]),
    .B(\V2/V1/V1/s2 [3]),
    .Z(\V2/V1/V1/A3/M2/s1 ));
 AND2_X1 \V2/V1/V1/A3/M2/M2/_0_  (.A1(\V2/V1/V1/A3/M2/s1 ),
    .A2(\V2/V1/V1/A3/c1 ),
    .ZN(\V2/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M2/M2/_1_  (.A(\V2/V1/V1/A3/M2/s1 ),
    .B(\V2/V1/V1/A3/c1 ),
    .Z(\V2/V1/v1 [5]));
 OR2_X1 \V2/V1/V1/A3/M2/_0_  (.A1(\V2/V1/V1/A3/M2/c1 ),
    .A2(\V2/V1/V1/A3/M2/c2 ),
    .ZN(\V2/V1/V1/A3/c2 ));
 AND2_X1 \V2/V1/V1/A3/M3/M1/_0_  (.A1(\V2/V1/V1/v4 [2]),
    .A2(\V2/V1/V1/c3 ),
    .ZN(\V2/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M3/M1/_1_  (.A(\V2/V1/V1/v4 [2]),
    .B(\V2/V1/V1/c3 ),
    .Z(\V2/V1/V1/A3/M3/s1 ));
 AND2_X1 \V2/V1/V1/A3/M3/M2/_0_  (.A1(\V2/V1/V1/A3/M3/s1 ),
    .A2(\V2/V1/V1/A3/c2 ),
    .ZN(\V2/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M3/M2/_1_  (.A(\V2/V1/V1/A3/M3/s1 ),
    .B(\V2/V1/V1/A3/c2 ),
    .Z(\V2/V1/v1 [6]));
 OR2_X1 \V2/V1/V1/A3/M3/_0_  (.A1(\V2/V1/V1/A3/M3/c1 ),
    .A2(\V2/V1/V1/A3/M3/c2 ),
    .ZN(\V2/V1/V1/A3/c3 ));
 AND2_X1 \V2/V1/V1/A3/M4/M1/_0_  (.A1(\V2/V1/V1/v4 [3]),
    .A2(net4),
    .ZN(\V2/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V1/A3/M4/M1/_1_  (.A(\V2/V1/V1/v4 [3]),
    .B(net4),
    .Z(\V2/V1/V1/A3/M4/s1 ));
 AND2_X1 \V2/V1/V1/A3/M4/M2/_0_  (.A1(\V2/V1/V1/A3/M4/s1 ),
    .A2(\V2/V1/V1/A3/c3 ),
    .ZN(\V2/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V1/A3/M4/M2/_1_  (.A(\V2/V1/V1/A3/M4/s1 ),
    .B(\V2/V1/V1/A3/c3 ),
    .Z(\V2/V1/v1 [7]));
 OR2_X1 \V2/V1/V1/A3/M4/_0_  (.A1(\V2/V1/V1/A3/M4/c1 ),
    .A2(\V2/V1/V1/A3/M4/c2 ),
    .ZN(\V2/V1/V1/overflow ));
 AND2_X1 \V2/V1/V1/V1/HA1/_0_  (.A1(\V2/V1/V1/V1/w2 ),
    .A2(\V2/V1/V1/V1/w1 ),
    .ZN(\V2/V1/V1/V1/w4 ));
 XOR2_X2 \V2/V1/V1/V1/HA1/_1_  (.A(\V2/V1/V1/V1/w2 ),
    .B(\V2/V1/V1/V1/w1 ),
    .Z(v2[1]));
 AND2_X1 \V2/V1/V1/V1/HA2/_0_  (.A1(\V2/V1/V1/V1/w4 ),
    .A2(\V2/V1/V1/V1/w3 ),
    .ZN(\V2/V1/V1/v1 [3]));
 XOR2_X2 \V2/V1/V1/V1/HA2/_1_  (.A(\V2/V1/V1/V1/w4 ),
    .B(\V2/V1/V1/V1/w3 ),
    .Z(\V2/V1/V1/v1 [2]));
 AND2_X1 \V2/V1/V1/V1/_0_  (.A1(net41),
    .A2(B[0]),
    .ZN(v2[0]));
 AND2_X1 \V2/V1/V1/V1/_1_  (.A1(net41),
    .A2(B[1]),
    .ZN(\V2/V1/V1/V1/w1 ));
 AND2_X1 \V2/V1/V1/V1/_2_  (.A1(B[0]),
    .A2(net40),
    .ZN(\V2/V1/V1/V1/w2 ));
 AND2_X1 \V2/V1/V1/V1/_3_  (.A1(B[1]),
    .A2(net40),
    .ZN(\V2/V1/V1/V1/w3 ));
 AND2_X1 \V2/V1/V1/V2/HA1/_0_  (.A1(\V2/V1/V1/V2/w2 ),
    .A2(\V2/V1/V1/V2/w1 ),
    .ZN(\V2/V1/V1/V2/w4 ));
 XOR2_X2 \V2/V1/V1/V2/HA1/_1_  (.A(\V2/V1/V1/V2/w2 ),
    .B(\V2/V1/V1/V2/w1 ),
    .Z(\V2/V1/V1/v2 [1]));
 AND2_X1 \V2/V1/V1/V2/HA2/_0_  (.A1(\V2/V1/V1/V2/w4 ),
    .A2(\V2/V1/V1/V2/w3 ),
    .ZN(\V2/V1/V1/v2 [3]));
 XOR2_X2 \V2/V1/V1/V2/HA2/_1_  (.A(\V2/V1/V1/V2/w4 ),
    .B(\V2/V1/V1/V2/w3 ),
    .Z(\V2/V1/V1/v2 [2]));
 AND2_X1 \V2/V1/V1/V2/_0_  (.A1(net39),
    .A2(B[0]),
    .ZN(\V2/V1/V1/v2 [0]));
 AND2_X1 \V2/V1/V1/V2/_1_  (.A1(A[18]),
    .A2(B[1]),
    .ZN(\V2/V1/V1/V2/w1 ));
 AND2_X1 \V2/V1/V1/V2/_2_  (.A1(B[0]),
    .A2(net38),
    .ZN(\V2/V1/V1/V2/w2 ));
 AND2_X1 \V2/V1/V1/V2/_3_  (.A1(B[1]),
    .A2(net38),
    .ZN(\V2/V1/V1/V2/w3 ));
 AND2_X1 \V2/V1/V1/V3/HA1/_0_  (.A1(\V2/V1/V1/V3/w2 ),
    .A2(\V2/V1/V1/V3/w1 ),
    .ZN(\V2/V1/V1/V3/w4 ));
 XOR2_X2 \V2/V1/V1/V3/HA1/_1_  (.A(\V2/V1/V1/V3/w2 ),
    .B(\V2/V1/V1/V3/w1 ),
    .Z(\V2/V1/V1/v3 [1]));
 AND2_X1 \V2/V1/V1/V3/HA2/_0_  (.A1(\V2/V1/V1/V3/w4 ),
    .A2(\V2/V1/V1/V3/w3 ),
    .ZN(\V2/V1/V1/v3 [3]));
 XOR2_X2 \V2/V1/V1/V3/HA2/_1_  (.A(\V2/V1/V1/V3/w4 ),
    .B(\V2/V1/V1/V3/w3 ),
    .Z(\V2/V1/V1/v3 [2]));
 AND2_X1 \V2/V1/V1/V3/_0_  (.A1(net41),
    .A2(B[2]),
    .ZN(\V2/V1/V1/v3 [0]));
 AND2_X1 \V2/V1/V1/V3/_1_  (.A1(net41),
    .A2(B[3]),
    .ZN(\V2/V1/V1/V3/w1 ));
 AND2_X1 \V2/V1/V1/V3/_2_  (.A1(B[2]),
    .A2(net40),
    .ZN(\V2/V1/V1/V3/w2 ));
 AND2_X1 \V2/V1/V1/V3/_3_  (.A1(B[3]),
    .A2(net40),
    .ZN(\V2/V1/V1/V3/w3 ));
 AND2_X1 \V2/V1/V1/V4/HA1/_0_  (.A1(\V2/V1/V1/V4/w2 ),
    .A2(\V2/V1/V1/V4/w1 ),
    .ZN(\V2/V1/V1/V4/w4 ));
 XOR2_X2 \V2/V1/V1/V4/HA1/_1_  (.A(\V2/V1/V1/V4/w2 ),
    .B(\V2/V1/V1/V4/w1 ),
    .Z(\V2/V1/V1/v4 [1]));
 AND2_X1 \V2/V1/V1/V4/HA2/_0_  (.A1(\V2/V1/V1/V4/w4 ),
    .A2(\V2/V1/V1/V4/w3 ),
    .ZN(\V2/V1/V1/v4 [3]));
 XOR2_X2 \V2/V1/V1/V4/HA2/_1_  (.A(\V2/V1/V1/V4/w4 ),
    .B(\V2/V1/V1/V4/w3 ),
    .Z(\V2/V1/V1/v4 [2]));
 AND2_X1 \V2/V1/V1/V4/_0_  (.A1(net39),
    .A2(B[2]),
    .ZN(\V2/V1/V1/v4 [0]));
 AND2_X1 \V2/V1/V1/V4/_1_  (.A1(net39),
    .A2(B[3]),
    .ZN(\V2/V1/V1/V4/w1 ));
 AND2_X1 \V2/V1/V1/V4/_2_  (.A1(B[2]),
    .A2(net38),
    .ZN(\V2/V1/V1/V4/w2 ));
 AND2_X1 \V2/V1/V1/V4/_3_  (.A1(B[3]),
    .A2(net38),
    .ZN(\V2/V1/V1/V4/w3 ));
 OR2_X1 \V2/V1/V1/_0_  (.A1(\V2/V1/V1/c1 ),
    .A2(\V2/V1/V1/c2 ),
    .ZN(\V2/V1/V1/c3 ));
 AND2_X1 \V2/V1/V2/A1/M1/M1/_0_  (.A1(\V2/V1/V2/v2 [0]),
    .A2(\V2/V1/V2/v3 [0]),
    .ZN(\V2/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M1/M1/_1_  (.A(\V2/V1/V2/v2 [0]),
    .B(\V2/V1/V2/v3 [0]),
    .Z(\V2/V1/V2/A1/M1/s1 ));
 AND2_X1 \V2/V1/V2/A1/M1/M2/_0_  (.A1(\V2/V1/V2/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M1/M2/_1_  (.A(\V2/V1/V2/A1/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/V2/s1 [0]));
 OR2_X1 \V2/V1/V2/A1/M1/_0_  (.A1(\V2/V1/V2/A1/M1/c1 ),
    .A2(\V2/V1/V2/A1/M1/c2 ),
    .ZN(\V2/V1/V2/A1/c1 ));
 AND2_X1 \V2/V1/V2/A1/M2/M1/_0_  (.A1(\V2/V1/V2/v2 [1]),
    .A2(\V2/V1/V2/v3 [1]),
    .ZN(\V2/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M2/M1/_1_  (.A(\V2/V1/V2/v2 [1]),
    .B(\V2/V1/V2/v3 [1]),
    .Z(\V2/V1/V2/A1/M2/s1 ));
 AND2_X1 \V2/V1/V2/A1/M2/M2/_0_  (.A1(\V2/V1/V2/A1/M2/s1 ),
    .A2(\V2/V1/V2/A1/c1 ),
    .ZN(\V2/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M2/M2/_1_  (.A(\V2/V1/V2/A1/M2/s1 ),
    .B(\V2/V1/V2/A1/c1 ),
    .Z(\V2/V1/V2/s1 [1]));
 OR2_X1 \V2/V1/V2/A1/M2/_0_  (.A1(\V2/V1/V2/A1/M2/c1 ),
    .A2(\V2/V1/V2/A1/M2/c2 ),
    .ZN(\V2/V1/V2/A1/c2 ));
 AND2_X1 \V2/V1/V2/A1/M3/M1/_0_  (.A1(\V2/V1/V2/v2 [2]),
    .A2(\V2/V1/V2/v3 [2]),
    .ZN(\V2/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M3/M1/_1_  (.A(\V2/V1/V2/v2 [2]),
    .B(\V2/V1/V2/v3 [2]),
    .Z(\V2/V1/V2/A1/M3/s1 ));
 AND2_X1 \V2/V1/V2/A1/M3/M2/_0_  (.A1(\V2/V1/V2/A1/M3/s1 ),
    .A2(\V2/V1/V2/A1/c2 ),
    .ZN(\V2/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M3/M2/_1_  (.A(\V2/V1/V2/A1/M3/s1 ),
    .B(\V2/V1/V2/A1/c2 ),
    .Z(\V2/V1/V2/s1 [2]));
 OR2_X1 \V2/V1/V2/A1/M3/_0_  (.A1(\V2/V1/V2/A1/M3/c1 ),
    .A2(\V2/V1/V2/A1/M3/c2 ),
    .ZN(\V2/V1/V2/A1/c3 ));
 AND2_X1 \V2/V1/V2/A1/M4/M1/_0_  (.A1(\V2/V1/V2/v2 [3]),
    .A2(\V2/V1/V2/v3 [3]),
    .ZN(\V2/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A1/M4/M1/_1_  (.A(\V2/V1/V2/v2 [3]),
    .B(\V2/V1/V2/v3 [3]),
    .Z(\V2/V1/V2/A1/M4/s1 ));
 AND2_X1 \V2/V1/V2/A1/M4/M2/_0_  (.A1(\V2/V1/V2/A1/M4/s1 ),
    .A2(\V2/V1/V2/A1/c3 ),
    .ZN(\V2/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A1/M4/M2/_1_  (.A(\V2/V1/V2/A1/M4/s1 ),
    .B(\V2/V1/V2/A1/c3 ),
    .Z(\V2/V1/V2/s1 [3]));
 OR2_X1 \V2/V1/V2/A1/M4/_0_  (.A1(\V2/V1/V2/A1/M4/c1 ),
    .A2(\V2/V1/V2/A1/M4/c2 ),
    .ZN(\V2/V1/V2/c1 ));
 AND2_X1 \V2/V1/V2/A2/M1/M1/_0_  (.A1(\V2/V1/V2/s1 [0]),
    .A2(\V2/V1/V2/v1 [2]),
    .ZN(\V2/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M1/M1/_1_  (.A(\V2/V1/V2/s1 [0]),
    .B(\V2/V1/V2/v1 [2]),
    .Z(\V2/V1/V2/A2/M1/s1 ));
 AND2_X1 \V2/V1/V2/A2/M1/M2/_0_  (.A1(\V2/V1/V2/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M1/M2/_1_  (.A(\V2/V1/V2/A2/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/v2 [2]));
 OR2_X1 \V2/V1/V2/A2/M1/_0_  (.A1(\V2/V1/V2/A2/M1/c1 ),
    .A2(\V2/V1/V2/A2/M1/c2 ),
    .ZN(\V2/V1/V2/A2/c1 ));
 AND2_X1 \V2/V1/V2/A2/M2/M1/_0_  (.A1(\V2/V1/V2/s1 [1]),
    .A2(\V2/V1/V2/v1 [3]),
    .ZN(\V2/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M2/M1/_1_  (.A(\V2/V1/V2/s1 [1]),
    .B(\V2/V1/V2/v1 [3]),
    .Z(\V2/V1/V2/A2/M2/s1 ));
 AND2_X1 \V2/V1/V2/A2/M2/M2/_0_  (.A1(\V2/V1/V2/A2/M2/s1 ),
    .A2(\V2/V1/V2/A2/c1 ),
    .ZN(\V2/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M2/M2/_1_  (.A(\V2/V1/V2/A2/M2/s1 ),
    .B(\V2/V1/V2/A2/c1 ),
    .Z(\V2/V1/v2 [3]));
 OR2_X1 \V2/V1/V2/A2/M2/_0_  (.A1(\V2/V1/V2/A2/M2/c1 ),
    .A2(\V2/V1/V2/A2/M2/c2 ),
    .ZN(\V2/V1/V2/A2/c2 ));
 AND2_X1 \V2/V1/V2/A2/M3/M1/_0_  (.A1(\V2/V1/V2/s1 [2]),
    .A2(net4),
    .ZN(\V2/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M3/M1/_1_  (.A(\V2/V1/V2/s1 [2]),
    .B(net4),
    .Z(\V2/V1/V2/A2/M3/s1 ));
 AND2_X1 \V2/V1/V2/A2/M3/M2/_0_  (.A1(\V2/V1/V2/A2/M3/s1 ),
    .A2(\V2/V1/V2/A2/c2 ),
    .ZN(\V2/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M3/M2/_1_  (.A(\V2/V1/V2/A2/M3/s1 ),
    .B(\V2/V1/V2/A2/c2 ),
    .Z(\V2/V1/V2/s2 [2]));
 OR2_X1 \V2/V1/V2/A2/M3/_0_  (.A1(\V2/V1/V2/A2/M3/c1 ),
    .A2(\V2/V1/V2/A2/M3/c2 ),
    .ZN(\V2/V1/V2/A2/c3 ));
 AND2_X1 \V2/V1/V2/A2/M4/M1/_0_  (.A1(\V2/V1/V2/s1 [3]),
    .A2(net4),
    .ZN(\V2/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A2/M4/M1/_1_  (.A(\V2/V1/V2/s1 [3]),
    .B(net4),
    .Z(\V2/V1/V2/A2/M4/s1 ));
 AND2_X1 \V2/V1/V2/A2/M4/M2/_0_  (.A1(\V2/V1/V2/A2/M4/s1 ),
    .A2(\V2/V1/V2/A2/c3 ),
    .ZN(\V2/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A2/M4/M2/_1_  (.A(\V2/V1/V2/A2/M4/s1 ),
    .B(\V2/V1/V2/A2/c3 ),
    .Z(\V2/V1/V2/s2 [3]));
 OR2_X1 \V2/V1/V2/A2/M4/_0_  (.A1(\V2/V1/V2/A2/M4/c1 ),
    .A2(\V2/V1/V2/A2/M4/c2 ),
    .ZN(\V2/V1/V2/c2 ));
 AND2_X1 \V2/V1/V2/A3/M1/M1/_0_  (.A1(\V2/V1/V2/v4 [0]),
    .A2(\V2/V1/V2/s2 [2]),
    .ZN(\V2/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M1/M1/_1_  (.A(\V2/V1/V2/v4 [0]),
    .B(\V2/V1/V2/s2 [2]),
    .Z(\V2/V1/V2/A3/M1/s1 ));
 AND2_X1 \V2/V1/V2/A3/M1/M2/_0_  (.A1(\V2/V1/V2/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M1/M2/_1_  (.A(\V2/V1/V2/A3/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/v2 [4]));
 OR2_X1 \V2/V1/V2/A3/M1/_0_  (.A1(\V2/V1/V2/A3/M1/c1 ),
    .A2(\V2/V1/V2/A3/M1/c2 ),
    .ZN(\V2/V1/V2/A3/c1 ));
 AND2_X1 \V2/V1/V2/A3/M2/M1/_0_  (.A1(\V2/V1/V2/v4 [1]),
    .A2(\V2/V1/V2/s2 [3]),
    .ZN(\V2/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M2/M1/_1_  (.A(\V2/V1/V2/v4 [1]),
    .B(\V2/V1/V2/s2 [3]),
    .Z(\V2/V1/V2/A3/M2/s1 ));
 AND2_X1 \V2/V1/V2/A3/M2/M2/_0_  (.A1(\V2/V1/V2/A3/M2/s1 ),
    .A2(\V2/V1/V2/A3/c1 ),
    .ZN(\V2/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M2/M2/_1_  (.A(\V2/V1/V2/A3/M2/s1 ),
    .B(\V2/V1/V2/A3/c1 ),
    .Z(\V2/V1/v2 [5]));
 OR2_X1 \V2/V1/V2/A3/M2/_0_  (.A1(\V2/V1/V2/A3/M2/c1 ),
    .A2(\V2/V1/V2/A3/M2/c2 ),
    .ZN(\V2/V1/V2/A3/c2 ));
 AND2_X1 \V2/V1/V2/A3/M3/M1/_0_  (.A1(\V2/V1/V2/v4 [2]),
    .A2(\V2/V1/V2/c3 ),
    .ZN(\V2/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M3/M1/_1_  (.A(\V2/V1/V2/v4 [2]),
    .B(\V2/V1/V2/c3 ),
    .Z(\V2/V1/V2/A3/M3/s1 ));
 AND2_X1 \V2/V1/V2/A3/M3/M2/_0_  (.A1(\V2/V1/V2/A3/M3/s1 ),
    .A2(\V2/V1/V2/A3/c2 ),
    .ZN(\V2/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M3/M2/_1_  (.A(\V2/V1/V2/A3/M3/s1 ),
    .B(\V2/V1/V2/A3/c2 ),
    .Z(\V2/V1/v2 [6]));
 OR2_X1 \V2/V1/V2/A3/M3/_0_  (.A1(\V2/V1/V2/A3/M3/c1 ),
    .A2(\V2/V1/V2/A3/M3/c2 ),
    .ZN(\V2/V1/V2/A3/c3 ));
 AND2_X1 \V2/V1/V2/A3/M4/M1/_0_  (.A1(\V2/V1/V2/v4 [3]),
    .A2(net4),
    .ZN(\V2/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V2/A3/M4/M1/_1_  (.A(\V2/V1/V2/v4 [3]),
    .B(net4),
    .Z(\V2/V1/V2/A3/M4/s1 ));
 AND2_X1 \V2/V1/V2/A3/M4/M2/_0_  (.A1(\V2/V1/V2/A3/M4/s1 ),
    .A2(\V2/V1/V2/A3/c3 ),
    .ZN(\V2/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V2/A3/M4/M2/_1_  (.A(\V2/V1/V2/A3/M4/s1 ),
    .B(\V2/V1/V2/A3/c3 ),
    .Z(\V2/V1/v2 [7]));
 OR2_X1 \V2/V1/V2/A3/M4/_0_  (.A1(\V2/V1/V2/A3/M4/c1 ),
    .A2(\V2/V1/V2/A3/M4/c2 ),
    .ZN(\V2/V1/V2/overflow ));
 AND2_X1 \V2/V1/V2/V1/HA1/_0_  (.A1(\V2/V1/V2/V1/w2 ),
    .A2(\V2/V1/V2/V1/w1 ),
    .ZN(\V2/V1/V2/V1/w4 ));
 XOR2_X2 \V2/V1/V2/V1/HA1/_1_  (.A(\V2/V1/V2/V1/w2 ),
    .B(\V2/V1/V2/V1/w1 ),
    .Z(\V2/V1/v2 [1]));
 AND2_X1 \V2/V1/V2/V1/HA2/_0_  (.A1(\V2/V1/V2/V1/w4 ),
    .A2(\V2/V1/V2/V1/w3 ),
    .ZN(\V2/V1/V2/v1 [3]));
 XOR2_X2 \V2/V1/V2/V1/HA2/_1_  (.A(\V2/V1/V2/V1/w4 ),
    .B(\V2/V1/V2/V1/w3 ),
    .Z(\V2/V1/V2/v1 [2]));
 AND2_X1 \V2/V1/V2/V1/_0_  (.A1(A[20]),
    .A2(B[0]),
    .ZN(\V2/V1/v2 [0]));
 AND2_X1 \V2/V1/V2/V1/_1_  (.A1(A[20]),
    .A2(B[1]),
    .ZN(\V2/V1/V2/V1/w1 ));
 AND2_X1 \V2/V1/V2/V1/_2_  (.A1(B[0]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V1/w2 ));
 AND2_X1 \V2/V1/V2/V1/_3_  (.A1(B[1]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V1/w3 ));
 AND2_X1 \V2/V1/V2/V2/HA1/_0_  (.A1(\V2/V1/V2/V2/w2 ),
    .A2(\V2/V1/V2/V2/w1 ),
    .ZN(\V2/V1/V2/V2/w4 ));
 XOR2_X2 \V2/V1/V2/V2/HA1/_1_  (.A(\V2/V1/V2/V2/w2 ),
    .B(\V2/V1/V2/V2/w1 ),
    .Z(\V2/V1/V2/v2 [1]));
 AND2_X1 \V2/V1/V2/V2/HA2/_0_  (.A1(\V2/V1/V2/V2/w4 ),
    .A2(\V2/V1/V2/V2/w3 ),
    .ZN(\V2/V1/V2/v2 [3]));
 XOR2_X2 \V2/V1/V2/V2/HA2/_1_  (.A(\V2/V1/V2/V2/w4 ),
    .B(\V2/V1/V2/V2/w3 ),
    .Z(\V2/V1/V2/v2 [2]));
 AND2_X1 \V2/V1/V2/V2/_0_  (.A1(net35),
    .A2(B[0]),
    .ZN(\V2/V1/V2/v2 [0]));
 AND2_X1 \V2/V1/V2/V2/_1_  (.A1(net35),
    .A2(B[1]),
    .ZN(\V2/V1/V2/V2/w1 ));
 AND2_X1 \V2/V1/V2/V2/_2_  (.A1(B[0]),
    .A2(net34),
    .ZN(\V2/V1/V2/V2/w2 ));
 AND2_X1 \V2/V1/V2/V2/_3_  (.A1(B[1]),
    .A2(net34),
    .ZN(\V2/V1/V2/V2/w3 ));
 AND2_X1 \V2/V1/V2/V3/HA1/_0_  (.A1(\V2/V1/V2/V3/w2 ),
    .A2(\V2/V1/V2/V3/w1 ),
    .ZN(\V2/V1/V2/V3/w4 ));
 XOR2_X2 \V2/V1/V2/V3/HA1/_1_  (.A(\V2/V1/V2/V3/w2 ),
    .B(\V2/V1/V2/V3/w1 ),
    .Z(\V2/V1/V2/v3 [1]));
 AND2_X1 \V2/V1/V2/V3/HA2/_0_  (.A1(\V2/V1/V2/V3/w4 ),
    .A2(\V2/V1/V2/V3/w3 ),
    .ZN(\V2/V1/V2/v3 [3]));
 XOR2_X2 \V2/V1/V2/V3/HA2/_1_  (.A(\V2/V1/V2/V3/w4 ),
    .B(\V2/V1/V2/V3/w3 ),
    .Z(\V2/V1/V2/v3 [2]));
 AND2_X1 \V2/V1/V2/V3/_0_  (.A1(A[20]),
    .A2(B[2]),
    .ZN(\V2/V1/V2/v3 [0]));
 AND2_X1 \V2/V1/V2/V3/_1_  (.A1(A[20]),
    .A2(B[3]),
    .ZN(\V2/V1/V2/V3/w1 ));
 AND2_X1 \V2/V1/V2/V3/_2_  (.A1(B[2]),
    .A2(A[21]),
    .ZN(\V2/V1/V2/V3/w2 ));
 AND2_X1 \V2/V1/V2/V3/_3_  (.A1(B[3]),
    .A2(net36),
    .ZN(\V2/V1/V2/V3/w3 ));
 AND2_X1 \V2/V1/V2/V4/HA1/_0_  (.A1(\V2/V1/V2/V4/w2 ),
    .A2(\V2/V1/V2/V4/w1 ),
    .ZN(\V2/V1/V2/V4/w4 ));
 XOR2_X2 \V2/V1/V2/V4/HA1/_1_  (.A(\V2/V1/V2/V4/w2 ),
    .B(\V2/V1/V2/V4/w1 ),
    .Z(\V2/V1/V2/v4 [1]));
 AND2_X1 \V2/V1/V2/V4/HA2/_0_  (.A1(\V2/V1/V2/V4/w4 ),
    .A2(\V2/V1/V2/V4/w3 ),
    .ZN(\V2/V1/V2/v4 [3]));
 XOR2_X2 \V2/V1/V2/V4/HA2/_1_  (.A(\V2/V1/V2/V4/w4 ),
    .B(\V2/V1/V2/V4/w3 ),
    .Z(\V2/V1/V2/v4 [2]));
 AND2_X1 \V2/V1/V2/V4/_0_  (.A1(net35),
    .A2(B[2]),
    .ZN(\V2/V1/V2/v4 [0]));
 AND2_X1 \V2/V1/V2/V4/_1_  (.A1(net35),
    .A2(B[3]),
    .ZN(\V2/V1/V2/V4/w1 ));
 AND2_X1 \V2/V1/V2/V4/_2_  (.A1(B[2]),
    .A2(net34),
    .ZN(\V2/V1/V2/V4/w2 ));
 AND2_X1 \V2/V1/V2/V4/_3_  (.A1(B[3]),
    .A2(net34),
    .ZN(\V2/V1/V2/V4/w3 ));
 OR2_X1 \V2/V1/V2/_0_  (.A1(\V2/V1/V2/c1 ),
    .A2(\V2/V1/V2/c2 ),
    .ZN(\V2/V1/V2/c3 ));
 AND2_X1 \V2/V1/V3/A1/M1/M1/_0_  (.A1(\V2/V1/V3/v2 [0]),
    .A2(\V2/V1/V3/v3 [0]),
    .ZN(\V2/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M1/M1/_1_  (.A(\V2/V1/V3/v2 [0]),
    .B(\V2/V1/V3/v3 [0]),
    .Z(\V2/V1/V3/A1/M1/s1 ));
 AND2_X1 \V2/V1/V3/A1/M1/M2/_0_  (.A1(\V2/V1/V3/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M1/M2/_1_  (.A(\V2/V1/V3/A1/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/V3/s1 [0]));
 OR2_X1 \V2/V1/V3/A1/M1/_0_  (.A1(\V2/V1/V3/A1/M1/c1 ),
    .A2(\V2/V1/V3/A1/M1/c2 ),
    .ZN(\V2/V1/V3/A1/c1 ));
 AND2_X1 \V2/V1/V3/A1/M2/M1/_0_  (.A1(\V2/V1/V3/v2 [1]),
    .A2(\V2/V1/V3/v3 [1]),
    .ZN(\V2/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M2/M1/_1_  (.A(\V2/V1/V3/v2 [1]),
    .B(\V2/V1/V3/v3 [1]),
    .Z(\V2/V1/V3/A1/M2/s1 ));
 AND2_X1 \V2/V1/V3/A1/M2/M2/_0_  (.A1(\V2/V1/V3/A1/M2/s1 ),
    .A2(\V2/V1/V3/A1/c1 ),
    .ZN(\V2/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M2/M2/_1_  (.A(\V2/V1/V3/A1/M2/s1 ),
    .B(\V2/V1/V3/A1/c1 ),
    .Z(\V2/V1/V3/s1 [1]));
 OR2_X1 \V2/V1/V3/A1/M2/_0_  (.A1(\V2/V1/V3/A1/M2/c1 ),
    .A2(\V2/V1/V3/A1/M2/c2 ),
    .ZN(\V2/V1/V3/A1/c2 ));
 AND2_X1 \V2/V1/V3/A1/M3/M1/_0_  (.A1(\V2/V1/V3/v2 [2]),
    .A2(\V2/V1/V3/v3 [2]),
    .ZN(\V2/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M3/M1/_1_  (.A(\V2/V1/V3/v2 [2]),
    .B(\V2/V1/V3/v3 [2]),
    .Z(\V2/V1/V3/A1/M3/s1 ));
 AND2_X1 \V2/V1/V3/A1/M3/M2/_0_  (.A1(\V2/V1/V3/A1/M3/s1 ),
    .A2(\V2/V1/V3/A1/c2 ),
    .ZN(\V2/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M3/M2/_1_  (.A(\V2/V1/V3/A1/M3/s1 ),
    .B(\V2/V1/V3/A1/c2 ),
    .Z(\V2/V1/V3/s1 [2]));
 OR2_X1 \V2/V1/V3/A1/M3/_0_  (.A1(\V2/V1/V3/A1/M3/c1 ),
    .A2(\V2/V1/V3/A1/M3/c2 ),
    .ZN(\V2/V1/V3/A1/c3 ));
 AND2_X1 \V2/V1/V3/A1/M4/M1/_0_  (.A1(\V2/V1/V3/v2 [3]),
    .A2(\V2/V1/V3/v3 [3]),
    .ZN(\V2/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A1/M4/M1/_1_  (.A(\V2/V1/V3/v2 [3]),
    .B(\V2/V1/V3/v3 [3]),
    .Z(\V2/V1/V3/A1/M4/s1 ));
 AND2_X1 \V2/V1/V3/A1/M4/M2/_0_  (.A1(\V2/V1/V3/A1/M4/s1 ),
    .A2(\V2/V1/V3/A1/c3 ),
    .ZN(\V2/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A1/M4/M2/_1_  (.A(\V2/V1/V3/A1/M4/s1 ),
    .B(\V2/V1/V3/A1/c3 ),
    .Z(\V2/V1/V3/s1 [3]));
 OR2_X1 \V2/V1/V3/A1/M4/_0_  (.A1(\V2/V1/V3/A1/M4/c1 ),
    .A2(\V2/V1/V3/A1/M4/c2 ),
    .ZN(\V2/V1/V3/c1 ));
 AND2_X1 \V2/V1/V3/A2/M1/M1/_0_  (.A1(\V2/V1/V3/s1 [0]),
    .A2(\V2/V1/V3/v1 [2]),
    .ZN(\V2/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M1/M1/_1_  (.A(\V2/V1/V3/s1 [0]),
    .B(\V2/V1/V3/v1 [2]),
    .Z(\V2/V1/V3/A2/M1/s1 ));
 AND2_X1 \V2/V1/V3/A2/M1/M2/_0_  (.A1(\V2/V1/V3/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M1/M2/_1_  (.A(\V2/V1/V3/A2/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/v3 [2]));
 OR2_X1 \V2/V1/V3/A2/M1/_0_  (.A1(\V2/V1/V3/A2/M1/c1 ),
    .A2(\V2/V1/V3/A2/M1/c2 ),
    .ZN(\V2/V1/V3/A2/c1 ));
 AND2_X1 \V2/V1/V3/A2/M2/M1/_0_  (.A1(\V2/V1/V3/s1 [1]),
    .A2(\V2/V1/V3/v1 [3]),
    .ZN(\V2/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M2/M1/_1_  (.A(\V2/V1/V3/s1 [1]),
    .B(\V2/V1/V3/v1 [3]),
    .Z(\V2/V1/V3/A2/M2/s1 ));
 AND2_X1 \V2/V1/V3/A2/M2/M2/_0_  (.A1(\V2/V1/V3/A2/M2/s1 ),
    .A2(\V2/V1/V3/A2/c1 ),
    .ZN(\V2/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M2/M2/_1_  (.A(\V2/V1/V3/A2/M2/s1 ),
    .B(\V2/V1/V3/A2/c1 ),
    .Z(\V2/V1/v3 [3]));
 OR2_X1 \V2/V1/V3/A2/M2/_0_  (.A1(\V2/V1/V3/A2/M2/c1 ),
    .A2(\V2/V1/V3/A2/M2/c2 ),
    .ZN(\V2/V1/V3/A2/c2 ));
 AND2_X1 \V2/V1/V3/A2/M3/M1/_0_  (.A1(\V2/V1/V3/s1 [2]),
    .A2(net4),
    .ZN(\V2/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M3/M1/_1_  (.A(\V2/V1/V3/s1 [2]),
    .B(net4),
    .Z(\V2/V1/V3/A2/M3/s1 ));
 AND2_X1 \V2/V1/V3/A2/M3/M2/_0_  (.A1(\V2/V1/V3/A2/M3/s1 ),
    .A2(\V2/V1/V3/A2/c2 ),
    .ZN(\V2/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M3/M2/_1_  (.A(\V2/V1/V3/A2/M3/s1 ),
    .B(\V2/V1/V3/A2/c2 ),
    .Z(\V2/V1/V3/s2 [2]));
 OR2_X1 \V2/V1/V3/A2/M3/_0_  (.A1(\V2/V1/V3/A2/M3/c1 ),
    .A2(\V2/V1/V3/A2/M3/c2 ),
    .ZN(\V2/V1/V3/A2/c3 ));
 AND2_X1 \V2/V1/V3/A2/M4/M1/_0_  (.A1(\V2/V1/V3/s1 [3]),
    .A2(net4),
    .ZN(\V2/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A2/M4/M1/_1_  (.A(\V2/V1/V3/s1 [3]),
    .B(net4),
    .Z(\V2/V1/V3/A2/M4/s1 ));
 AND2_X1 \V2/V1/V3/A2/M4/M2/_0_  (.A1(\V2/V1/V3/A2/M4/s1 ),
    .A2(\V2/V1/V3/A2/c3 ),
    .ZN(\V2/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A2/M4/M2/_1_  (.A(\V2/V1/V3/A2/M4/s1 ),
    .B(\V2/V1/V3/A2/c3 ),
    .Z(\V2/V1/V3/s2 [3]));
 OR2_X1 \V2/V1/V3/A2/M4/_0_  (.A1(\V2/V1/V3/A2/M4/c1 ),
    .A2(\V2/V1/V3/A2/M4/c2 ),
    .ZN(\V2/V1/V3/c2 ));
 AND2_X1 \V2/V1/V3/A3/M1/M1/_0_  (.A1(\V2/V1/V3/v4 [0]),
    .A2(\V2/V1/V3/s2 [2]),
    .ZN(\V2/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M1/M1/_1_  (.A(\V2/V1/V3/v4 [0]),
    .B(\V2/V1/V3/s2 [2]),
    .Z(\V2/V1/V3/A3/M1/s1 ));
 AND2_X1 \V2/V1/V3/A3/M1/M2/_0_  (.A1(\V2/V1/V3/A3/M1/s1 ),
    .A2(net4),
    .ZN(\V2/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M1/M2/_1_  (.A(\V2/V1/V3/A3/M1/s1 ),
    .B(net4),
    .Z(\V2/V1/v3 [4]));
 OR2_X1 \V2/V1/V3/A3/M1/_0_  (.A1(\V2/V1/V3/A3/M1/c1 ),
    .A2(\V2/V1/V3/A3/M1/c2 ),
    .ZN(\V2/V1/V3/A3/c1 ));
 AND2_X1 \V2/V1/V3/A3/M2/M1/_0_  (.A1(\V2/V1/V3/v4 [1]),
    .A2(\V2/V1/V3/s2 [3]),
    .ZN(\V2/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M2/M1/_1_  (.A(\V2/V1/V3/v4 [1]),
    .B(\V2/V1/V3/s2 [3]),
    .Z(\V2/V1/V3/A3/M2/s1 ));
 AND2_X1 \V2/V1/V3/A3/M2/M2/_0_  (.A1(\V2/V1/V3/A3/M2/s1 ),
    .A2(\V2/V1/V3/A3/c1 ),
    .ZN(\V2/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M2/M2/_1_  (.A(\V2/V1/V3/A3/M2/s1 ),
    .B(\V2/V1/V3/A3/c1 ),
    .Z(\V2/V1/v3 [5]));
 OR2_X1 \V2/V1/V3/A3/M2/_0_  (.A1(\V2/V1/V3/A3/M2/c1 ),
    .A2(\V2/V1/V3/A3/M2/c2 ),
    .ZN(\V2/V1/V3/A3/c2 ));
 AND2_X1 \V2/V1/V3/A3/M3/M1/_0_  (.A1(\V2/V1/V3/v4 [2]),
    .A2(\V2/V1/V3/c3 ),
    .ZN(\V2/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M3/M1/_1_  (.A(\V2/V1/V3/v4 [2]),
    .B(\V2/V1/V3/c3 ),
    .Z(\V2/V1/V3/A3/M3/s1 ));
 AND2_X1 \V2/V1/V3/A3/M3/M2/_0_  (.A1(\V2/V1/V3/A3/M3/s1 ),
    .A2(\V2/V1/V3/A3/c2 ),
    .ZN(\V2/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M3/M2/_1_  (.A(\V2/V1/V3/A3/M3/s1 ),
    .B(\V2/V1/V3/A3/c2 ),
    .Z(\V2/V1/v3 [6]));
 OR2_X1 \V2/V1/V3/A3/M3/_0_  (.A1(\V2/V1/V3/A3/M3/c1 ),
    .A2(\V2/V1/V3/A3/M3/c2 ),
    .ZN(\V2/V1/V3/A3/c3 ));
 AND2_X1 \V2/V1/V3/A3/M4/M1/_0_  (.A1(\V2/V1/V3/v4 [3]),
    .A2(net4),
    .ZN(\V2/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V3/A3/M4/M1/_1_  (.A(\V2/V1/V3/v4 [3]),
    .B(net4),
    .Z(\V2/V1/V3/A3/M4/s1 ));
 AND2_X1 \V2/V1/V3/A3/M4/M2/_0_  (.A1(\V2/V1/V3/A3/M4/s1 ),
    .A2(\V2/V1/V3/A3/c3 ),
    .ZN(\V2/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V3/A3/M4/M2/_1_  (.A(\V2/V1/V3/A3/M4/s1 ),
    .B(\V2/V1/V3/A3/c3 ),
    .Z(\V2/V1/v3 [7]));
 OR2_X1 \V2/V1/V3/A3/M4/_0_  (.A1(\V2/V1/V3/A3/M4/c1 ),
    .A2(\V2/V1/V3/A3/M4/c2 ),
    .ZN(\V2/V1/V3/overflow ));
 AND2_X1 \V2/V1/V3/V1/HA1/_0_  (.A1(\V2/V1/V3/V1/w2 ),
    .A2(\V2/V1/V3/V1/w1 ),
    .ZN(\V2/V1/V3/V1/w4 ));
 XOR2_X2 \V2/V1/V3/V1/HA1/_1_  (.A(\V2/V1/V3/V1/w2 ),
    .B(\V2/V1/V3/V1/w1 ),
    .Z(\V2/V1/v3 [1]));
 AND2_X1 \V2/V1/V3/V1/HA2/_0_  (.A1(\V2/V1/V3/V1/w4 ),
    .A2(\V2/V1/V3/V1/w3 ),
    .ZN(\V2/V1/V3/v1 [3]));
 XOR2_X2 \V2/V1/V3/V1/HA2/_1_  (.A(\V2/V1/V3/V1/w4 ),
    .B(\V2/V1/V3/V1/w3 ),
    .Z(\V2/V1/V3/v1 [2]));
 AND2_X1 \V2/V1/V3/V1/_0_  (.A1(net41),
    .A2(B[4]),
    .ZN(\V2/V1/v3 [0]));
 AND2_X1 \V2/V1/V3/V1/_1_  (.A1(net41),
    .A2(B[5]),
    .ZN(\V2/V1/V3/V1/w1 ));
 AND2_X1 \V2/V1/V3/V1/_2_  (.A1(B[4]),
    .A2(net40),
    .ZN(\V2/V1/V3/V1/w2 ));
 AND2_X1 \V2/V1/V3/V1/_3_  (.A1(B[5]),
    .A2(net40),
    .ZN(\V2/V1/V3/V1/w3 ));
 AND2_X1 \V2/V1/V3/V2/HA1/_0_  (.A1(\V2/V1/V3/V2/w2 ),
    .A2(\V2/V1/V3/V2/w1 ),
    .ZN(\V2/V1/V3/V2/w4 ));
 XOR2_X2 \V2/V1/V3/V2/HA1/_1_  (.A(\V2/V1/V3/V2/w2 ),
    .B(\V2/V1/V3/V2/w1 ),
    .Z(\V2/V1/V3/v2 [1]));
 AND2_X1 \V2/V1/V3/V2/HA2/_0_  (.A1(\V2/V1/V3/V2/w4 ),
    .A2(\V2/V1/V3/V2/w3 ),
    .ZN(\V2/V1/V3/v2 [3]));
 XOR2_X2 \V2/V1/V3/V2/HA2/_1_  (.A(\V2/V1/V3/V2/w4 ),
    .B(\V2/V1/V3/V2/w3 ),
    .Z(\V2/V1/V3/v2 [2]));
 AND2_X1 \V2/V1/V3/V2/_0_  (.A1(A[18]),
    .A2(B[4]),
    .ZN(\V2/V1/V3/v2 [0]));
 AND2_X1 \V2/V1/V3/V2/_1_  (.A1(A[18]),
    .A2(B[5]),
    .ZN(\V2/V1/V3/V2/w1 ));
 AND2_X1 \V2/V1/V3/V2/_2_  (.A1(B[4]),
    .A2(net38),
    .ZN(\V2/V1/V3/V2/w2 ));
 AND2_X1 \V2/V1/V3/V2/_3_  (.A1(B[5]),
    .A2(net38),
    .ZN(\V2/V1/V3/V2/w3 ));
 AND2_X1 \V2/V1/V3/V3/HA1/_0_  (.A1(\V2/V1/V3/V3/w2 ),
    .A2(\V2/V1/V3/V3/w1 ),
    .ZN(\V2/V1/V3/V3/w4 ));
 XOR2_X2 \V2/V1/V3/V3/HA1/_1_  (.A(\V2/V1/V3/V3/w2 ),
    .B(\V2/V1/V3/V3/w1 ),
    .Z(\V2/V1/V3/v3 [1]));
 AND2_X1 \V2/V1/V3/V3/HA2/_0_  (.A1(\V2/V1/V3/V3/w4 ),
    .A2(\V2/V1/V3/V3/w3 ),
    .ZN(\V2/V1/V3/v3 [3]));
 XOR2_X2 \V2/V1/V3/V3/HA2/_1_  (.A(\V2/V1/V3/V3/w4 ),
    .B(\V2/V1/V3/V3/w3 ),
    .Z(\V2/V1/V3/v3 [2]));
 AND2_X1 \V2/V1/V3/V3/_0_  (.A1(net41),
    .A2(B[6]),
    .ZN(\V2/V1/V3/v3 [0]));
 AND2_X1 \V2/V1/V3/V3/_1_  (.A1(net41),
    .A2(B[7]),
    .ZN(\V2/V1/V3/V3/w1 ));
 AND2_X1 \V2/V1/V3/V3/_2_  (.A1(B[6]),
    .A2(net40),
    .ZN(\V2/V1/V3/V3/w2 ));
 AND2_X1 \V2/V1/V3/V3/_3_  (.A1(B[7]),
    .A2(net40),
    .ZN(\V2/V1/V3/V3/w3 ));
 AND2_X1 \V2/V1/V3/V4/HA1/_0_  (.A1(\V2/V1/V3/V4/w2 ),
    .A2(\V2/V1/V3/V4/w1 ),
    .ZN(\V2/V1/V3/V4/w4 ));
 XOR2_X2 \V2/V1/V3/V4/HA1/_1_  (.A(\V2/V1/V3/V4/w2 ),
    .B(\V2/V1/V3/V4/w1 ),
    .Z(\V2/V1/V3/v4 [1]));
 AND2_X1 \V2/V1/V3/V4/HA2/_0_  (.A1(\V2/V1/V3/V4/w4 ),
    .A2(\V2/V1/V3/V4/w3 ),
    .ZN(\V2/V1/V3/v4 [3]));
 XOR2_X2 \V2/V1/V3/V4/HA2/_1_  (.A(\V2/V1/V3/V4/w4 ),
    .B(\V2/V1/V3/V4/w3 ),
    .Z(\V2/V1/V3/v4 [2]));
 AND2_X1 \V2/V1/V3/V4/_0_  (.A1(net39),
    .A2(B[6]),
    .ZN(\V2/V1/V3/v4 [0]));
 AND2_X1 \V2/V1/V3/V4/_1_  (.A1(net39),
    .A2(B[7]),
    .ZN(\V2/V1/V3/V4/w1 ));
 AND2_X1 \V2/V1/V3/V4/_2_  (.A1(B[6]),
    .A2(net38),
    .ZN(\V2/V1/V3/V4/w2 ));
 AND2_X1 \V2/V1/V3/V4/_3_  (.A1(B[7]),
    .A2(net38),
    .ZN(\V2/V1/V3/V4/w3 ));
 OR2_X1 \V2/V1/V3/_0_  (.A1(\V2/V1/V3/c1 ),
    .A2(\V2/V1/V3/c2 ),
    .ZN(\V2/V1/V3/c3 ));
 AND2_X1 \V2/V1/V4/A1/M1/M1/_0_  (.A1(\V2/V1/V4/v2 [0]),
    .A2(\V2/V1/V4/v3 [0]),
    .ZN(\V2/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M1/M1/_1_  (.A(\V2/V1/V4/v2 [0]),
    .B(\V2/V1/V4/v3 [0]),
    .Z(\V2/V1/V4/A1/M1/s1 ));
 AND2_X1 \V2/V1/V4/A1/M1/M2/_0_  (.A1(\V2/V1/V4/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M1/M2/_1_  (.A(\V2/V1/V4/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/V1/V4/s1 [0]));
 OR2_X1 \V2/V1/V4/A1/M1/_0_  (.A1(\V2/V1/V4/A1/M1/c1 ),
    .A2(\V2/V1/V4/A1/M1/c2 ),
    .ZN(\V2/V1/V4/A1/c1 ));
 AND2_X1 \V2/V1/V4/A1/M2/M1/_0_  (.A1(\V2/V1/V4/v2 [1]),
    .A2(\V2/V1/V4/v3 [1]),
    .ZN(\V2/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M2/M1/_1_  (.A(\V2/V1/V4/v2 [1]),
    .B(\V2/V1/V4/v3 [1]),
    .Z(\V2/V1/V4/A1/M2/s1 ));
 AND2_X1 \V2/V1/V4/A1/M2/M2/_0_  (.A1(\V2/V1/V4/A1/M2/s1 ),
    .A2(\V2/V1/V4/A1/c1 ),
    .ZN(\V2/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M2/M2/_1_  (.A(\V2/V1/V4/A1/M2/s1 ),
    .B(\V2/V1/V4/A1/c1 ),
    .Z(\V2/V1/V4/s1 [1]));
 OR2_X1 \V2/V1/V4/A1/M2/_0_  (.A1(\V2/V1/V4/A1/M2/c1 ),
    .A2(\V2/V1/V4/A1/M2/c2 ),
    .ZN(\V2/V1/V4/A1/c2 ));
 AND2_X1 \V2/V1/V4/A1/M3/M1/_0_  (.A1(\V2/V1/V4/v2 [2]),
    .A2(\V2/V1/V4/v3 [2]),
    .ZN(\V2/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M3/M1/_1_  (.A(\V2/V1/V4/v2 [2]),
    .B(\V2/V1/V4/v3 [2]),
    .Z(\V2/V1/V4/A1/M3/s1 ));
 AND2_X1 \V2/V1/V4/A1/M3/M2/_0_  (.A1(\V2/V1/V4/A1/M3/s1 ),
    .A2(\V2/V1/V4/A1/c2 ),
    .ZN(\V2/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M3/M2/_1_  (.A(\V2/V1/V4/A1/M3/s1 ),
    .B(\V2/V1/V4/A1/c2 ),
    .Z(\V2/V1/V4/s1 [2]));
 OR2_X1 \V2/V1/V4/A1/M3/_0_  (.A1(\V2/V1/V4/A1/M3/c1 ),
    .A2(\V2/V1/V4/A1/M3/c2 ),
    .ZN(\V2/V1/V4/A1/c3 ));
 AND2_X1 \V2/V1/V4/A1/M4/M1/_0_  (.A1(\V2/V1/V4/v2 [3]),
    .A2(\V2/V1/V4/v3 [3]),
    .ZN(\V2/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A1/M4/M1/_1_  (.A(\V2/V1/V4/v2 [3]),
    .B(\V2/V1/V4/v3 [3]),
    .Z(\V2/V1/V4/A1/M4/s1 ));
 AND2_X1 \V2/V1/V4/A1/M4/M2/_0_  (.A1(\V2/V1/V4/A1/M4/s1 ),
    .A2(\V2/V1/V4/A1/c3 ),
    .ZN(\V2/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A1/M4/M2/_1_  (.A(\V2/V1/V4/A1/M4/s1 ),
    .B(\V2/V1/V4/A1/c3 ),
    .Z(\V2/V1/V4/s1 [3]));
 OR2_X1 \V2/V1/V4/A1/M4/_0_  (.A1(\V2/V1/V4/A1/M4/c1 ),
    .A2(\V2/V1/V4/A1/M4/c2 ),
    .ZN(\V2/V1/V4/c1 ));
 AND2_X1 \V2/V1/V4/A2/M1/M1/_0_  (.A1(\V2/V1/V4/s1 [0]),
    .A2(\V2/V1/V4/v1 [2]),
    .ZN(\V2/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M1/M1/_1_  (.A(\V2/V1/V4/s1 [0]),
    .B(\V2/V1/V4/v1 [2]),
    .Z(\V2/V1/V4/A2/M1/s1 ));
 AND2_X1 \V2/V1/V4/A2/M1/M2/_0_  (.A1(\V2/V1/V4/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M1/M2/_1_  (.A(\V2/V1/V4/A2/M1/s1 ),
    .B(net2),
    .Z(\V2/V1/v4 [2]));
 OR2_X1 \V2/V1/V4/A2/M1/_0_  (.A1(\V2/V1/V4/A2/M1/c1 ),
    .A2(\V2/V1/V4/A2/M1/c2 ),
    .ZN(\V2/V1/V4/A2/c1 ));
 AND2_X1 \V2/V1/V4/A2/M2/M1/_0_  (.A1(\V2/V1/V4/s1 [1]),
    .A2(\V2/V1/V4/v1 [3]),
    .ZN(\V2/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M2/M1/_1_  (.A(\V2/V1/V4/s1 [1]),
    .B(\V2/V1/V4/v1 [3]),
    .Z(\V2/V1/V4/A2/M2/s1 ));
 AND2_X1 \V2/V1/V4/A2/M2/M2/_0_  (.A1(\V2/V1/V4/A2/M2/s1 ),
    .A2(\V2/V1/V4/A2/c1 ),
    .ZN(\V2/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M2/M2/_1_  (.A(\V2/V1/V4/A2/M2/s1 ),
    .B(\V2/V1/V4/A2/c1 ),
    .Z(\V2/V1/v4 [3]));
 OR2_X1 \V2/V1/V4/A2/M2/_0_  (.A1(\V2/V1/V4/A2/M2/c1 ),
    .A2(\V2/V1/V4/A2/M2/c2 ),
    .ZN(\V2/V1/V4/A2/c2 ));
 AND2_X1 \V2/V1/V4/A2/M3/M1/_0_  (.A1(\V2/V1/V4/s1 [2]),
    .A2(net2),
    .ZN(\V2/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M3/M1/_1_  (.A(\V2/V1/V4/s1 [2]),
    .B(net2),
    .Z(\V2/V1/V4/A2/M3/s1 ));
 AND2_X1 \V2/V1/V4/A2/M3/M2/_0_  (.A1(\V2/V1/V4/A2/M3/s1 ),
    .A2(\V2/V1/V4/A2/c2 ),
    .ZN(\V2/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M3/M2/_1_  (.A(\V2/V1/V4/A2/M3/s1 ),
    .B(\V2/V1/V4/A2/c2 ),
    .Z(\V2/V1/V4/s2 [2]));
 OR2_X1 \V2/V1/V4/A2/M3/_0_  (.A1(\V2/V1/V4/A2/M3/c1 ),
    .A2(\V2/V1/V4/A2/M3/c2 ),
    .ZN(\V2/V1/V4/A2/c3 ));
 AND2_X1 \V2/V1/V4/A2/M4/M1/_0_  (.A1(\V2/V1/V4/s1 [3]),
    .A2(net2),
    .ZN(\V2/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A2/M4/M1/_1_  (.A(\V2/V1/V4/s1 [3]),
    .B(net2),
    .Z(\V2/V1/V4/A2/M4/s1 ));
 AND2_X1 \V2/V1/V4/A2/M4/M2/_0_  (.A1(\V2/V1/V4/A2/M4/s1 ),
    .A2(\V2/V1/V4/A2/c3 ),
    .ZN(\V2/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A2/M4/M2/_1_  (.A(\V2/V1/V4/A2/M4/s1 ),
    .B(\V2/V1/V4/A2/c3 ),
    .Z(\V2/V1/V4/s2 [3]));
 OR2_X1 \V2/V1/V4/A2/M4/_0_  (.A1(\V2/V1/V4/A2/M4/c1 ),
    .A2(\V2/V1/V4/A2/M4/c2 ),
    .ZN(\V2/V1/V4/c2 ));
 AND2_X1 \V2/V1/V4/A3/M1/M1/_0_  (.A1(\V2/V1/V4/v4 [0]),
    .A2(\V2/V1/V4/s2 [2]),
    .ZN(\V2/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M1/M1/_1_  (.A(\V2/V1/V4/v4 [0]),
    .B(\V2/V1/V4/s2 [2]),
    .Z(\V2/V1/V4/A3/M1/s1 ));
 AND2_X1 \V2/V1/V4/A3/M1/M2/_0_  (.A1(\V2/V1/V4/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M1/M2/_1_  (.A(\V2/V1/V4/A3/M1/s1 ),
    .B(net2),
    .Z(\V2/V1/v4 [4]));
 OR2_X1 \V2/V1/V4/A3/M1/_0_  (.A1(\V2/V1/V4/A3/M1/c1 ),
    .A2(\V2/V1/V4/A3/M1/c2 ),
    .ZN(\V2/V1/V4/A3/c1 ));
 AND2_X1 \V2/V1/V4/A3/M2/M1/_0_  (.A1(\V2/V1/V4/v4 [1]),
    .A2(\V2/V1/V4/s2 [3]),
    .ZN(\V2/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M2/M1/_1_  (.A(\V2/V1/V4/v4 [1]),
    .B(\V2/V1/V4/s2 [3]),
    .Z(\V2/V1/V4/A3/M2/s1 ));
 AND2_X1 \V2/V1/V4/A3/M2/M2/_0_  (.A1(\V2/V1/V4/A3/M2/s1 ),
    .A2(\V2/V1/V4/A3/c1 ),
    .ZN(\V2/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M2/M2/_1_  (.A(\V2/V1/V4/A3/M2/s1 ),
    .B(\V2/V1/V4/A3/c1 ),
    .Z(\V2/V1/v4 [5]));
 OR2_X1 \V2/V1/V4/A3/M2/_0_  (.A1(\V2/V1/V4/A3/M2/c1 ),
    .A2(\V2/V1/V4/A3/M2/c2 ),
    .ZN(\V2/V1/V4/A3/c2 ));
 AND2_X1 \V2/V1/V4/A3/M3/M1/_0_  (.A1(\V2/V1/V4/v4 [2]),
    .A2(\V2/V1/V4/c3 ),
    .ZN(\V2/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M3/M1/_1_  (.A(\V2/V1/V4/v4 [2]),
    .B(\V2/V1/V4/c3 ),
    .Z(\V2/V1/V4/A3/M3/s1 ));
 AND2_X1 \V2/V1/V4/A3/M3/M2/_0_  (.A1(\V2/V1/V4/A3/M3/s1 ),
    .A2(\V2/V1/V4/A3/c2 ),
    .ZN(\V2/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M3/M2/_1_  (.A(\V2/V1/V4/A3/M3/s1 ),
    .B(\V2/V1/V4/A3/c2 ),
    .Z(\V2/V1/v4 [6]));
 OR2_X1 \V2/V1/V4/A3/M3/_0_  (.A1(\V2/V1/V4/A3/M3/c1 ),
    .A2(\V2/V1/V4/A3/M3/c2 ),
    .ZN(\V2/V1/V4/A3/c3 ));
 AND2_X1 \V2/V1/V4/A3/M4/M1/_0_  (.A1(\V2/V1/V4/v4 [3]),
    .A2(net2),
    .ZN(\V2/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V1/V4/A3/M4/M1/_1_  (.A(\V2/V1/V4/v4 [3]),
    .B(net2),
    .Z(\V2/V1/V4/A3/M4/s1 ));
 AND2_X1 \V2/V1/V4/A3/M4/M2/_0_  (.A1(\V2/V1/V4/A3/M4/s1 ),
    .A2(\V2/V1/V4/A3/c3 ),
    .ZN(\V2/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V1/V4/A3/M4/M2/_1_  (.A(\V2/V1/V4/A3/M4/s1 ),
    .B(\V2/V1/V4/A3/c3 ),
    .Z(\V2/V1/v4 [7]));
 OR2_X1 \V2/V1/V4/A3/M4/_0_  (.A1(\V2/V1/V4/A3/M4/c1 ),
    .A2(\V2/V1/V4/A3/M4/c2 ),
    .ZN(\V2/V1/V4/overflow ));
 AND2_X1 \V2/V1/V4/V1/HA1/_0_  (.A1(\V2/V1/V4/V1/w2 ),
    .A2(\V2/V1/V4/V1/w1 ),
    .ZN(\V2/V1/V4/V1/w4 ));
 XOR2_X2 \V2/V1/V4/V1/HA1/_1_  (.A(\V2/V1/V4/V1/w2 ),
    .B(\V2/V1/V4/V1/w1 ),
    .Z(\V2/V1/v4 [1]));
 AND2_X1 \V2/V1/V4/V1/HA2/_0_  (.A1(\V2/V1/V4/V1/w4 ),
    .A2(\V2/V1/V4/V1/w3 ),
    .ZN(\V2/V1/V4/v1 [3]));
 XOR2_X2 \V2/V1/V4/V1/HA2/_1_  (.A(\V2/V1/V4/V1/w4 ),
    .B(\V2/V1/V4/V1/w3 ),
    .Z(\V2/V1/V4/v1 [2]));
 AND2_X1 \V2/V1/V4/V1/_0_  (.A1(net37),
    .A2(B[4]),
    .ZN(\V2/V1/v4 [0]));
 AND2_X1 \V2/V1/V4/V1/_1_  (.A1(net37),
    .A2(B[5]),
    .ZN(\V2/V1/V4/V1/w1 ));
 AND2_X1 \V2/V1/V4/V1/_2_  (.A1(B[4]),
    .A2(net36),
    .ZN(\V2/V1/V4/V1/w2 ));
 AND2_X1 \V2/V1/V4/V1/_3_  (.A1(B[5]),
    .A2(net36),
    .ZN(\V2/V1/V4/V1/w3 ));
 AND2_X1 \V2/V1/V4/V2/HA1/_0_  (.A1(\V2/V1/V4/V2/w2 ),
    .A2(\V2/V1/V4/V2/w1 ),
    .ZN(\V2/V1/V4/V2/w4 ));
 XOR2_X2 \V2/V1/V4/V2/HA1/_1_  (.A(\V2/V1/V4/V2/w2 ),
    .B(\V2/V1/V4/V2/w1 ),
    .Z(\V2/V1/V4/v2 [1]));
 AND2_X1 \V2/V1/V4/V2/HA2/_0_  (.A1(\V2/V1/V4/V2/w4 ),
    .A2(\V2/V1/V4/V2/w3 ),
    .ZN(\V2/V1/V4/v2 [3]));
 XOR2_X2 \V2/V1/V4/V2/HA2/_1_  (.A(\V2/V1/V4/V2/w4 ),
    .B(\V2/V1/V4/V2/w3 ),
    .Z(\V2/V1/V4/v2 [2]));
 AND2_X1 \V2/V1/V4/V2/_0_  (.A1(net35),
    .A2(B[4]),
    .ZN(\V2/V1/V4/v2 [0]));
 AND2_X1 \V2/V1/V4/V2/_1_  (.A1(net35),
    .A2(B[5]),
    .ZN(\V2/V1/V4/V2/w1 ));
 AND2_X1 \V2/V1/V4/V2/_2_  (.A1(B[4]),
    .A2(net34),
    .ZN(\V2/V1/V4/V2/w2 ));
 AND2_X1 \V2/V1/V4/V2/_3_  (.A1(B[5]),
    .A2(net34),
    .ZN(\V2/V1/V4/V2/w3 ));
 AND2_X1 \V2/V1/V4/V3/HA1/_0_  (.A1(\V2/V1/V4/V3/w2 ),
    .A2(\V2/V1/V4/V3/w1 ),
    .ZN(\V2/V1/V4/V3/w4 ));
 XOR2_X2 \V2/V1/V4/V3/HA1/_1_  (.A(\V2/V1/V4/V3/w2 ),
    .B(\V2/V1/V4/V3/w1 ),
    .Z(\V2/V1/V4/v3 [1]));
 AND2_X1 \V2/V1/V4/V3/HA2/_0_  (.A1(\V2/V1/V4/V3/w4 ),
    .A2(\V2/V1/V4/V3/w3 ),
    .ZN(\V2/V1/V4/v3 [3]));
 XOR2_X2 \V2/V1/V4/V3/HA2/_1_  (.A(\V2/V1/V4/V3/w4 ),
    .B(\V2/V1/V4/V3/w3 ),
    .Z(\V2/V1/V4/v3 [2]));
 AND2_X1 \V2/V1/V4/V3/_0_  (.A1(net37),
    .A2(B[6]),
    .ZN(\V2/V1/V4/v3 [0]));
 AND2_X1 \V2/V1/V4/V3/_1_  (.A1(net37),
    .A2(B[7]),
    .ZN(\V2/V1/V4/V3/w1 ));
 AND2_X1 \V2/V1/V4/V3/_2_  (.A1(B[6]),
    .A2(net36),
    .ZN(\V2/V1/V4/V3/w2 ));
 AND2_X1 \V2/V1/V4/V3/_3_  (.A1(B[7]),
    .A2(net36),
    .ZN(\V2/V1/V4/V3/w3 ));
 AND2_X1 \V2/V1/V4/V4/HA1/_0_  (.A1(\V2/V1/V4/V4/w2 ),
    .A2(\V2/V1/V4/V4/w1 ),
    .ZN(\V2/V1/V4/V4/w4 ));
 XOR2_X2 \V2/V1/V4/V4/HA1/_1_  (.A(\V2/V1/V4/V4/w2 ),
    .B(\V2/V1/V4/V4/w1 ),
    .Z(\V2/V1/V4/v4 [1]));
 AND2_X1 \V2/V1/V4/V4/HA2/_0_  (.A1(\V2/V1/V4/V4/w4 ),
    .A2(\V2/V1/V4/V4/w3 ),
    .ZN(\V2/V1/V4/v4 [3]));
 XOR2_X2 \V2/V1/V4/V4/HA2/_1_  (.A(\V2/V1/V4/V4/w4 ),
    .B(\V2/V1/V4/V4/w3 ),
    .Z(\V2/V1/V4/v4 [2]));
 AND2_X1 \V2/V1/V4/V4/_0_  (.A1(net35),
    .A2(B[6]),
    .ZN(\V2/V1/V4/v4 [0]));
 AND2_X1 \V2/V1/V4/V4/_1_  (.A1(net35),
    .A2(B[7]),
    .ZN(\V2/V1/V4/V4/w1 ));
 AND2_X1 \V2/V1/V4/V4/_2_  (.A1(B[6]),
    .A2(net34),
    .ZN(\V2/V1/V4/V4/w2 ));
 AND2_X1 \V2/V1/V4/V4/_3_  (.A1(B[7]),
    .A2(net34),
    .ZN(\V2/V1/V4/V4/w3 ));
 OR2_X1 \V2/V1/V4/_0_  (.A1(\V2/V1/V4/c1 ),
    .A2(\V2/V1/V4/c2 ),
    .ZN(\V2/V1/V4/c3 ));
 OR2_X2 \V2/V1/_0_  (.A1(\V2/V1/c1 ),
    .A2(\V2/V1/c2 ),
    .ZN(\V2/V1/c3 ));
 AND2_X1 \V2/V2/A1/A1/M1/M1/_0_  (.A1(\V2/V2/v2 [0]),
    .A2(\V2/V2/v3 [0]),
    .ZN(\V2/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M1/M1/_1_  (.A(\V2/V2/v2 [0]),
    .B(\V2/V2/v3 [0]),
    .Z(\V2/V2/A1/A1/M1/s1 ));
 AND2_X1 \V2/V2/A1/A1/M1/M2/_0_  (.A1(\V2/V2/A1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M1/M2/_1_  (.A(\V2/V2/A1/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/V2/s1 [0]));
 OR2_X1 \V2/V2/A1/A1/M1/_0_  (.A1(\V2/V2/A1/A1/M1/c1 ),
    .A2(\V2/V2/A1/A1/M1/c2 ),
    .ZN(\V2/V2/A1/A1/c1 ));
 AND2_X1 \V2/V2/A1/A1/M2/M1/_0_  (.A1(\V2/V2/v2 [1]),
    .A2(\V2/V2/v3 [1]),
    .ZN(\V2/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M2/M1/_1_  (.A(\V2/V2/v2 [1]),
    .B(\V2/V2/v3 [1]),
    .Z(\V2/V2/A1/A1/M2/s1 ));
 AND2_X1 \V2/V2/A1/A1/M2/M2/_0_  (.A1(\V2/V2/A1/A1/M2/s1 ),
    .A2(\V2/V2/A1/A1/c1 ),
    .ZN(\V2/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M2/M2/_1_  (.A(\V2/V2/A1/A1/M2/s1 ),
    .B(\V2/V2/A1/A1/c1 ),
    .Z(\V2/V2/s1 [1]));
 OR2_X1 \V2/V2/A1/A1/M2/_0_  (.A1(\V2/V2/A1/A1/M2/c1 ),
    .A2(\V2/V2/A1/A1/M2/c2 ),
    .ZN(\V2/V2/A1/A1/c2 ));
 AND2_X1 \V2/V2/A1/A1/M3/M1/_0_  (.A1(\V2/V2/v2 [2]),
    .A2(\V2/V2/v3 [2]),
    .ZN(\V2/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M3/M1/_1_  (.A(\V2/V2/v2 [2]),
    .B(\V2/V2/v3 [2]),
    .Z(\V2/V2/A1/A1/M3/s1 ));
 AND2_X1 \V2/V2/A1/A1/M3/M2/_0_  (.A1(\V2/V2/A1/A1/M3/s1 ),
    .A2(\V2/V2/A1/A1/c2 ),
    .ZN(\V2/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M3/M2/_1_  (.A(\V2/V2/A1/A1/M3/s1 ),
    .B(\V2/V2/A1/A1/c2 ),
    .Z(\V2/V2/s1 [2]));
 OR2_X1 \V2/V2/A1/A1/M3/_0_  (.A1(\V2/V2/A1/A1/M3/c1 ),
    .A2(\V2/V2/A1/A1/M3/c2 ),
    .ZN(\V2/V2/A1/A1/c3 ));
 AND2_X1 \V2/V2/A1/A1/M4/M1/_0_  (.A1(\V2/V2/v2 [3]),
    .A2(\V2/V2/v3 [3]),
    .ZN(\V2/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A1/A1/M4/M1/_1_  (.A(\V2/V2/v2 [3]),
    .B(\V2/V2/v3 [3]),
    .Z(\V2/V2/A1/A1/M4/s1 ));
 AND2_X1 \V2/V2/A1/A1/M4/M2/_0_  (.A1(\V2/V2/A1/A1/M4/s1 ),
    .A2(\V2/V2/A1/A1/c3 ),
    .ZN(\V2/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A1/A1/M4/M2/_1_  (.A(\V2/V2/A1/A1/M4/s1 ),
    .B(\V2/V2/A1/A1/c3 ),
    .Z(\V2/V2/s1 [3]));
 OR2_X1 \V2/V2/A1/A1/M4/_0_  (.A1(\V2/V2/A1/A1/M4/c1 ),
    .A2(\V2/V2/A1/A1/M4/c2 ),
    .ZN(\V2/V2/A1/c1 ));
 AND2_X1 \V2/V2/A1/A2/M1/M1/_0_  (.A1(\V2/V2/v2 [4]),
    .A2(\V2/V2/v3 [4]),
    .ZN(\V2/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M1/M1/_1_  (.A(\V2/V2/v2 [4]),
    .B(\V2/V2/v3 [4]),
    .Z(\V2/V2/A1/A2/M1/s1 ));
 AND2_X1 \V2/V2/A1/A2/M1/M2/_0_  (.A1(\V2/V2/A1/A2/M1/s1 ),
    .A2(\V2/V2/A1/c1 ),
    .ZN(\V2/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M1/M2/_1_  (.A(\V2/V2/A1/A2/M1/s1 ),
    .B(\V2/V2/A1/c1 ),
    .Z(\V2/V2/s1 [4]));
 OR2_X1 \V2/V2/A1/A2/M1/_0_  (.A1(\V2/V2/A1/A2/M1/c1 ),
    .A2(\V2/V2/A1/A2/M1/c2 ),
    .ZN(\V2/V2/A1/A2/c1 ));
 AND2_X1 \V2/V2/A1/A2/M2/M1/_0_  (.A1(\V2/V2/v2 [5]),
    .A2(\V2/V2/v3 [5]),
    .ZN(\V2/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M2/M1/_1_  (.A(\V2/V2/v2 [5]),
    .B(\V2/V2/v3 [5]),
    .Z(\V2/V2/A1/A2/M2/s1 ));
 AND2_X1 \V2/V2/A1/A2/M2/M2/_0_  (.A1(\V2/V2/A1/A2/M2/s1 ),
    .A2(\V2/V2/A1/A2/c1 ),
    .ZN(\V2/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M2/M2/_1_  (.A(\V2/V2/A1/A2/M2/s1 ),
    .B(\V2/V2/A1/A2/c1 ),
    .Z(\V2/V2/s1 [5]));
 OR2_X1 \V2/V2/A1/A2/M2/_0_  (.A1(\V2/V2/A1/A2/M2/c1 ),
    .A2(\V2/V2/A1/A2/M2/c2 ),
    .ZN(\V2/V2/A1/A2/c2 ));
 AND2_X1 \V2/V2/A1/A2/M3/M1/_0_  (.A1(\V2/V2/v2 [6]),
    .A2(\V2/V2/v3 [6]),
    .ZN(\V2/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M3/M1/_1_  (.A(\V2/V2/v2 [6]),
    .B(\V2/V2/v3 [6]),
    .Z(\V2/V2/A1/A2/M3/s1 ));
 AND2_X1 \V2/V2/A1/A2/M3/M2/_0_  (.A1(\V2/V2/A1/A2/M3/s1 ),
    .A2(\V2/V2/A1/A2/c2 ),
    .ZN(\V2/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M3/M2/_1_  (.A(\V2/V2/A1/A2/M3/s1 ),
    .B(\V2/V2/A1/A2/c2 ),
    .Z(\V2/V2/s1 [6]));
 OR2_X1 \V2/V2/A1/A2/M3/_0_  (.A1(\V2/V2/A1/A2/M3/c1 ),
    .A2(\V2/V2/A1/A2/M3/c2 ),
    .ZN(\V2/V2/A1/A2/c3 ));
 AND2_X1 \V2/V2/A1/A2/M4/M1/_0_  (.A1(\V2/V2/v2 [7]),
    .A2(\V2/V2/v3 [7]),
    .ZN(\V2/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A1/A2/M4/M1/_1_  (.A(\V2/V2/v2 [7]),
    .B(\V2/V2/v3 [7]),
    .Z(\V2/V2/A1/A2/M4/s1 ));
 AND2_X1 \V2/V2/A1/A2/M4/M2/_0_  (.A1(\V2/V2/A1/A2/M4/s1 ),
    .A2(\V2/V2/A1/A2/c3 ),
    .ZN(\V2/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A1/A2/M4/M2/_1_  (.A(\V2/V2/A1/A2/M4/s1 ),
    .B(\V2/V2/A1/A2/c3 ),
    .Z(\V2/V2/s1 [7]));
 OR2_X1 \V2/V2/A1/A2/M4/_0_  (.A1(\V2/V2/A1/A2/M4/c1 ),
    .A2(\V2/V2/A1/A2/M4/c2 ),
    .ZN(\V2/V2/c1 ));
 AND2_X1 \V2/V2/A2/A1/M1/M1/_0_  (.A1(\V2/V2/s1 [0]),
    .A2(\V2/V2/v1 [4]),
    .ZN(\V2/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M1/M1/_1_  (.A(\V2/V2/s1 [0]),
    .B(\V2/V2/v1 [4]),
    .Z(\V2/V2/A2/A1/M1/s1 ));
 AND2_X1 \V2/V2/A2/A1/M1/M2/_0_  (.A1(\V2/V2/A2/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M1/M2/_1_  (.A(\V2/V2/A2/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/v2 [4]));
 OR2_X1 \V2/V2/A2/A1/M1/_0_  (.A1(\V2/V2/A2/A1/M1/c1 ),
    .A2(\V2/V2/A2/A1/M1/c2 ),
    .ZN(\V2/V2/A2/A1/c1 ));
 AND2_X1 \V2/V2/A2/A1/M2/M1/_0_  (.A1(\V2/V2/s1 [1]),
    .A2(\V2/V2/v1 [5]),
    .ZN(\V2/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M2/M1/_1_  (.A(\V2/V2/s1 [1]),
    .B(\V2/V2/v1 [5]),
    .Z(\V2/V2/A2/A1/M2/s1 ));
 AND2_X1 \V2/V2/A2/A1/M2/M2/_0_  (.A1(\V2/V2/A2/A1/M2/s1 ),
    .A2(\V2/V2/A2/A1/c1 ),
    .ZN(\V2/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M2/M2/_1_  (.A(\V2/V2/A2/A1/M2/s1 ),
    .B(\V2/V2/A2/A1/c1 ),
    .Z(\V2/v2 [5]));
 OR2_X1 \V2/V2/A2/A1/M2/_0_  (.A1(\V2/V2/A2/A1/M2/c1 ),
    .A2(\V2/V2/A2/A1/M2/c2 ),
    .ZN(\V2/V2/A2/A1/c2 ));
 AND2_X1 \V2/V2/A2/A1/M3/M1/_0_  (.A1(\V2/V2/s1 [2]),
    .A2(\V2/V2/v1 [6]),
    .ZN(\V2/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M3/M1/_1_  (.A(\V2/V2/s1 [2]),
    .B(\V2/V2/v1 [6]),
    .Z(\V2/V2/A2/A1/M3/s1 ));
 AND2_X1 \V2/V2/A2/A1/M3/M2/_0_  (.A1(\V2/V2/A2/A1/M3/s1 ),
    .A2(\V2/V2/A2/A1/c2 ),
    .ZN(\V2/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M3/M2/_1_  (.A(\V2/V2/A2/A1/M3/s1 ),
    .B(\V2/V2/A2/A1/c2 ),
    .Z(\V2/v2 [6]));
 OR2_X1 \V2/V2/A2/A1/M3/_0_  (.A1(\V2/V2/A2/A1/M3/c1 ),
    .A2(\V2/V2/A2/A1/M3/c2 ),
    .ZN(\V2/V2/A2/A1/c3 ));
 AND2_X1 \V2/V2/A2/A1/M4/M1/_0_  (.A1(\V2/V2/s1 [3]),
    .A2(\V2/V2/v1 [7]),
    .ZN(\V2/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A2/A1/M4/M1/_1_  (.A(\V2/V2/s1 [3]),
    .B(\V2/V2/v1 [7]),
    .Z(\V2/V2/A2/A1/M4/s1 ));
 AND2_X1 \V2/V2/A2/A1/M4/M2/_0_  (.A1(\V2/V2/A2/A1/M4/s1 ),
    .A2(\V2/V2/A2/A1/c3 ),
    .ZN(\V2/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A2/A1/M4/M2/_1_  (.A(\V2/V2/A2/A1/M4/s1 ),
    .B(\V2/V2/A2/A1/c3 ),
    .Z(\V2/v2 [7]));
 OR2_X1 \V2/V2/A2/A1/M4/_0_  (.A1(\V2/V2/A2/A1/M4/c1 ),
    .A2(\V2/V2/A2/A1/M4/c2 ),
    .ZN(\V2/V2/A2/c1 ));
 AND2_X1 \V2/V2/A2/A2/M1/M1/_0_  (.A1(\V2/V2/s1 [4]),
    .A2(net7),
    .ZN(\V2/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M1/M1/_1_  (.A(\V2/V2/s1 [4]),
    .B(net7),
    .Z(\V2/V2/A2/A2/M1/s1 ));
 AND2_X1 \V2/V2/A2/A2/M1/M2/_0_  (.A1(\V2/V2/A2/A2/M1/s1 ),
    .A2(\V2/V2/A2/c1 ),
    .ZN(\V2/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M1/M2/_1_  (.A(\V2/V2/A2/A2/M1/s1 ),
    .B(\V2/V2/A2/c1 ),
    .Z(\V2/V2/s2 [4]));
 OR2_X1 \V2/V2/A2/A2/M1/_0_  (.A1(\V2/V2/A2/A2/M1/c1 ),
    .A2(\V2/V2/A2/A2/M1/c2 ),
    .ZN(\V2/V2/A2/A2/c1 ));
 AND2_X1 \V2/V2/A2/A2/M2/M1/_0_  (.A1(\V2/V2/s1 [5]),
    .A2(net7),
    .ZN(\V2/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M2/M1/_1_  (.A(\V2/V2/s1 [5]),
    .B(net7),
    .Z(\V2/V2/A2/A2/M2/s1 ));
 AND2_X1 \V2/V2/A2/A2/M2/M2/_0_  (.A1(\V2/V2/A2/A2/M2/s1 ),
    .A2(\V2/V2/A2/A2/c1 ),
    .ZN(\V2/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M2/M2/_1_  (.A(\V2/V2/A2/A2/M2/s1 ),
    .B(\V2/V2/A2/A2/c1 ),
    .Z(\V2/V2/s2 [5]));
 OR2_X1 \V2/V2/A2/A2/M2/_0_  (.A1(\V2/V2/A2/A2/M2/c1 ),
    .A2(\V2/V2/A2/A2/M2/c2 ),
    .ZN(\V2/V2/A2/A2/c2 ));
 AND2_X1 \V2/V2/A2/A2/M3/M1/_0_  (.A1(\V2/V2/s1 [6]),
    .A2(net7),
    .ZN(\V2/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M3/M1/_1_  (.A(\V2/V2/s1 [6]),
    .B(net7),
    .Z(\V2/V2/A2/A2/M3/s1 ));
 AND2_X1 \V2/V2/A2/A2/M3/M2/_0_  (.A1(\V2/V2/A2/A2/M3/s1 ),
    .A2(\V2/V2/A2/A2/c2 ),
    .ZN(\V2/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M3/M2/_1_  (.A(\V2/V2/A2/A2/M3/s1 ),
    .B(\V2/V2/A2/A2/c2 ),
    .Z(\V2/V2/s2 [6]));
 OR2_X1 \V2/V2/A2/A2/M3/_0_  (.A1(\V2/V2/A2/A2/M3/c1 ),
    .A2(\V2/V2/A2/A2/M3/c2 ),
    .ZN(\V2/V2/A2/A2/c3 ));
 AND2_X1 \V2/V2/A2/A2/M4/M1/_0_  (.A1(\V2/V2/s1 [7]),
    .A2(net7),
    .ZN(\V2/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A2/A2/M4/M1/_1_  (.A(\V2/V2/s1 [7]),
    .B(net7),
    .Z(\V2/V2/A2/A2/M4/s1 ));
 AND2_X1 \V2/V2/A2/A2/M4/M2/_0_  (.A1(\V2/V2/A2/A2/M4/s1 ),
    .A2(\V2/V2/A2/A2/c3 ),
    .ZN(\V2/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A2/A2/M4/M2/_1_  (.A(\V2/V2/A2/A2/M4/s1 ),
    .B(\V2/V2/A2/A2/c3 ),
    .Z(\V2/V2/s2 [7]));
 OR2_X1 \V2/V2/A2/A2/M4/_0_  (.A1(\V2/V2/A2/A2/M4/c1 ),
    .A2(\V2/V2/A2/A2/M4/c2 ),
    .ZN(\V2/V2/c2 ));
 AND2_X1 \V2/V2/A3/A1/M1/M1/_0_  (.A1(\V2/V2/v4 [0]),
    .A2(\V2/V2/s2 [4]),
    .ZN(\V2/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M1/M1/_1_  (.A(\V2/V2/v4 [0]),
    .B(\V2/V2/s2 [4]),
    .Z(\V2/V2/A3/A1/M1/s1 ));
 AND2_X1 \V2/V2/A3/A1/M1/M2/_0_  (.A1(\V2/V2/A3/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M1/M2/_1_  (.A(\V2/V2/A3/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/v2 [8]));
 OR2_X1 \V2/V2/A3/A1/M1/_0_  (.A1(\V2/V2/A3/A1/M1/c1 ),
    .A2(\V2/V2/A3/A1/M1/c2 ),
    .ZN(\V2/V2/A3/A1/c1 ));
 AND2_X1 \V2/V2/A3/A1/M2/M1/_0_  (.A1(\V2/V2/v4 [1]),
    .A2(\V2/V2/s2 [5]),
    .ZN(\V2/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M2/M1/_1_  (.A(\V2/V2/v4 [1]),
    .B(\V2/V2/s2 [5]),
    .Z(\V2/V2/A3/A1/M2/s1 ));
 AND2_X1 \V2/V2/A3/A1/M2/M2/_0_  (.A1(\V2/V2/A3/A1/M2/s1 ),
    .A2(\V2/V2/A3/A1/c1 ),
    .ZN(\V2/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M2/M2/_1_  (.A(\V2/V2/A3/A1/M2/s1 ),
    .B(\V2/V2/A3/A1/c1 ),
    .Z(\V2/v2 [9]));
 OR2_X1 \V2/V2/A3/A1/M2/_0_  (.A1(\V2/V2/A3/A1/M2/c1 ),
    .A2(\V2/V2/A3/A1/M2/c2 ),
    .ZN(\V2/V2/A3/A1/c2 ));
 AND2_X1 \V2/V2/A3/A1/M3/M1/_0_  (.A1(\V2/V2/v4 [2]),
    .A2(\V2/V2/s2 [6]),
    .ZN(\V2/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M3/M1/_1_  (.A(\V2/V2/v4 [2]),
    .B(\V2/V2/s2 [6]),
    .Z(\V2/V2/A3/A1/M3/s1 ));
 AND2_X1 \V2/V2/A3/A1/M3/M2/_0_  (.A1(\V2/V2/A3/A1/M3/s1 ),
    .A2(\V2/V2/A3/A1/c2 ),
    .ZN(\V2/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M3/M2/_1_  (.A(\V2/V2/A3/A1/M3/s1 ),
    .B(\V2/V2/A3/A1/c2 ),
    .Z(\V2/v2 [10]));
 OR2_X1 \V2/V2/A3/A1/M3/_0_  (.A1(\V2/V2/A3/A1/M3/c1 ),
    .A2(\V2/V2/A3/A1/M3/c2 ),
    .ZN(\V2/V2/A3/A1/c3 ));
 AND2_X1 \V2/V2/A3/A1/M4/M1/_0_  (.A1(\V2/V2/v4 [3]),
    .A2(\V2/V2/s2 [7]),
    .ZN(\V2/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V2/A3/A1/M4/M1/_1_  (.A(\V2/V2/v4 [3]),
    .B(\V2/V2/s2 [7]),
    .Z(\V2/V2/A3/A1/M4/s1 ));
 AND2_X1 \V2/V2/A3/A1/M4/M2/_0_  (.A1(\V2/V2/A3/A1/M4/s1 ),
    .A2(\V2/V2/A3/A1/c3 ),
    .ZN(\V2/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V2/A3/A1/M4/M2/_1_  (.A(\V2/V2/A3/A1/M4/s1 ),
    .B(\V2/V2/A3/A1/c3 ),
    .Z(\V2/v2 [11]));
 OR2_X1 \V2/V2/A3/A1/M4/_0_  (.A1(\V2/V2/A3/A1/M4/c1 ),
    .A2(\V2/V2/A3/A1/M4/c2 ),
    .ZN(\V2/V2/A3/c1 ));
 AND2_X1 \V2/V2/A3/A2/M1/M1/_0_  (.A1(\V2/V2/v4 [4]),
    .A2(\V2/V2/c3 ),
    .ZN(\V2/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M1/M1/_1_  (.A(\V2/V2/v4 [4]),
    .B(\V2/V2/c3 ),
    .Z(\V2/V2/A3/A2/M1/s1 ));
 AND2_X1 \V2/V2/A3/A2/M1/M2/_0_  (.A1(\V2/V2/A3/A2/M1/s1 ),
    .A2(\V2/V2/A3/c1 ),
    .ZN(\V2/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M1/M2/_1_  (.A(\V2/V2/A3/A2/M1/s1 ),
    .B(\V2/V2/A3/c1 ),
    .Z(\V2/v2 [12]));
 OR2_X1 \V2/V2/A3/A2/M1/_0_  (.A1(\V2/V2/A3/A2/M1/c1 ),
    .A2(\V2/V2/A3/A2/M1/c2 ),
    .ZN(\V2/V2/A3/A2/c1 ));
 AND2_X1 \V2/V2/A3/A2/M2/M1/_0_  (.A1(\V2/V2/v4 [5]),
    .A2(net9),
    .ZN(\V2/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M2/M1/_1_  (.A(\V2/V2/v4 [5]),
    .B(net9),
    .Z(\V2/V2/A3/A2/M2/s1 ));
 AND2_X1 \V2/V2/A3/A2/M2/M2/_0_  (.A1(\V2/V2/A3/A2/M2/s1 ),
    .A2(\V2/V2/A3/A2/c1 ),
    .ZN(\V2/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M2/M2/_1_  (.A(\V2/V2/A3/A2/M2/s1 ),
    .B(\V2/V2/A3/A2/c1 ),
    .Z(\V2/v2 [13]));
 OR2_X1 \V2/V2/A3/A2/M2/_0_  (.A1(\V2/V2/A3/A2/M2/c1 ),
    .A2(\V2/V2/A3/A2/M2/c2 ),
    .ZN(\V2/V2/A3/A2/c2 ));
 AND2_X1 \V2/V2/A3/A2/M3/M1/_0_  (.A1(\V2/V2/v4 [6]),
    .A2(net9),
    .ZN(\V2/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M3/M1/_1_  (.A(\V2/V2/v4 [6]),
    .B(net9),
    .Z(\V2/V2/A3/A2/M3/s1 ));
 AND2_X1 \V2/V2/A3/A2/M3/M2/_0_  (.A1(\V2/V2/A3/A2/M3/s1 ),
    .A2(\V2/V2/A3/A2/c2 ),
    .ZN(\V2/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M3/M2/_1_  (.A(\V2/V2/A3/A2/M3/s1 ),
    .B(\V2/V2/A3/A2/c2 ),
    .Z(\V2/v2 [14]));
 OR2_X1 \V2/V2/A3/A2/M3/_0_  (.A1(\V2/V2/A3/A2/M3/c1 ),
    .A2(\V2/V2/A3/A2/M3/c2 ),
    .ZN(\V2/V2/A3/A2/c3 ));
 AND2_X1 \V2/V2/A3/A2/M4/M1/_0_  (.A1(\V2/V2/v4 [7]),
    .A2(net9),
    .ZN(\V2/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V2/A3/A2/M4/M1/_1_  (.A(\V2/V2/v4 [7]),
    .B(net9),
    .Z(\V2/V2/A3/A2/M4/s1 ));
 AND2_X1 \V2/V2/A3/A2/M4/M2/_0_  (.A1(\V2/V2/A3/A2/M4/s1 ),
    .A2(\V2/V2/A3/A2/c3 ),
    .ZN(\V2/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V2/A3/A2/M4/M2/_1_  (.A(\V2/V2/A3/A2/M4/s1 ),
    .B(\V2/V2/A3/A2/c3 ),
    .Z(\V2/v2 [15]));
 OR2_X1 \V2/V2/A3/A2/M4/_0_  (.A1(\V2/V2/A3/A2/M4/c1 ),
    .A2(\V2/V2/A3/A2/M4/c2 ),
    .ZN(\V2/V2/overflow ));
 AND2_X1 \V2/V2/V1/A1/M1/M1/_0_  (.A1(\V2/V2/V1/v2 [0]),
    .A2(\V2/V2/V1/v3 [0]),
    .ZN(\V2/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M1/M1/_1_  (.A(\V2/V2/V1/v2 [0]),
    .B(\V2/V2/V1/v3 [0]),
    .Z(\V2/V2/V1/A1/M1/s1 ));
 AND2_X1 \V2/V2/V1/A1/M1/M2/_0_  (.A1(\V2/V2/V1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M1/M2/_1_  (.A(\V2/V2/V1/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/V2/V1/s1 [0]));
 OR2_X1 \V2/V2/V1/A1/M1/_0_  (.A1(\V2/V2/V1/A1/M1/c1 ),
    .A2(\V2/V2/V1/A1/M1/c2 ),
    .ZN(\V2/V2/V1/A1/c1 ));
 AND2_X1 \V2/V2/V1/A1/M2/M1/_0_  (.A1(\V2/V2/V1/v2 [1]),
    .A2(\V2/V2/V1/v3 [1]),
    .ZN(\V2/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M2/M1/_1_  (.A(\V2/V2/V1/v2 [1]),
    .B(\V2/V2/V1/v3 [1]),
    .Z(\V2/V2/V1/A1/M2/s1 ));
 AND2_X1 \V2/V2/V1/A1/M2/M2/_0_  (.A1(\V2/V2/V1/A1/M2/s1 ),
    .A2(\V2/V2/V1/A1/c1 ),
    .ZN(\V2/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M2/M2/_1_  (.A(\V2/V2/V1/A1/M2/s1 ),
    .B(\V2/V2/V1/A1/c1 ),
    .Z(\V2/V2/V1/s1 [1]));
 OR2_X1 \V2/V2/V1/A1/M2/_0_  (.A1(\V2/V2/V1/A1/M2/c1 ),
    .A2(\V2/V2/V1/A1/M2/c2 ),
    .ZN(\V2/V2/V1/A1/c2 ));
 AND2_X1 \V2/V2/V1/A1/M3/M1/_0_  (.A1(\V2/V2/V1/v2 [2]),
    .A2(\V2/V2/V1/v3 [2]),
    .ZN(\V2/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M3/M1/_1_  (.A(\V2/V2/V1/v2 [2]),
    .B(\V2/V2/V1/v3 [2]),
    .Z(\V2/V2/V1/A1/M3/s1 ));
 AND2_X1 \V2/V2/V1/A1/M3/M2/_0_  (.A1(\V2/V2/V1/A1/M3/s1 ),
    .A2(\V2/V2/V1/A1/c2 ),
    .ZN(\V2/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M3/M2/_1_  (.A(\V2/V2/V1/A1/M3/s1 ),
    .B(\V2/V2/V1/A1/c2 ),
    .Z(\V2/V2/V1/s1 [2]));
 OR2_X1 \V2/V2/V1/A1/M3/_0_  (.A1(\V2/V2/V1/A1/M3/c1 ),
    .A2(\V2/V2/V1/A1/M3/c2 ),
    .ZN(\V2/V2/V1/A1/c3 ));
 AND2_X1 \V2/V2/V1/A1/M4/M1/_0_  (.A1(\V2/V2/V1/v2 [3]),
    .A2(\V2/V2/V1/v3 [3]),
    .ZN(\V2/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A1/M4/M1/_1_  (.A(\V2/V2/V1/v2 [3]),
    .B(\V2/V2/V1/v3 [3]),
    .Z(\V2/V2/V1/A1/M4/s1 ));
 AND2_X1 \V2/V2/V1/A1/M4/M2/_0_  (.A1(\V2/V2/V1/A1/M4/s1 ),
    .A2(\V2/V2/V1/A1/c3 ),
    .ZN(\V2/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A1/M4/M2/_1_  (.A(\V2/V2/V1/A1/M4/s1 ),
    .B(\V2/V2/V1/A1/c3 ),
    .Z(\V2/V2/V1/s1 [3]));
 OR2_X1 \V2/V2/V1/A1/M4/_0_  (.A1(\V2/V2/V1/A1/M4/c1 ),
    .A2(\V2/V2/V1/A1/M4/c2 ),
    .ZN(\V2/V2/V1/c1 ));
 AND2_X1 \V2/V2/V1/A2/M1/M1/_0_  (.A1(\V2/V2/V1/s1 [0]),
    .A2(\V2/V2/V1/v1 [2]),
    .ZN(\V2/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M1/M1/_1_  (.A(\V2/V2/V1/s1 [0]),
    .B(\V2/V2/V1/v1 [2]),
    .Z(\V2/V2/V1/A2/M1/s1 ));
 AND2_X1 \V2/V2/V1/A2/M1/M2/_0_  (.A1(\V2/V2/V1/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M1/M2/_1_  (.A(\V2/V2/V1/A2/M1/s1 ),
    .B(net2),
    .Z(\V2/v2 [2]));
 OR2_X1 \V2/V2/V1/A2/M1/_0_  (.A1(\V2/V2/V1/A2/M1/c1 ),
    .A2(\V2/V2/V1/A2/M1/c2 ),
    .ZN(\V2/V2/V1/A2/c1 ));
 AND2_X1 \V2/V2/V1/A2/M2/M1/_0_  (.A1(\V2/V2/V1/s1 [1]),
    .A2(\V2/V2/V1/v1 [3]),
    .ZN(\V2/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M2/M1/_1_  (.A(\V2/V2/V1/s1 [1]),
    .B(\V2/V2/V1/v1 [3]),
    .Z(\V2/V2/V1/A2/M2/s1 ));
 AND2_X1 \V2/V2/V1/A2/M2/M2/_0_  (.A1(\V2/V2/V1/A2/M2/s1 ),
    .A2(\V2/V2/V1/A2/c1 ),
    .ZN(\V2/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M2/M2/_1_  (.A(\V2/V2/V1/A2/M2/s1 ),
    .B(\V2/V2/V1/A2/c1 ),
    .Z(\V2/v2 [3]));
 OR2_X1 \V2/V2/V1/A2/M2/_0_  (.A1(\V2/V2/V1/A2/M2/c1 ),
    .A2(\V2/V2/V1/A2/M2/c2 ),
    .ZN(\V2/V2/V1/A2/c2 ));
 AND2_X1 \V2/V2/V1/A2/M3/M1/_0_  (.A1(\V2/V2/V1/s1 [2]),
    .A2(net2),
    .ZN(\V2/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M3/M1/_1_  (.A(\V2/V2/V1/s1 [2]),
    .B(net2),
    .Z(\V2/V2/V1/A2/M3/s1 ));
 AND2_X1 \V2/V2/V1/A2/M3/M2/_0_  (.A1(\V2/V2/V1/A2/M3/s1 ),
    .A2(\V2/V2/V1/A2/c2 ),
    .ZN(\V2/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M3/M2/_1_  (.A(\V2/V2/V1/A2/M3/s1 ),
    .B(\V2/V2/V1/A2/c2 ),
    .Z(\V2/V2/V1/s2 [2]));
 OR2_X1 \V2/V2/V1/A2/M3/_0_  (.A1(\V2/V2/V1/A2/M3/c1 ),
    .A2(\V2/V2/V1/A2/M3/c2 ),
    .ZN(\V2/V2/V1/A2/c3 ));
 AND2_X1 \V2/V2/V1/A2/M4/M1/_0_  (.A1(\V2/V2/V1/s1 [3]),
    .A2(net2),
    .ZN(\V2/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A2/M4/M1/_1_  (.A(\V2/V2/V1/s1 [3]),
    .B(net2),
    .Z(\V2/V2/V1/A2/M4/s1 ));
 AND2_X1 \V2/V2/V1/A2/M4/M2/_0_  (.A1(\V2/V2/V1/A2/M4/s1 ),
    .A2(\V2/V2/V1/A2/c3 ),
    .ZN(\V2/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A2/M4/M2/_1_  (.A(\V2/V2/V1/A2/M4/s1 ),
    .B(\V2/V2/V1/A2/c3 ),
    .Z(\V2/V2/V1/s2 [3]));
 OR2_X1 \V2/V2/V1/A2/M4/_0_  (.A1(\V2/V2/V1/A2/M4/c1 ),
    .A2(\V2/V2/V1/A2/M4/c2 ),
    .ZN(\V2/V2/V1/c2 ));
 AND2_X1 \V2/V2/V1/A3/M1/M1/_0_  (.A1(\V2/V2/V1/v4 [0]),
    .A2(\V2/V2/V1/s2 [2]),
    .ZN(\V2/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M1/M1/_1_  (.A(\V2/V2/V1/v4 [0]),
    .B(\V2/V2/V1/s2 [2]),
    .Z(\V2/V2/V1/A3/M1/s1 ));
 AND2_X1 \V2/V2/V1/A3/M1/M2/_0_  (.A1(\V2/V2/V1/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M1/M2/_1_  (.A(\V2/V2/V1/A3/M1/s1 ),
    .B(net2),
    .Z(\V2/V2/v1 [4]));
 OR2_X1 \V2/V2/V1/A3/M1/_0_  (.A1(\V2/V2/V1/A3/M1/c1 ),
    .A2(\V2/V2/V1/A3/M1/c2 ),
    .ZN(\V2/V2/V1/A3/c1 ));
 AND2_X1 \V2/V2/V1/A3/M2/M1/_0_  (.A1(\V2/V2/V1/v4 [1]),
    .A2(\V2/V2/V1/s2 [3]),
    .ZN(\V2/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M2/M1/_1_  (.A(\V2/V2/V1/v4 [1]),
    .B(\V2/V2/V1/s2 [3]),
    .Z(\V2/V2/V1/A3/M2/s1 ));
 AND2_X1 \V2/V2/V1/A3/M2/M2/_0_  (.A1(\V2/V2/V1/A3/M2/s1 ),
    .A2(\V2/V2/V1/A3/c1 ),
    .ZN(\V2/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M2/M2/_1_  (.A(\V2/V2/V1/A3/M2/s1 ),
    .B(\V2/V2/V1/A3/c1 ),
    .Z(\V2/V2/v1 [5]));
 OR2_X1 \V2/V2/V1/A3/M2/_0_  (.A1(\V2/V2/V1/A3/M2/c1 ),
    .A2(\V2/V2/V1/A3/M2/c2 ),
    .ZN(\V2/V2/V1/A3/c2 ));
 AND2_X1 \V2/V2/V1/A3/M3/M1/_0_  (.A1(\V2/V2/V1/v4 [2]),
    .A2(\V2/V2/V1/c3 ),
    .ZN(\V2/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M3/M1/_1_  (.A(\V2/V2/V1/v4 [2]),
    .B(\V2/V2/V1/c3 ),
    .Z(\V2/V2/V1/A3/M3/s1 ));
 AND2_X1 \V2/V2/V1/A3/M3/M2/_0_  (.A1(\V2/V2/V1/A3/M3/s1 ),
    .A2(\V2/V2/V1/A3/c2 ),
    .ZN(\V2/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M3/M2/_1_  (.A(\V2/V2/V1/A3/M3/s1 ),
    .B(\V2/V2/V1/A3/c2 ),
    .Z(\V2/V2/v1 [6]));
 OR2_X1 \V2/V2/V1/A3/M3/_0_  (.A1(\V2/V2/V1/A3/M3/c1 ),
    .A2(\V2/V2/V1/A3/M3/c2 ),
    .ZN(\V2/V2/V1/A3/c3 ));
 AND2_X1 \V2/V2/V1/A3/M4/M1/_0_  (.A1(\V2/V2/V1/v4 [3]),
    .A2(net2),
    .ZN(\V2/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V1/A3/M4/M1/_1_  (.A(\V2/V2/V1/v4 [3]),
    .B(net2),
    .Z(\V2/V2/V1/A3/M4/s1 ));
 AND2_X1 \V2/V2/V1/A3/M4/M2/_0_  (.A1(\V2/V2/V1/A3/M4/s1 ),
    .A2(\V2/V2/V1/A3/c3 ),
    .ZN(\V2/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V1/A3/M4/M2/_1_  (.A(\V2/V2/V1/A3/M4/s1 ),
    .B(\V2/V2/V1/A3/c3 ),
    .Z(\V2/V2/v1 [7]));
 OR2_X1 \V2/V2/V1/A3/M4/_0_  (.A1(\V2/V2/V1/A3/M4/c1 ),
    .A2(\V2/V2/V1/A3/M4/c2 ),
    .ZN(\V2/V2/V1/overflow ));
 AND2_X1 \V2/V2/V1/V1/HA1/_0_  (.A1(\V2/V2/V1/V1/w2 ),
    .A2(\V2/V2/V1/V1/w1 ),
    .ZN(\V2/V2/V1/V1/w4 ));
 XOR2_X2 \V2/V2/V1/V1/HA1/_1_  (.A(\V2/V2/V1/V1/w2 ),
    .B(\V2/V2/V1/V1/w1 ),
    .Z(\V2/v2 [1]));
 AND2_X1 \V2/V2/V1/V1/HA2/_0_  (.A1(\V2/V2/V1/V1/w4 ),
    .A2(\V2/V2/V1/V1/w3 ),
    .ZN(\V2/V2/V1/v1 [3]));
 XOR2_X2 \V2/V2/V1/V1/HA2/_1_  (.A(\V2/V2/V1/V1/w4 ),
    .B(\V2/V2/V1/V1/w3 ),
    .Z(\V2/V2/V1/v1 [2]));
 AND2_X1 \V2/V2/V1/V1/_0_  (.A1(net33),
    .A2(net23),
    .ZN(\V2/v2 [0]));
 AND2_X1 \V2/V2/V1/V1/_1_  (.A1(net33),
    .A2(B[1]),
    .ZN(\V2/V2/V1/V1/w1 ));
 AND2_X1 \V2/V2/V1/V1/_2_  (.A1(net23),
    .A2(net32),
    .ZN(\V2/V2/V1/V1/w2 ));
 AND2_X1 \V2/V2/V1/V1/_3_  (.A1(B[1]),
    .A2(net32),
    .ZN(\V2/V2/V1/V1/w3 ));
 AND2_X1 \V2/V2/V1/V2/HA1/_0_  (.A1(\V2/V2/V1/V2/w2 ),
    .A2(\V2/V2/V1/V2/w1 ),
    .ZN(\V2/V2/V1/V2/w4 ));
 XOR2_X2 \V2/V2/V1/V2/HA1/_1_  (.A(\V2/V2/V1/V2/w2 ),
    .B(\V2/V2/V1/V2/w1 ),
    .Z(\V2/V2/V1/v2 [1]));
 AND2_X1 \V2/V2/V1/V2/HA2/_0_  (.A1(\V2/V2/V1/V2/w4 ),
    .A2(\V2/V2/V1/V2/w3 ),
    .ZN(\V2/V2/V1/v2 [3]));
 XOR2_X2 \V2/V2/V1/V2/HA2/_1_  (.A(\V2/V2/V1/V2/w4 ),
    .B(\V2/V2/V1/V2/w3 ),
    .Z(\V2/V2/V1/v2 [2]));
 AND2_X1 \V2/V2/V1/V2/_0_  (.A1(net31),
    .A2(net23),
    .ZN(\V2/V2/V1/v2 [0]));
 AND2_X1 \V2/V2/V1/V2/_1_  (.A1(net31),
    .A2(B[1]),
    .ZN(\V2/V2/V1/V2/w1 ));
 AND2_X1 \V2/V2/V1/V2/_2_  (.A1(net23),
    .A2(net30),
    .ZN(\V2/V2/V1/V2/w2 ));
 AND2_X1 \V2/V2/V1/V2/_3_  (.A1(B[1]),
    .A2(net30),
    .ZN(\V2/V2/V1/V2/w3 ));
 AND2_X1 \V2/V2/V1/V3/HA1/_0_  (.A1(\V2/V2/V1/V3/w2 ),
    .A2(\V2/V2/V1/V3/w1 ),
    .ZN(\V2/V2/V1/V3/w4 ));
 XOR2_X2 \V2/V2/V1/V3/HA1/_1_  (.A(\V2/V2/V1/V3/w2 ),
    .B(\V2/V2/V1/V3/w1 ),
    .Z(\V2/V2/V1/v3 [1]));
 AND2_X1 \V2/V2/V1/V3/HA2/_0_  (.A1(\V2/V2/V1/V3/w4 ),
    .A2(\V2/V2/V1/V3/w3 ),
    .ZN(\V2/V2/V1/v3 [3]));
 XOR2_X2 \V2/V2/V1/V3/HA2/_1_  (.A(\V2/V2/V1/V3/w4 ),
    .B(\V2/V2/V1/V3/w3 ),
    .Z(\V2/V2/V1/v3 [2]));
 AND2_X1 \V2/V2/V1/V3/_0_  (.A1(net33),
    .A2(B[2]),
    .ZN(\V2/V2/V1/v3 [0]));
 AND2_X1 \V2/V2/V1/V3/_1_  (.A1(net33),
    .A2(B[3]),
    .ZN(\V2/V2/V1/V3/w1 ));
 AND2_X1 \V2/V2/V1/V3/_2_  (.A1(B[2]),
    .A2(net32),
    .ZN(\V2/V2/V1/V3/w2 ));
 AND2_X1 \V2/V2/V1/V3/_3_  (.A1(B[3]),
    .A2(net32),
    .ZN(\V2/V2/V1/V3/w3 ));
 AND2_X1 \V2/V2/V1/V4/HA1/_0_  (.A1(\V2/V2/V1/V4/w2 ),
    .A2(\V2/V2/V1/V4/w1 ),
    .ZN(\V2/V2/V1/V4/w4 ));
 XOR2_X2 \V2/V2/V1/V4/HA1/_1_  (.A(\V2/V2/V1/V4/w2 ),
    .B(\V2/V2/V1/V4/w1 ),
    .Z(\V2/V2/V1/v4 [1]));
 AND2_X1 \V2/V2/V1/V4/HA2/_0_  (.A1(\V2/V2/V1/V4/w4 ),
    .A2(\V2/V2/V1/V4/w3 ),
    .ZN(\V2/V2/V1/v4 [3]));
 XOR2_X2 \V2/V2/V1/V4/HA2/_1_  (.A(\V2/V2/V1/V4/w4 ),
    .B(\V2/V2/V1/V4/w3 ),
    .Z(\V2/V2/V1/v4 [2]));
 AND2_X1 \V2/V2/V1/V4/_0_  (.A1(net31),
    .A2(B[2]),
    .ZN(\V2/V2/V1/v4 [0]));
 AND2_X1 \V2/V2/V1/V4/_1_  (.A1(net31),
    .A2(B[3]),
    .ZN(\V2/V2/V1/V4/w1 ));
 AND2_X1 \V2/V2/V1/V4/_2_  (.A1(B[2]),
    .A2(net30),
    .ZN(\V2/V2/V1/V4/w2 ));
 AND2_X1 \V2/V2/V1/V4/_3_  (.A1(B[3]),
    .A2(net30),
    .ZN(\V2/V2/V1/V4/w3 ));
 OR2_X1 \V2/V2/V1/_0_  (.A1(\V2/V2/V1/c1 ),
    .A2(\V2/V2/V1/c2 ),
    .ZN(\V2/V2/V1/c3 ));
 AND2_X1 \V2/V2/V2/A1/M1/M1/_0_  (.A1(\V2/V2/V2/v2 [0]),
    .A2(\V2/V2/V2/v3 [0]),
    .ZN(\V2/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M1/M1/_1_  (.A(\V2/V2/V2/v2 [0]),
    .B(\V2/V2/V2/v3 [0]),
    .Z(\V2/V2/V2/A1/M1/s1 ));
 AND2_X1 \V2/V2/V2/A1/M1/M2/_0_  (.A1(\V2/V2/V2/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M1/M2/_1_  (.A(\V2/V2/V2/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/V2/s1 [0]));
 OR2_X1 \V2/V2/V2/A1/M1/_0_  (.A1(\V2/V2/V2/A1/M1/c1 ),
    .A2(\V2/V2/V2/A1/M1/c2 ),
    .ZN(\V2/V2/V2/A1/c1 ));
 AND2_X1 \V2/V2/V2/A1/M2/M1/_0_  (.A1(\V2/V2/V2/v2 [1]),
    .A2(\V2/V2/V2/v3 [1]),
    .ZN(\V2/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M2/M1/_1_  (.A(\V2/V2/V2/v2 [1]),
    .B(\V2/V2/V2/v3 [1]),
    .Z(\V2/V2/V2/A1/M2/s1 ));
 AND2_X1 \V2/V2/V2/A1/M2/M2/_0_  (.A1(\V2/V2/V2/A1/M2/s1 ),
    .A2(\V2/V2/V2/A1/c1 ),
    .ZN(\V2/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M2/M2/_1_  (.A(\V2/V2/V2/A1/M2/s1 ),
    .B(\V2/V2/V2/A1/c1 ),
    .Z(\V2/V2/V2/s1 [1]));
 OR2_X1 \V2/V2/V2/A1/M2/_0_  (.A1(\V2/V2/V2/A1/M2/c1 ),
    .A2(\V2/V2/V2/A1/M2/c2 ),
    .ZN(\V2/V2/V2/A1/c2 ));
 AND2_X1 \V2/V2/V2/A1/M3/M1/_0_  (.A1(\V2/V2/V2/v2 [2]),
    .A2(\V2/V2/V2/v3 [2]),
    .ZN(\V2/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M3/M1/_1_  (.A(\V2/V2/V2/v2 [2]),
    .B(\V2/V2/V2/v3 [2]),
    .Z(\V2/V2/V2/A1/M3/s1 ));
 AND2_X1 \V2/V2/V2/A1/M3/M2/_0_  (.A1(\V2/V2/V2/A1/M3/s1 ),
    .A2(\V2/V2/V2/A1/c2 ),
    .ZN(\V2/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M3/M2/_1_  (.A(\V2/V2/V2/A1/M3/s1 ),
    .B(\V2/V2/V2/A1/c2 ),
    .Z(\V2/V2/V2/s1 [2]));
 OR2_X1 \V2/V2/V2/A1/M3/_0_  (.A1(\V2/V2/V2/A1/M3/c1 ),
    .A2(\V2/V2/V2/A1/M3/c2 ),
    .ZN(\V2/V2/V2/A1/c3 ));
 AND2_X1 \V2/V2/V2/A1/M4/M1/_0_  (.A1(\V2/V2/V2/v2 [3]),
    .A2(\V2/V2/V2/v3 [3]),
    .ZN(\V2/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A1/M4/M1/_1_  (.A(\V2/V2/V2/v2 [3]),
    .B(\V2/V2/V2/v3 [3]),
    .Z(\V2/V2/V2/A1/M4/s1 ));
 AND2_X1 \V2/V2/V2/A1/M4/M2/_0_  (.A1(\V2/V2/V2/A1/M4/s1 ),
    .A2(\V2/V2/V2/A1/c3 ),
    .ZN(\V2/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A1/M4/M2/_1_  (.A(\V2/V2/V2/A1/M4/s1 ),
    .B(\V2/V2/V2/A1/c3 ),
    .Z(\V2/V2/V2/s1 [3]));
 OR2_X1 \V2/V2/V2/A1/M4/_0_  (.A1(\V2/V2/V2/A1/M4/c1 ),
    .A2(\V2/V2/V2/A1/M4/c2 ),
    .ZN(\V2/V2/V2/c1 ));
 AND2_X1 \V2/V2/V2/A2/M1/M1/_0_  (.A1(\V2/V2/V2/s1 [0]),
    .A2(\V2/V2/V2/v1 [2]),
    .ZN(\V2/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M1/M1/_1_  (.A(\V2/V2/V2/s1 [0]),
    .B(\V2/V2/V2/v1 [2]),
    .Z(\V2/V2/V2/A2/M1/s1 ));
 AND2_X1 \V2/V2/V2/A2/M1/M2/_0_  (.A1(\V2/V2/V2/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M1/M2/_1_  (.A(\V2/V2/V2/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/v2 [2]));
 OR2_X1 \V2/V2/V2/A2/M1/_0_  (.A1(\V2/V2/V2/A2/M1/c1 ),
    .A2(\V2/V2/V2/A2/M1/c2 ),
    .ZN(\V2/V2/V2/A2/c1 ));
 AND2_X1 \V2/V2/V2/A2/M2/M1/_0_  (.A1(\V2/V2/V2/s1 [1]),
    .A2(\V2/V2/V2/v1 [3]),
    .ZN(\V2/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M2/M1/_1_  (.A(\V2/V2/V2/s1 [1]),
    .B(\V2/V2/V2/v1 [3]),
    .Z(\V2/V2/V2/A2/M2/s1 ));
 AND2_X1 \V2/V2/V2/A2/M2/M2/_0_  (.A1(\V2/V2/V2/A2/M2/s1 ),
    .A2(\V2/V2/V2/A2/c1 ),
    .ZN(\V2/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M2/M2/_1_  (.A(\V2/V2/V2/A2/M2/s1 ),
    .B(\V2/V2/V2/A2/c1 ),
    .Z(\V2/V2/v2 [3]));
 OR2_X1 \V2/V2/V2/A2/M2/_0_  (.A1(\V2/V2/V2/A2/M2/c1 ),
    .A2(\V2/V2/V2/A2/M2/c2 ),
    .ZN(\V2/V2/V2/A2/c2 ));
 AND2_X1 \V2/V2/V2/A2/M3/M1/_0_  (.A1(\V2/V2/V2/s1 [2]),
    .A2(net9),
    .ZN(\V2/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M3/M1/_1_  (.A(\V2/V2/V2/s1 [2]),
    .B(net9),
    .Z(\V2/V2/V2/A2/M3/s1 ));
 AND2_X1 \V2/V2/V2/A2/M3/M2/_0_  (.A1(\V2/V2/V2/A2/M3/s1 ),
    .A2(\V2/V2/V2/A2/c2 ),
    .ZN(\V2/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M3/M2/_1_  (.A(\V2/V2/V2/A2/M3/s1 ),
    .B(\V2/V2/V2/A2/c2 ),
    .Z(\V2/V2/V2/s2 [2]));
 OR2_X1 \V2/V2/V2/A2/M3/_0_  (.A1(\V2/V2/V2/A2/M3/c1 ),
    .A2(\V2/V2/V2/A2/M3/c2 ),
    .ZN(\V2/V2/V2/A2/c3 ));
 AND2_X1 \V2/V2/V2/A2/M4/M1/_0_  (.A1(\V2/V2/V2/s1 [3]),
    .A2(net9),
    .ZN(\V2/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A2/M4/M1/_1_  (.A(\V2/V2/V2/s1 [3]),
    .B(net9),
    .Z(\V2/V2/V2/A2/M4/s1 ));
 AND2_X1 \V2/V2/V2/A2/M4/M2/_0_  (.A1(\V2/V2/V2/A2/M4/s1 ),
    .A2(\V2/V2/V2/A2/c3 ),
    .ZN(\V2/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A2/M4/M2/_1_  (.A(\V2/V2/V2/A2/M4/s1 ),
    .B(\V2/V2/V2/A2/c3 ),
    .Z(\V2/V2/V2/s2 [3]));
 OR2_X1 \V2/V2/V2/A2/M4/_0_  (.A1(\V2/V2/V2/A2/M4/c1 ),
    .A2(\V2/V2/V2/A2/M4/c2 ),
    .ZN(\V2/V2/V2/c2 ));
 AND2_X1 \V2/V2/V2/A3/M1/M1/_0_  (.A1(\V2/V2/V2/v4 [0]),
    .A2(\V2/V2/V2/s2 [2]),
    .ZN(\V2/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M1/M1/_1_  (.A(\V2/V2/V2/v4 [0]),
    .B(\V2/V2/V2/s2 [2]),
    .Z(\V2/V2/V2/A3/M1/s1 ));
 AND2_X1 \V2/V2/V2/A3/M1/M2/_0_  (.A1(\V2/V2/V2/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M1/M2/_1_  (.A(\V2/V2/V2/A3/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/v2 [4]));
 OR2_X1 \V2/V2/V2/A3/M1/_0_  (.A1(\V2/V2/V2/A3/M1/c1 ),
    .A2(\V2/V2/V2/A3/M1/c2 ),
    .ZN(\V2/V2/V2/A3/c1 ));
 AND2_X1 \V2/V2/V2/A3/M2/M1/_0_  (.A1(\V2/V2/V2/v4 [1]),
    .A2(\V2/V2/V2/s2 [3]),
    .ZN(\V2/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M2/M1/_1_  (.A(\V2/V2/V2/v4 [1]),
    .B(\V2/V2/V2/s2 [3]),
    .Z(\V2/V2/V2/A3/M2/s1 ));
 AND2_X1 \V2/V2/V2/A3/M2/M2/_0_  (.A1(\V2/V2/V2/A3/M2/s1 ),
    .A2(\V2/V2/V2/A3/c1 ),
    .ZN(\V2/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M2/M2/_1_  (.A(\V2/V2/V2/A3/M2/s1 ),
    .B(\V2/V2/V2/A3/c1 ),
    .Z(\V2/V2/v2 [5]));
 OR2_X1 \V2/V2/V2/A3/M2/_0_  (.A1(\V2/V2/V2/A3/M2/c1 ),
    .A2(\V2/V2/V2/A3/M2/c2 ),
    .ZN(\V2/V2/V2/A3/c2 ));
 AND2_X1 \V2/V2/V2/A3/M3/M1/_0_  (.A1(\V2/V2/V2/v4 [2]),
    .A2(\V2/V2/V2/c3 ),
    .ZN(\V2/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M3/M1/_1_  (.A(\V2/V2/V2/v4 [2]),
    .B(\V2/V2/V2/c3 ),
    .Z(\V2/V2/V2/A3/M3/s1 ));
 AND2_X1 \V2/V2/V2/A3/M3/M2/_0_  (.A1(\V2/V2/V2/A3/M3/s1 ),
    .A2(\V2/V2/V2/A3/c2 ),
    .ZN(\V2/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M3/M2/_1_  (.A(\V2/V2/V2/A3/M3/s1 ),
    .B(\V2/V2/V2/A3/c2 ),
    .Z(\V2/V2/v2 [6]));
 OR2_X1 \V2/V2/V2/A3/M3/_0_  (.A1(\V2/V2/V2/A3/M3/c1 ),
    .A2(\V2/V2/V2/A3/M3/c2 ),
    .ZN(\V2/V2/V2/A3/c3 ));
 AND2_X1 \V2/V2/V2/A3/M4/M1/_0_  (.A1(\V2/V2/V2/v4 [3]),
    .A2(net9),
    .ZN(\V2/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V2/A3/M4/M1/_1_  (.A(\V2/V2/V2/v4 [3]),
    .B(net9),
    .Z(\V2/V2/V2/A3/M4/s1 ));
 AND2_X1 \V2/V2/V2/A3/M4/M2/_0_  (.A1(\V2/V2/V2/A3/M4/s1 ),
    .A2(\V2/V2/V2/A3/c3 ),
    .ZN(\V2/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V2/A3/M4/M2/_1_  (.A(\V2/V2/V2/A3/M4/s1 ),
    .B(\V2/V2/V2/A3/c3 ),
    .Z(\V2/V2/v2 [7]));
 OR2_X1 \V2/V2/V2/A3/M4/_0_  (.A1(\V2/V2/V2/A3/M4/c1 ),
    .A2(\V2/V2/V2/A3/M4/c2 ),
    .ZN(\V2/V2/V2/overflow ));
 AND2_X1 \V2/V2/V2/V1/HA1/_0_  (.A1(\V2/V2/V2/V1/w2 ),
    .A2(\V2/V2/V2/V1/w1 ),
    .ZN(\V2/V2/V2/V1/w4 ));
 XOR2_X2 \V2/V2/V2/V1/HA1/_1_  (.A(\V2/V2/V2/V1/w2 ),
    .B(\V2/V2/V2/V1/w1 ),
    .Z(\V2/V2/v2 [1]));
 AND2_X1 \V2/V2/V2/V1/HA2/_0_  (.A1(\V2/V2/V2/V1/w4 ),
    .A2(\V2/V2/V2/V1/w3 ),
    .ZN(\V2/V2/V2/v1 [3]));
 XOR2_X2 \V2/V2/V2/V1/HA2/_1_  (.A(\V2/V2/V2/V1/w4 ),
    .B(\V2/V2/V2/V1/w3 ),
    .Z(\V2/V2/V2/v1 [2]));
 AND2_X1 \V2/V2/V2/V1/_0_  (.A1(net29),
    .A2(net23),
    .ZN(\V2/V2/v2 [0]));
 AND2_X1 \V2/V2/V2/V1/_1_  (.A1(net29),
    .A2(B[1]),
    .ZN(\V2/V2/V2/V1/w1 ));
 AND2_X1 \V2/V2/V2/V1/_2_  (.A1(net23),
    .A2(net28),
    .ZN(\V2/V2/V2/V1/w2 ));
 AND2_X1 \V2/V2/V2/V1/_3_  (.A1(B[1]),
    .A2(net28),
    .ZN(\V2/V2/V2/V1/w3 ));
 AND2_X1 \V2/V2/V2/V2/HA1/_0_  (.A1(\V2/V2/V2/V2/w2 ),
    .A2(\V2/V2/V2/V2/w1 ),
    .ZN(\V2/V2/V2/V2/w4 ));
 XOR2_X2 \V2/V2/V2/V2/HA1/_1_  (.A(\V2/V2/V2/V2/w2 ),
    .B(\V2/V2/V2/V2/w1 ),
    .Z(\V2/V2/V2/v2 [1]));
 AND2_X1 \V2/V2/V2/V2/HA2/_0_  (.A1(\V2/V2/V2/V2/w4 ),
    .A2(\V2/V2/V2/V2/w3 ),
    .ZN(\V2/V2/V2/v2 [3]));
 XOR2_X2 \V2/V2/V2/V2/HA2/_1_  (.A(\V2/V2/V2/V2/w4 ),
    .B(\V2/V2/V2/V2/w3 ),
    .Z(\V2/V2/V2/v2 [2]));
 AND2_X1 \V2/V2/V2/V2/_0_  (.A1(net27),
    .A2(net23),
    .ZN(\V2/V2/V2/v2 [0]));
 AND2_X1 \V2/V2/V2/V2/_1_  (.A1(net27),
    .A2(B[1]),
    .ZN(\V2/V2/V2/V2/w1 ));
 AND2_X1 \V2/V2/V2/V2/_2_  (.A1(net23),
    .A2(net26),
    .ZN(\V2/V2/V2/V2/w2 ));
 AND2_X1 \V2/V2/V2/V2/_3_  (.A1(B[1]),
    .A2(net26),
    .ZN(\V2/V2/V2/V2/w3 ));
 AND2_X1 \V2/V2/V2/V3/HA1/_0_  (.A1(\V2/V2/V2/V3/w2 ),
    .A2(\V2/V2/V2/V3/w1 ),
    .ZN(\V2/V2/V2/V3/w4 ));
 XOR2_X2 \V2/V2/V2/V3/HA1/_1_  (.A(\V2/V2/V2/V3/w2 ),
    .B(\V2/V2/V2/V3/w1 ),
    .Z(\V2/V2/V2/v3 [1]));
 AND2_X1 \V2/V2/V2/V3/HA2/_0_  (.A1(\V2/V2/V2/V3/w4 ),
    .A2(\V2/V2/V2/V3/w3 ),
    .ZN(\V2/V2/V2/v3 [3]));
 XOR2_X2 \V2/V2/V2/V3/HA2/_1_  (.A(\V2/V2/V2/V3/w4 ),
    .B(\V2/V2/V2/V3/w3 ),
    .Z(\V2/V2/V2/v3 [2]));
 AND2_X1 \V2/V2/V2/V3/_0_  (.A1(net29),
    .A2(B[2]),
    .ZN(\V2/V2/V2/v3 [0]));
 AND2_X1 \V2/V2/V2/V3/_1_  (.A1(net29),
    .A2(B[3]),
    .ZN(\V2/V2/V2/V3/w1 ));
 AND2_X1 \V2/V2/V2/V3/_2_  (.A1(B[2]),
    .A2(net28),
    .ZN(\V2/V2/V2/V3/w2 ));
 AND2_X1 \V2/V2/V2/V3/_3_  (.A1(B[3]),
    .A2(net28),
    .ZN(\V2/V2/V2/V3/w3 ));
 AND2_X1 \V2/V2/V2/V4/HA1/_0_  (.A1(\V2/V2/V2/V4/w2 ),
    .A2(\V2/V2/V2/V4/w1 ),
    .ZN(\V2/V2/V2/V4/w4 ));
 XOR2_X2 \V2/V2/V2/V4/HA1/_1_  (.A(\V2/V2/V2/V4/w2 ),
    .B(\V2/V2/V2/V4/w1 ),
    .Z(\V2/V2/V2/v4 [1]));
 AND2_X1 \V2/V2/V2/V4/HA2/_0_  (.A1(\V2/V2/V2/V4/w4 ),
    .A2(\V2/V2/V2/V4/w3 ),
    .ZN(\V2/V2/V2/v4 [3]));
 XOR2_X2 \V2/V2/V2/V4/HA2/_1_  (.A(\V2/V2/V2/V4/w4 ),
    .B(\V2/V2/V2/V4/w3 ),
    .Z(\V2/V2/V2/v4 [2]));
 AND2_X1 \V2/V2/V2/V4/_0_  (.A1(net27),
    .A2(B[2]),
    .ZN(\V2/V2/V2/v4 [0]));
 AND2_X1 \V2/V2/V2/V4/_1_  (.A1(net27),
    .A2(B[3]),
    .ZN(\V2/V2/V2/V4/w1 ));
 AND2_X1 \V2/V2/V2/V4/_2_  (.A1(B[2]),
    .A2(net26),
    .ZN(\V2/V2/V2/V4/w2 ));
 AND2_X1 \V2/V2/V2/V4/_3_  (.A1(B[3]),
    .A2(net26),
    .ZN(\V2/V2/V2/V4/w3 ));
 OR2_X1 \V2/V2/V2/_0_  (.A1(\V2/V2/V2/c1 ),
    .A2(\V2/V2/V2/c2 ),
    .ZN(\V2/V2/V2/c3 ));
 AND2_X1 \V2/V2/V3/A1/M1/M1/_0_  (.A1(\V2/V2/V3/v2 [0]),
    .A2(\V2/V2/V3/v3 [0]),
    .ZN(\V2/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M1/M1/_1_  (.A(\V2/V2/V3/v2 [0]),
    .B(\V2/V2/V3/v3 [0]),
    .Z(\V2/V2/V3/A1/M1/s1 ));
 AND2_X1 \V2/V2/V3/A1/M1/M2/_0_  (.A1(\V2/V2/V3/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M1/M2/_1_  (.A(\V2/V2/V3/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/V3/s1 [0]));
 OR2_X1 \V2/V2/V3/A1/M1/_0_  (.A1(\V2/V2/V3/A1/M1/c1 ),
    .A2(\V2/V2/V3/A1/M1/c2 ),
    .ZN(\V2/V2/V3/A1/c1 ));
 AND2_X1 \V2/V2/V3/A1/M2/M1/_0_  (.A1(\V2/V2/V3/v2 [1]),
    .A2(\V2/V2/V3/v3 [1]),
    .ZN(\V2/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M2/M1/_1_  (.A(\V2/V2/V3/v2 [1]),
    .B(\V2/V2/V3/v3 [1]),
    .Z(\V2/V2/V3/A1/M2/s1 ));
 AND2_X1 \V2/V2/V3/A1/M2/M2/_0_  (.A1(\V2/V2/V3/A1/M2/s1 ),
    .A2(\V2/V2/V3/A1/c1 ),
    .ZN(\V2/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M2/M2/_1_  (.A(\V2/V2/V3/A1/M2/s1 ),
    .B(\V2/V2/V3/A1/c1 ),
    .Z(\V2/V2/V3/s1 [1]));
 OR2_X1 \V2/V2/V3/A1/M2/_0_  (.A1(\V2/V2/V3/A1/M2/c1 ),
    .A2(\V2/V2/V3/A1/M2/c2 ),
    .ZN(\V2/V2/V3/A1/c2 ));
 AND2_X1 \V2/V2/V3/A1/M3/M1/_0_  (.A1(\V2/V2/V3/v2 [2]),
    .A2(\V2/V2/V3/v3 [2]),
    .ZN(\V2/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M3/M1/_1_  (.A(\V2/V2/V3/v2 [2]),
    .B(\V2/V2/V3/v3 [2]),
    .Z(\V2/V2/V3/A1/M3/s1 ));
 AND2_X1 \V2/V2/V3/A1/M3/M2/_0_  (.A1(\V2/V2/V3/A1/M3/s1 ),
    .A2(\V2/V2/V3/A1/c2 ),
    .ZN(\V2/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M3/M2/_1_  (.A(\V2/V2/V3/A1/M3/s1 ),
    .B(\V2/V2/V3/A1/c2 ),
    .Z(\V2/V2/V3/s1 [2]));
 OR2_X1 \V2/V2/V3/A1/M3/_0_  (.A1(\V2/V2/V3/A1/M3/c1 ),
    .A2(\V2/V2/V3/A1/M3/c2 ),
    .ZN(\V2/V2/V3/A1/c3 ));
 AND2_X1 \V2/V2/V3/A1/M4/M1/_0_  (.A1(\V2/V2/V3/v2 [3]),
    .A2(\V2/V2/V3/v3 [3]),
    .ZN(\V2/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A1/M4/M1/_1_  (.A(\V2/V2/V3/v2 [3]),
    .B(\V2/V2/V3/v3 [3]),
    .Z(\V2/V2/V3/A1/M4/s1 ));
 AND2_X1 \V2/V2/V3/A1/M4/M2/_0_  (.A1(\V2/V2/V3/A1/M4/s1 ),
    .A2(\V2/V2/V3/A1/c3 ),
    .ZN(\V2/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A1/M4/M2/_1_  (.A(\V2/V2/V3/A1/M4/s1 ),
    .B(\V2/V2/V3/A1/c3 ),
    .Z(\V2/V2/V3/s1 [3]));
 OR2_X1 \V2/V2/V3/A1/M4/_0_  (.A1(\V2/V2/V3/A1/M4/c1 ),
    .A2(\V2/V2/V3/A1/M4/c2 ),
    .ZN(\V2/V2/V3/c1 ));
 AND2_X1 \V2/V2/V3/A2/M1/M1/_0_  (.A1(\V2/V2/V3/s1 [0]),
    .A2(\V2/V2/V3/v1 [2]),
    .ZN(\V2/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M1/M1/_1_  (.A(\V2/V2/V3/s1 [0]),
    .B(\V2/V2/V3/v1 [2]),
    .Z(\V2/V2/V3/A2/M1/s1 ));
 AND2_X1 \V2/V2/V3/A2/M1/M2/_0_  (.A1(\V2/V2/V3/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M1/M2/_1_  (.A(\V2/V2/V3/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/v3 [2]));
 OR2_X1 \V2/V2/V3/A2/M1/_0_  (.A1(\V2/V2/V3/A2/M1/c1 ),
    .A2(\V2/V2/V3/A2/M1/c2 ),
    .ZN(\V2/V2/V3/A2/c1 ));
 AND2_X1 \V2/V2/V3/A2/M2/M1/_0_  (.A1(\V2/V2/V3/s1 [1]),
    .A2(\V2/V2/V3/v1 [3]),
    .ZN(\V2/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M2/M1/_1_  (.A(\V2/V2/V3/s1 [1]),
    .B(\V2/V2/V3/v1 [3]),
    .Z(\V2/V2/V3/A2/M2/s1 ));
 AND2_X1 \V2/V2/V3/A2/M2/M2/_0_  (.A1(\V2/V2/V3/A2/M2/s1 ),
    .A2(\V2/V2/V3/A2/c1 ),
    .ZN(\V2/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M2/M2/_1_  (.A(\V2/V2/V3/A2/M2/s1 ),
    .B(\V2/V2/V3/A2/c1 ),
    .Z(\V2/V2/v3 [3]));
 OR2_X1 \V2/V2/V3/A2/M2/_0_  (.A1(\V2/V2/V3/A2/M2/c1 ),
    .A2(\V2/V2/V3/A2/M2/c2 ),
    .ZN(\V2/V2/V3/A2/c2 ));
 AND2_X1 \V2/V2/V3/A2/M3/M1/_0_  (.A1(\V2/V2/V3/s1 [2]),
    .A2(net7),
    .ZN(\V2/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M3/M1/_1_  (.A(\V2/V2/V3/s1 [2]),
    .B(net7),
    .Z(\V2/V2/V3/A2/M3/s1 ));
 AND2_X1 \V2/V2/V3/A2/M3/M2/_0_  (.A1(\V2/V2/V3/A2/M3/s1 ),
    .A2(\V2/V2/V3/A2/c2 ),
    .ZN(\V2/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M3/M2/_1_  (.A(\V2/V2/V3/A2/M3/s1 ),
    .B(\V2/V2/V3/A2/c2 ),
    .Z(\V2/V2/V3/s2 [2]));
 OR2_X1 \V2/V2/V3/A2/M3/_0_  (.A1(\V2/V2/V3/A2/M3/c1 ),
    .A2(\V2/V2/V3/A2/M3/c2 ),
    .ZN(\V2/V2/V3/A2/c3 ));
 AND2_X1 \V2/V2/V3/A2/M4/M1/_0_  (.A1(\V2/V2/V3/s1 [3]),
    .A2(net7),
    .ZN(\V2/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A2/M4/M1/_1_  (.A(\V2/V2/V3/s1 [3]),
    .B(net7),
    .Z(\V2/V2/V3/A2/M4/s1 ));
 AND2_X1 \V2/V2/V3/A2/M4/M2/_0_  (.A1(\V2/V2/V3/A2/M4/s1 ),
    .A2(\V2/V2/V3/A2/c3 ),
    .ZN(\V2/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A2/M4/M2/_1_  (.A(\V2/V2/V3/A2/M4/s1 ),
    .B(\V2/V2/V3/A2/c3 ),
    .Z(\V2/V2/V3/s2 [3]));
 OR2_X1 \V2/V2/V3/A2/M4/_0_  (.A1(\V2/V2/V3/A2/M4/c1 ),
    .A2(\V2/V2/V3/A2/M4/c2 ),
    .ZN(\V2/V2/V3/c2 ));
 AND2_X1 \V2/V2/V3/A3/M1/M1/_0_  (.A1(\V2/V2/V3/v4 [0]),
    .A2(\V2/V2/V3/s2 [2]),
    .ZN(\V2/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M1/M1/_1_  (.A(\V2/V2/V3/v4 [0]),
    .B(\V2/V2/V3/s2 [2]),
    .Z(\V2/V2/V3/A3/M1/s1 ));
 AND2_X1 \V2/V2/V3/A3/M1/M2/_0_  (.A1(\V2/V2/V3/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M1/M2/_1_  (.A(\V2/V2/V3/A3/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/v3 [4]));
 OR2_X1 \V2/V2/V3/A3/M1/_0_  (.A1(\V2/V2/V3/A3/M1/c1 ),
    .A2(\V2/V2/V3/A3/M1/c2 ),
    .ZN(\V2/V2/V3/A3/c1 ));
 AND2_X1 \V2/V2/V3/A3/M2/M1/_0_  (.A1(\V2/V2/V3/v4 [1]),
    .A2(\V2/V2/V3/s2 [3]),
    .ZN(\V2/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M2/M1/_1_  (.A(\V2/V2/V3/v4 [1]),
    .B(\V2/V2/V3/s2 [3]),
    .Z(\V2/V2/V3/A3/M2/s1 ));
 AND2_X1 \V2/V2/V3/A3/M2/M2/_0_  (.A1(\V2/V2/V3/A3/M2/s1 ),
    .A2(\V2/V2/V3/A3/c1 ),
    .ZN(\V2/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M2/M2/_1_  (.A(\V2/V2/V3/A3/M2/s1 ),
    .B(\V2/V2/V3/A3/c1 ),
    .Z(\V2/V2/v3 [5]));
 OR2_X1 \V2/V2/V3/A3/M2/_0_  (.A1(\V2/V2/V3/A3/M2/c1 ),
    .A2(\V2/V2/V3/A3/M2/c2 ),
    .ZN(\V2/V2/V3/A3/c2 ));
 AND2_X1 \V2/V2/V3/A3/M3/M1/_0_  (.A1(\V2/V2/V3/v4 [2]),
    .A2(\V2/V2/V3/c3 ),
    .ZN(\V2/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M3/M1/_1_  (.A(\V2/V2/V3/v4 [2]),
    .B(\V2/V2/V3/c3 ),
    .Z(\V2/V2/V3/A3/M3/s1 ));
 AND2_X1 \V2/V2/V3/A3/M3/M2/_0_  (.A1(\V2/V2/V3/A3/M3/s1 ),
    .A2(\V2/V2/V3/A3/c2 ),
    .ZN(\V2/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M3/M2/_1_  (.A(\V2/V2/V3/A3/M3/s1 ),
    .B(\V2/V2/V3/A3/c2 ),
    .Z(\V2/V2/v3 [6]));
 OR2_X1 \V2/V2/V3/A3/M3/_0_  (.A1(\V2/V2/V3/A3/M3/c1 ),
    .A2(\V2/V2/V3/A3/M3/c2 ),
    .ZN(\V2/V2/V3/A3/c3 ));
 AND2_X1 \V2/V2/V3/A3/M4/M1/_0_  (.A1(\V2/V2/V3/v4 [3]),
    .A2(net7),
    .ZN(\V2/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V3/A3/M4/M1/_1_  (.A(\V2/V2/V3/v4 [3]),
    .B(net7),
    .Z(\V2/V2/V3/A3/M4/s1 ));
 AND2_X1 \V2/V2/V3/A3/M4/M2/_0_  (.A1(\V2/V2/V3/A3/M4/s1 ),
    .A2(\V2/V2/V3/A3/c3 ),
    .ZN(\V2/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V3/A3/M4/M2/_1_  (.A(\V2/V2/V3/A3/M4/s1 ),
    .B(\V2/V2/V3/A3/c3 ),
    .Z(\V2/V2/v3 [7]));
 OR2_X1 \V2/V2/V3/A3/M4/_0_  (.A1(\V2/V2/V3/A3/M4/c1 ),
    .A2(\V2/V2/V3/A3/M4/c2 ),
    .ZN(\V2/V2/V3/overflow ));
 AND2_X1 \V2/V2/V3/V1/HA1/_0_  (.A1(\V2/V2/V3/V1/w2 ),
    .A2(\V2/V2/V3/V1/w1 ),
    .ZN(\V2/V2/V3/V1/w4 ));
 XOR2_X2 \V2/V2/V3/V1/HA1/_1_  (.A(\V2/V2/V3/V1/w2 ),
    .B(\V2/V2/V3/V1/w1 ),
    .Z(\V2/V2/v3 [1]));
 AND2_X1 \V2/V2/V3/V1/HA2/_0_  (.A1(\V2/V2/V3/V1/w4 ),
    .A2(\V2/V2/V3/V1/w3 ),
    .ZN(\V2/V2/V3/v1 [3]));
 XOR2_X2 \V2/V2/V3/V1/HA2/_1_  (.A(\V2/V2/V3/V1/w4 ),
    .B(\V2/V2/V3/V1/w3 ),
    .Z(\V2/V2/V3/v1 [2]));
 AND2_X1 \V2/V2/V3/V1/_0_  (.A1(net33),
    .A2(B[4]),
    .ZN(\V2/V2/v3 [0]));
 AND2_X1 \V2/V2/V3/V1/_1_  (.A1(net33),
    .A2(B[5]),
    .ZN(\V2/V2/V3/V1/w1 ));
 AND2_X1 \V2/V2/V3/V1/_2_  (.A1(B[4]),
    .A2(net32),
    .ZN(\V2/V2/V3/V1/w2 ));
 AND2_X1 \V2/V2/V3/V1/_3_  (.A1(B[5]),
    .A2(net32),
    .ZN(\V2/V2/V3/V1/w3 ));
 AND2_X1 \V2/V2/V3/V2/HA1/_0_  (.A1(\V2/V2/V3/V2/w2 ),
    .A2(\V2/V2/V3/V2/w1 ),
    .ZN(\V2/V2/V3/V2/w4 ));
 XOR2_X2 \V2/V2/V3/V2/HA1/_1_  (.A(\V2/V2/V3/V2/w2 ),
    .B(\V2/V2/V3/V2/w1 ),
    .Z(\V2/V2/V3/v2 [1]));
 AND2_X1 \V2/V2/V3/V2/HA2/_0_  (.A1(\V2/V2/V3/V2/w4 ),
    .A2(\V2/V2/V3/V2/w3 ),
    .ZN(\V2/V2/V3/v2 [3]));
 XOR2_X2 \V2/V2/V3/V2/HA2/_1_  (.A(\V2/V2/V3/V2/w4 ),
    .B(\V2/V2/V3/V2/w3 ),
    .Z(\V2/V2/V3/v2 [2]));
 AND2_X1 \V2/V2/V3/V2/_0_  (.A1(net31),
    .A2(B[4]),
    .ZN(\V2/V2/V3/v2 [0]));
 AND2_X1 \V2/V2/V3/V2/_1_  (.A1(net31),
    .A2(B[5]),
    .ZN(\V2/V2/V3/V2/w1 ));
 AND2_X1 \V2/V2/V3/V2/_2_  (.A1(B[4]),
    .A2(net30),
    .ZN(\V2/V2/V3/V2/w2 ));
 AND2_X1 \V2/V2/V3/V2/_3_  (.A1(B[5]),
    .A2(net30),
    .ZN(\V2/V2/V3/V2/w3 ));
 AND2_X1 \V2/V2/V3/V3/HA1/_0_  (.A1(\V2/V2/V3/V3/w2 ),
    .A2(\V2/V2/V3/V3/w1 ),
    .ZN(\V2/V2/V3/V3/w4 ));
 XOR2_X2 \V2/V2/V3/V3/HA1/_1_  (.A(\V2/V2/V3/V3/w2 ),
    .B(\V2/V2/V3/V3/w1 ),
    .Z(\V2/V2/V3/v3 [1]));
 AND2_X1 \V2/V2/V3/V3/HA2/_0_  (.A1(\V2/V2/V3/V3/w4 ),
    .A2(\V2/V2/V3/V3/w3 ),
    .ZN(\V2/V2/V3/v3 [3]));
 XOR2_X2 \V2/V2/V3/V3/HA2/_1_  (.A(\V2/V2/V3/V3/w4 ),
    .B(\V2/V2/V3/V3/w3 ),
    .Z(\V2/V2/V3/v3 [2]));
 AND2_X1 \V2/V2/V3/V3/_0_  (.A1(net33),
    .A2(B[6]),
    .ZN(\V2/V2/V3/v3 [0]));
 AND2_X1 \V2/V2/V3/V3/_1_  (.A1(net33),
    .A2(B[7]),
    .ZN(\V2/V2/V3/V3/w1 ));
 AND2_X1 \V2/V2/V3/V3/_2_  (.A1(B[6]),
    .A2(net32),
    .ZN(\V2/V2/V3/V3/w2 ));
 AND2_X1 \V2/V2/V3/V3/_3_  (.A1(B[7]),
    .A2(net32),
    .ZN(\V2/V2/V3/V3/w3 ));
 AND2_X1 \V2/V2/V3/V4/HA1/_0_  (.A1(\V2/V2/V3/V4/w2 ),
    .A2(\V2/V2/V3/V4/w1 ),
    .ZN(\V2/V2/V3/V4/w4 ));
 XOR2_X2 \V2/V2/V3/V4/HA1/_1_  (.A(\V2/V2/V3/V4/w2 ),
    .B(\V2/V2/V3/V4/w1 ),
    .Z(\V2/V2/V3/v4 [1]));
 AND2_X1 \V2/V2/V3/V4/HA2/_0_  (.A1(\V2/V2/V3/V4/w4 ),
    .A2(\V2/V2/V3/V4/w3 ),
    .ZN(\V2/V2/V3/v4 [3]));
 XOR2_X2 \V2/V2/V3/V4/HA2/_1_  (.A(\V2/V2/V3/V4/w4 ),
    .B(\V2/V2/V3/V4/w3 ),
    .Z(\V2/V2/V3/v4 [2]));
 AND2_X1 \V2/V2/V3/V4/_0_  (.A1(net31),
    .A2(B[6]),
    .ZN(\V2/V2/V3/v4 [0]));
 AND2_X1 \V2/V2/V3/V4/_1_  (.A1(net31),
    .A2(B[7]),
    .ZN(\V2/V2/V3/V4/w1 ));
 AND2_X1 \V2/V2/V3/V4/_2_  (.A1(B[6]),
    .A2(net30),
    .ZN(\V2/V2/V3/V4/w2 ));
 AND2_X1 \V2/V2/V3/V4/_3_  (.A1(B[7]),
    .A2(net30),
    .ZN(\V2/V2/V3/V4/w3 ));
 OR2_X1 \V2/V2/V3/_0_  (.A1(\V2/V2/V3/c1 ),
    .A2(\V2/V2/V3/c2 ),
    .ZN(\V2/V2/V3/c3 ));
 AND2_X1 \V2/V2/V4/A1/M1/M1/_0_  (.A1(\V2/V2/V4/v2 [0]),
    .A2(\V2/V2/V4/v3 [0]),
    .ZN(\V2/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M1/M1/_1_  (.A(\V2/V2/V4/v2 [0]),
    .B(\V2/V2/V4/v3 [0]),
    .Z(\V2/V2/V4/A1/M1/s1 ));
 AND2_X1 \V2/V2/V4/A1/M1/M2/_0_  (.A1(\V2/V2/V4/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M1/M2/_1_  (.A(\V2/V2/V4/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/V4/s1 [0]));
 OR2_X1 \V2/V2/V4/A1/M1/_0_  (.A1(\V2/V2/V4/A1/M1/c1 ),
    .A2(\V2/V2/V4/A1/M1/c2 ),
    .ZN(\V2/V2/V4/A1/c1 ));
 AND2_X1 \V2/V2/V4/A1/M2/M1/_0_  (.A1(\V2/V2/V4/v2 [1]),
    .A2(\V2/V2/V4/v3 [1]),
    .ZN(\V2/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M2/M1/_1_  (.A(\V2/V2/V4/v2 [1]),
    .B(\V2/V2/V4/v3 [1]),
    .Z(\V2/V2/V4/A1/M2/s1 ));
 AND2_X1 \V2/V2/V4/A1/M2/M2/_0_  (.A1(\V2/V2/V4/A1/M2/s1 ),
    .A2(\V2/V2/V4/A1/c1 ),
    .ZN(\V2/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M2/M2/_1_  (.A(\V2/V2/V4/A1/M2/s1 ),
    .B(\V2/V2/V4/A1/c1 ),
    .Z(\V2/V2/V4/s1 [1]));
 OR2_X1 \V2/V2/V4/A1/M2/_0_  (.A1(\V2/V2/V4/A1/M2/c1 ),
    .A2(\V2/V2/V4/A1/M2/c2 ),
    .ZN(\V2/V2/V4/A1/c2 ));
 AND2_X1 \V2/V2/V4/A1/M3/M1/_0_  (.A1(\V2/V2/V4/v2 [2]),
    .A2(\V2/V2/V4/v3 [2]),
    .ZN(\V2/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M3/M1/_1_  (.A(\V2/V2/V4/v2 [2]),
    .B(\V2/V2/V4/v3 [2]),
    .Z(\V2/V2/V4/A1/M3/s1 ));
 AND2_X1 \V2/V2/V4/A1/M3/M2/_0_  (.A1(\V2/V2/V4/A1/M3/s1 ),
    .A2(\V2/V2/V4/A1/c2 ),
    .ZN(\V2/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M3/M2/_1_  (.A(\V2/V2/V4/A1/M3/s1 ),
    .B(\V2/V2/V4/A1/c2 ),
    .Z(\V2/V2/V4/s1 [2]));
 OR2_X1 \V2/V2/V4/A1/M3/_0_  (.A1(\V2/V2/V4/A1/M3/c1 ),
    .A2(\V2/V2/V4/A1/M3/c2 ),
    .ZN(\V2/V2/V4/A1/c3 ));
 AND2_X1 \V2/V2/V4/A1/M4/M1/_0_  (.A1(\V2/V2/V4/v2 [3]),
    .A2(\V2/V2/V4/v3 [3]),
    .ZN(\V2/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A1/M4/M1/_1_  (.A(\V2/V2/V4/v2 [3]),
    .B(\V2/V2/V4/v3 [3]),
    .Z(\V2/V2/V4/A1/M4/s1 ));
 AND2_X1 \V2/V2/V4/A1/M4/M2/_0_  (.A1(\V2/V2/V4/A1/M4/s1 ),
    .A2(\V2/V2/V4/A1/c3 ),
    .ZN(\V2/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A1/M4/M2/_1_  (.A(\V2/V2/V4/A1/M4/s1 ),
    .B(\V2/V2/V4/A1/c3 ),
    .Z(\V2/V2/V4/s1 [3]));
 OR2_X1 \V2/V2/V4/A1/M4/_0_  (.A1(\V2/V2/V4/A1/M4/c1 ),
    .A2(\V2/V2/V4/A1/M4/c2 ),
    .ZN(\V2/V2/V4/c1 ));
 AND2_X1 \V2/V2/V4/A2/M1/M1/_0_  (.A1(\V2/V2/V4/s1 [0]),
    .A2(\V2/V2/V4/v1 [2]),
    .ZN(\V2/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M1/M1/_1_  (.A(\V2/V2/V4/s1 [0]),
    .B(\V2/V2/V4/v1 [2]),
    .Z(\V2/V2/V4/A2/M1/s1 ));
 AND2_X1 \V2/V2/V4/A2/M1/M2/_0_  (.A1(\V2/V2/V4/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M1/M2/_1_  (.A(\V2/V2/V4/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V2/v4 [2]));
 OR2_X1 \V2/V2/V4/A2/M1/_0_  (.A1(\V2/V2/V4/A2/M1/c1 ),
    .A2(\V2/V2/V4/A2/M1/c2 ),
    .ZN(\V2/V2/V4/A2/c1 ));
 AND2_X1 \V2/V2/V4/A2/M2/M1/_0_  (.A1(\V2/V2/V4/s1 [1]),
    .A2(\V2/V2/V4/v1 [3]),
    .ZN(\V2/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M2/M1/_1_  (.A(\V2/V2/V4/s1 [1]),
    .B(\V2/V2/V4/v1 [3]),
    .Z(\V2/V2/V4/A2/M2/s1 ));
 AND2_X1 \V2/V2/V4/A2/M2/M2/_0_  (.A1(\V2/V2/V4/A2/M2/s1 ),
    .A2(\V2/V2/V4/A2/c1 ),
    .ZN(\V2/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M2/M2/_1_  (.A(\V2/V2/V4/A2/M2/s1 ),
    .B(\V2/V2/V4/A2/c1 ),
    .Z(\V2/V2/v4 [3]));
 OR2_X1 \V2/V2/V4/A2/M2/_0_  (.A1(\V2/V2/V4/A2/M2/c1 ),
    .A2(\V2/V2/V4/A2/M2/c2 ),
    .ZN(\V2/V2/V4/A2/c2 ));
 AND2_X1 \V2/V2/V4/A2/M3/M1/_0_  (.A1(\V2/V2/V4/s1 [2]),
    .A2(net9),
    .ZN(\V2/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M3/M1/_1_  (.A(\V2/V2/V4/s1 [2]),
    .B(net9),
    .Z(\V2/V2/V4/A2/M3/s1 ));
 AND2_X1 \V2/V2/V4/A2/M3/M2/_0_  (.A1(\V2/V2/V4/A2/M3/s1 ),
    .A2(\V2/V2/V4/A2/c2 ),
    .ZN(\V2/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M3/M2/_1_  (.A(\V2/V2/V4/A2/M3/s1 ),
    .B(\V2/V2/V4/A2/c2 ),
    .Z(\V2/V2/V4/s2 [2]));
 OR2_X1 \V2/V2/V4/A2/M3/_0_  (.A1(\V2/V2/V4/A2/M3/c1 ),
    .A2(\V2/V2/V4/A2/M3/c2 ),
    .ZN(\V2/V2/V4/A2/c3 ));
 AND2_X1 \V2/V2/V4/A2/M4/M1/_0_  (.A1(\V2/V2/V4/s1 [3]),
    .A2(net9),
    .ZN(\V2/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A2/M4/M1/_1_  (.A(\V2/V2/V4/s1 [3]),
    .B(net9),
    .Z(\V2/V2/V4/A2/M4/s1 ));
 AND2_X1 \V2/V2/V4/A2/M4/M2/_0_  (.A1(\V2/V2/V4/A2/M4/s1 ),
    .A2(\V2/V2/V4/A2/c3 ),
    .ZN(\V2/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A2/M4/M2/_1_  (.A(\V2/V2/V4/A2/M4/s1 ),
    .B(\V2/V2/V4/A2/c3 ),
    .Z(\V2/V2/V4/s2 [3]));
 OR2_X1 \V2/V2/V4/A2/M4/_0_  (.A1(\V2/V2/V4/A2/M4/c1 ),
    .A2(\V2/V2/V4/A2/M4/c2 ),
    .ZN(\V2/V2/V4/c2 ));
 AND2_X1 \V2/V2/V4/A3/M1/M1/_0_  (.A1(\V2/V2/V4/v4 [0]),
    .A2(\V2/V2/V4/s2 [2]),
    .ZN(\V2/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M1/M1/_1_  (.A(\V2/V2/V4/v4 [0]),
    .B(\V2/V2/V4/s2 [2]),
    .Z(\V2/V2/V4/A3/M1/s1 ));
 AND2_X1 \V2/V2/V4/A3/M1/M2/_0_  (.A1(\V2/V2/V4/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M1/M2/_1_  (.A(\V2/V2/V4/A3/M1/s1 ),
    .B(net9),
    .Z(\V2/V2/v4 [4]));
 OR2_X1 \V2/V2/V4/A3/M1/_0_  (.A1(\V2/V2/V4/A3/M1/c1 ),
    .A2(\V2/V2/V4/A3/M1/c2 ),
    .ZN(\V2/V2/V4/A3/c1 ));
 AND2_X1 \V2/V2/V4/A3/M2/M1/_0_  (.A1(\V2/V2/V4/v4 [1]),
    .A2(\V2/V2/V4/s2 [3]),
    .ZN(\V2/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M2/M1/_1_  (.A(\V2/V2/V4/v4 [1]),
    .B(\V2/V2/V4/s2 [3]),
    .Z(\V2/V2/V4/A3/M2/s1 ));
 AND2_X1 \V2/V2/V4/A3/M2/M2/_0_  (.A1(\V2/V2/V4/A3/M2/s1 ),
    .A2(\V2/V2/V4/A3/c1 ),
    .ZN(\V2/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M2/M2/_1_  (.A(\V2/V2/V4/A3/M2/s1 ),
    .B(\V2/V2/V4/A3/c1 ),
    .Z(\V2/V2/v4 [5]));
 OR2_X1 \V2/V2/V4/A3/M2/_0_  (.A1(\V2/V2/V4/A3/M2/c1 ),
    .A2(\V2/V2/V4/A3/M2/c2 ),
    .ZN(\V2/V2/V4/A3/c2 ));
 AND2_X1 \V2/V2/V4/A3/M3/M1/_0_  (.A1(\V2/V2/V4/v4 [2]),
    .A2(\V2/V2/V4/c3 ),
    .ZN(\V2/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M3/M1/_1_  (.A(\V2/V2/V4/v4 [2]),
    .B(\V2/V2/V4/c3 ),
    .Z(\V2/V2/V4/A3/M3/s1 ));
 AND2_X1 \V2/V2/V4/A3/M3/M2/_0_  (.A1(\V2/V2/V4/A3/M3/s1 ),
    .A2(\V2/V2/V4/A3/c2 ),
    .ZN(\V2/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M3/M2/_1_  (.A(\V2/V2/V4/A3/M3/s1 ),
    .B(\V2/V2/V4/A3/c2 ),
    .Z(\V2/V2/v4 [6]));
 OR2_X1 \V2/V2/V4/A3/M3/_0_  (.A1(\V2/V2/V4/A3/M3/c1 ),
    .A2(\V2/V2/V4/A3/M3/c2 ),
    .ZN(\V2/V2/V4/A3/c3 ));
 AND2_X1 \V2/V2/V4/A3/M4/M1/_0_  (.A1(\V2/V2/V4/v4 [3]),
    .A2(net9),
    .ZN(\V2/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V2/V4/A3/M4/M1/_1_  (.A(\V2/V2/V4/v4 [3]),
    .B(net9),
    .Z(\V2/V2/V4/A3/M4/s1 ));
 AND2_X1 \V2/V2/V4/A3/M4/M2/_0_  (.A1(\V2/V2/V4/A3/M4/s1 ),
    .A2(\V2/V2/V4/A3/c3 ),
    .ZN(\V2/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V2/V4/A3/M4/M2/_1_  (.A(\V2/V2/V4/A3/M4/s1 ),
    .B(\V2/V2/V4/A3/c3 ),
    .Z(\V2/V2/v4 [7]));
 OR2_X1 \V2/V2/V4/A3/M4/_0_  (.A1(\V2/V2/V4/A3/M4/c1 ),
    .A2(\V2/V2/V4/A3/M4/c2 ),
    .ZN(\V2/V2/V4/overflow ));
 AND2_X1 \V2/V2/V4/V1/HA1/_0_  (.A1(\V2/V2/V4/V1/w2 ),
    .A2(\V2/V2/V4/V1/w1 ),
    .ZN(\V2/V2/V4/V1/w4 ));
 XOR2_X2 \V2/V2/V4/V1/HA1/_1_  (.A(\V2/V2/V4/V1/w2 ),
    .B(\V2/V2/V4/V1/w1 ),
    .Z(\V2/V2/v4 [1]));
 AND2_X1 \V2/V2/V4/V1/HA2/_0_  (.A1(\V2/V2/V4/V1/w4 ),
    .A2(\V2/V2/V4/V1/w3 ),
    .ZN(\V2/V2/V4/v1 [3]));
 XOR2_X2 \V2/V2/V4/V1/HA2/_1_  (.A(\V2/V2/V4/V1/w4 ),
    .B(\V2/V2/V4/V1/w3 ),
    .Z(\V2/V2/V4/v1 [2]));
 AND2_X1 \V2/V2/V4/V1/_0_  (.A1(net29),
    .A2(B[4]),
    .ZN(\V2/V2/v4 [0]));
 AND2_X1 \V2/V2/V4/V1/_1_  (.A1(net29),
    .A2(B[5]),
    .ZN(\V2/V2/V4/V1/w1 ));
 AND2_X1 \V2/V2/V4/V1/_2_  (.A1(B[4]),
    .A2(net28),
    .ZN(\V2/V2/V4/V1/w2 ));
 AND2_X1 \V2/V2/V4/V1/_3_  (.A1(B[5]),
    .A2(net28),
    .ZN(\V2/V2/V4/V1/w3 ));
 AND2_X1 \V2/V2/V4/V2/HA1/_0_  (.A1(\V2/V2/V4/V2/w2 ),
    .A2(\V2/V2/V4/V2/w1 ),
    .ZN(\V2/V2/V4/V2/w4 ));
 XOR2_X2 \V2/V2/V4/V2/HA1/_1_  (.A(\V2/V2/V4/V2/w2 ),
    .B(\V2/V2/V4/V2/w1 ),
    .Z(\V2/V2/V4/v2 [1]));
 AND2_X1 \V2/V2/V4/V2/HA2/_0_  (.A1(\V2/V2/V4/V2/w4 ),
    .A2(\V2/V2/V4/V2/w3 ),
    .ZN(\V2/V2/V4/v2 [3]));
 XOR2_X2 \V2/V2/V4/V2/HA2/_1_  (.A(\V2/V2/V4/V2/w4 ),
    .B(\V2/V2/V4/V2/w3 ),
    .Z(\V2/V2/V4/v2 [2]));
 AND2_X1 \V2/V2/V4/V2/_0_  (.A1(net27),
    .A2(B[4]),
    .ZN(\V2/V2/V4/v2 [0]));
 AND2_X1 \V2/V2/V4/V2/_1_  (.A1(net27),
    .A2(B[5]),
    .ZN(\V2/V2/V4/V2/w1 ));
 AND2_X1 \V2/V2/V4/V2/_2_  (.A1(B[4]),
    .A2(net26),
    .ZN(\V2/V2/V4/V2/w2 ));
 AND2_X1 \V2/V2/V4/V2/_3_  (.A1(B[5]),
    .A2(net26),
    .ZN(\V2/V2/V4/V2/w3 ));
 AND2_X1 \V2/V2/V4/V3/HA1/_0_  (.A1(\V2/V2/V4/V3/w2 ),
    .A2(\V2/V2/V4/V3/w1 ),
    .ZN(\V2/V2/V4/V3/w4 ));
 XOR2_X2 \V2/V2/V4/V3/HA1/_1_  (.A(\V2/V2/V4/V3/w2 ),
    .B(\V2/V2/V4/V3/w1 ),
    .Z(\V2/V2/V4/v3 [1]));
 AND2_X1 \V2/V2/V4/V3/HA2/_0_  (.A1(\V2/V2/V4/V3/w4 ),
    .A2(\V2/V2/V4/V3/w3 ),
    .ZN(\V2/V2/V4/v3 [3]));
 XOR2_X2 \V2/V2/V4/V3/HA2/_1_  (.A(\V2/V2/V4/V3/w4 ),
    .B(\V2/V2/V4/V3/w3 ),
    .Z(\V2/V2/V4/v3 [2]));
 AND2_X1 \V2/V2/V4/V3/_0_  (.A1(net29),
    .A2(B[6]),
    .ZN(\V2/V2/V4/v3 [0]));
 AND2_X1 \V2/V2/V4/V3/_1_  (.A1(net29),
    .A2(B[7]),
    .ZN(\V2/V2/V4/V3/w1 ));
 AND2_X1 \V2/V2/V4/V3/_2_  (.A1(B[6]),
    .A2(net28),
    .ZN(\V2/V2/V4/V3/w2 ));
 AND2_X1 \V2/V2/V4/V3/_3_  (.A1(B[7]),
    .A2(net28),
    .ZN(\V2/V2/V4/V3/w3 ));
 AND2_X1 \V2/V2/V4/V4/HA1/_0_  (.A1(\V2/V2/V4/V4/w2 ),
    .A2(\V2/V2/V4/V4/w1 ),
    .ZN(\V2/V2/V4/V4/w4 ));
 XOR2_X2 \V2/V2/V4/V4/HA1/_1_  (.A(\V2/V2/V4/V4/w2 ),
    .B(\V2/V2/V4/V4/w1 ),
    .Z(\V2/V2/V4/v4 [1]));
 AND2_X1 \V2/V2/V4/V4/HA2/_0_  (.A1(\V2/V2/V4/V4/w4 ),
    .A2(\V2/V2/V4/V4/w3 ),
    .ZN(\V2/V2/V4/v4 [3]));
 XOR2_X2 \V2/V2/V4/V4/HA2/_1_  (.A(\V2/V2/V4/V4/w4 ),
    .B(\V2/V2/V4/V4/w3 ),
    .Z(\V2/V2/V4/v4 [2]));
 AND2_X1 \V2/V2/V4/V4/_0_  (.A1(net27),
    .A2(B[6]),
    .ZN(\V2/V2/V4/v4 [0]));
 AND2_X1 \V2/V2/V4/V4/_1_  (.A1(net27),
    .A2(B[7]),
    .ZN(\V2/V2/V4/V4/w1 ));
 AND2_X1 \V2/V2/V4/V4/_2_  (.A1(B[6]),
    .A2(net26),
    .ZN(\V2/V2/V4/V4/w2 ));
 AND2_X1 \V2/V2/V4/V4/_3_  (.A1(B[7]),
    .A2(net26),
    .ZN(\V2/V2/V4/V4/w3 ));
 OR2_X1 \V2/V2/V4/_0_  (.A1(\V2/V2/V4/c1 ),
    .A2(\V2/V2/V4/c2 ),
    .ZN(\V2/V2/V4/c3 ));
 OR2_X1 \V2/V2/_0_  (.A1(\V2/V2/c1 ),
    .A2(\V2/V2/c2 ),
    .ZN(\V2/V2/c3 ));
 AND2_X1 \V2/V3/A1/A1/M1/M1/_0_  (.A1(\V2/V3/v2 [0]),
    .A2(\V2/V3/v3 [0]),
    .ZN(\V2/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M1/M1/_1_  (.A(\V2/V3/v2 [0]),
    .B(\V2/V3/v3 [0]),
    .Z(\V2/V3/A1/A1/M1/s1 ));
 AND2_X1 \V2/V3/A1/A1/M1/M2/_0_  (.A1(\V2/V3/A1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M1/M2/_1_  (.A(\V2/V3/A1/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/V3/s1 [0]));
 OR2_X1 \V2/V3/A1/A1/M1/_0_  (.A1(\V2/V3/A1/A1/M1/c1 ),
    .A2(\V2/V3/A1/A1/M1/c2 ),
    .ZN(\V2/V3/A1/A1/c1 ));
 AND2_X1 \V2/V3/A1/A1/M2/M1/_0_  (.A1(\V2/V3/v2 [1]),
    .A2(\V2/V3/v3 [1]),
    .ZN(\V2/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M2/M1/_1_  (.A(\V2/V3/v2 [1]),
    .B(\V2/V3/v3 [1]),
    .Z(\V2/V3/A1/A1/M2/s1 ));
 AND2_X1 \V2/V3/A1/A1/M2/M2/_0_  (.A1(\V2/V3/A1/A1/M2/s1 ),
    .A2(\V2/V3/A1/A1/c1 ),
    .ZN(\V2/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M2/M2/_1_  (.A(\V2/V3/A1/A1/M2/s1 ),
    .B(\V2/V3/A1/A1/c1 ),
    .Z(\V2/V3/s1 [1]));
 OR2_X1 \V2/V3/A1/A1/M2/_0_  (.A1(\V2/V3/A1/A1/M2/c1 ),
    .A2(\V2/V3/A1/A1/M2/c2 ),
    .ZN(\V2/V3/A1/A1/c2 ));
 AND2_X1 \V2/V3/A1/A1/M3/M1/_0_  (.A1(\V2/V3/v2 [2]),
    .A2(\V2/V3/v3 [2]),
    .ZN(\V2/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M3/M1/_1_  (.A(\V2/V3/v2 [2]),
    .B(\V2/V3/v3 [2]),
    .Z(\V2/V3/A1/A1/M3/s1 ));
 AND2_X1 \V2/V3/A1/A1/M3/M2/_0_  (.A1(\V2/V3/A1/A1/M3/s1 ),
    .A2(\V2/V3/A1/A1/c2 ),
    .ZN(\V2/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M3/M2/_1_  (.A(\V2/V3/A1/A1/M3/s1 ),
    .B(\V2/V3/A1/A1/c2 ),
    .Z(\V2/V3/s1 [2]));
 OR2_X1 \V2/V3/A1/A1/M3/_0_  (.A1(\V2/V3/A1/A1/M3/c1 ),
    .A2(\V2/V3/A1/A1/M3/c2 ),
    .ZN(\V2/V3/A1/A1/c3 ));
 AND2_X1 \V2/V3/A1/A1/M4/M1/_0_  (.A1(\V2/V3/v2 [3]),
    .A2(\V2/V3/v3 [3]),
    .ZN(\V2/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A1/A1/M4/M1/_1_  (.A(\V2/V3/v2 [3]),
    .B(\V2/V3/v3 [3]),
    .Z(\V2/V3/A1/A1/M4/s1 ));
 AND2_X1 \V2/V3/A1/A1/M4/M2/_0_  (.A1(\V2/V3/A1/A1/M4/s1 ),
    .A2(\V2/V3/A1/A1/c3 ),
    .ZN(\V2/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A1/A1/M4/M2/_1_  (.A(\V2/V3/A1/A1/M4/s1 ),
    .B(\V2/V3/A1/A1/c3 ),
    .Z(\V2/V3/s1 [3]));
 OR2_X1 \V2/V3/A1/A1/M4/_0_  (.A1(\V2/V3/A1/A1/M4/c1 ),
    .A2(\V2/V3/A1/A1/M4/c2 ),
    .ZN(\V2/V3/A1/c1 ));
 AND2_X1 \V2/V3/A1/A2/M1/M1/_0_  (.A1(\V2/V3/v2 [4]),
    .A2(\V2/V3/v3 [4]),
    .ZN(\V2/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M1/M1/_1_  (.A(\V2/V3/v2 [4]),
    .B(\V2/V3/v3 [4]),
    .Z(\V2/V3/A1/A2/M1/s1 ));
 AND2_X1 \V2/V3/A1/A2/M1/M2/_0_  (.A1(\V2/V3/A1/A2/M1/s1 ),
    .A2(\V2/V3/A1/c1 ),
    .ZN(\V2/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M1/M2/_1_  (.A(\V2/V3/A1/A2/M1/s1 ),
    .B(\V2/V3/A1/c1 ),
    .Z(\V2/V3/s1 [4]));
 OR2_X1 \V2/V3/A1/A2/M1/_0_  (.A1(\V2/V3/A1/A2/M1/c1 ),
    .A2(\V2/V3/A1/A2/M1/c2 ),
    .ZN(\V2/V3/A1/A2/c1 ));
 AND2_X1 \V2/V3/A1/A2/M2/M1/_0_  (.A1(\V2/V3/v2 [5]),
    .A2(\V2/V3/v3 [5]),
    .ZN(\V2/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M2/M1/_1_  (.A(\V2/V3/v2 [5]),
    .B(\V2/V3/v3 [5]),
    .Z(\V2/V3/A1/A2/M2/s1 ));
 AND2_X1 \V2/V3/A1/A2/M2/M2/_0_  (.A1(\V2/V3/A1/A2/M2/s1 ),
    .A2(\V2/V3/A1/A2/c1 ),
    .ZN(\V2/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M2/M2/_1_  (.A(\V2/V3/A1/A2/M2/s1 ),
    .B(\V2/V3/A1/A2/c1 ),
    .Z(\V2/V3/s1 [5]));
 OR2_X1 \V2/V3/A1/A2/M2/_0_  (.A1(\V2/V3/A1/A2/M2/c1 ),
    .A2(\V2/V3/A1/A2/M2/c2 ),
    .ZN(\V2/V3/A1/A2/c2 ));
 AND2_X1 \V2/V3/A1/A2/M3/M1/_0_  (.A1(\V2/V3/v2 [6]),
    .A2(\V2/V3/v3 [6]),
    .ZN(\V2/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M3/M1/_1_  (.A(\V2/V3/v2 [6]),
    .B(\V2/V3/v3 [6]),
    .Z(\V2/V3/A1/A2/M3/s1 ));
 AND2_X1 \V2/V3/A1/A2/M3/M2/_0_  (.A1(\V2/V3/A1/A2/M3/s1 ),
    .A2(\V2/V3/A1/A2/c2 ),
    .ZN(\V2/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M3/M2/_1_  (.A(\V2/V3/A1/A2/M3/s1 ),
    .B(\V2/V3/A1/A2/c2 ),
    .Z(\V2/V3/s1 [6]));
 OR2_X1 \V2/V3/A1/A2/M3/_0_  (.A1(\V2/V3/A1/A2/M3/c1 ),
    .A2(\V2/V3/A1/A2/M3/c2 ),
    .ZN(\V2/V3/A1/A2/c3 ));
 AND2_X1 \V2/V3/A1/A2/M4/M1/_0_  (.A1(\V2/V3/v2 [7]),
    .A2(\V2/V3/v3 [7]),
    .ZN(\V2/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A1/A2/M4/M1/_1_  (.A(\V2/V3/v2 [7]),
    .B(\V2/V3/v3 [7]),
    .Z(\V2/V3/A1/A2/M4/s1 ));
 AND2_X1 \V2/V3/A1/A2/M4/M2/_0_  (.A1(\V2/V3/A1/A2/M4/s1 ),
    .A2(\V2/V3/A1/A2/c3 ),
    .ZN(\V2/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A1/A2/M4/M2/_1_  (.A(\V2/V3/A1/A2/M4/s1 ),
    .B(\V2/V3/A1/A2/c3 ),
    .Z(\V2/V3/s1 [7]));
 OR2_X1 \V2/V3/A1/A2/M4/_0_  (.A1(\V2/V3/A1/A2/M4/c1 ),
    .A2(\V2/V3/A1/A2/M4/c2 ),
    .ZN(\V2/V3/c1 ));
 AND2_X1 \V2/V3/A2/A1/M1/M1/_0_  (.A1(\V2/V3/s1 [0]),
    .A2(\V2/V3/v1 [4]),
    .ZN(\V2/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M1/M1/_1_  (.A(\V2/V3/s1 [0]),
    .B(\V2/V3/v1 [4]),
    .Z(\V2/V3/A2/A1/M1/s1 ));
 AND2_X1 \V2/V3/A2/A1/M1/M2/_0_  (.A1(\V2/V3/A2/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M1/M2/_1_  (.A(\V2/V3/A2/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/v3 [4]));
 OR2_X1 \V2/V3/A2/A1/M1/_0_  (.A1(\V2/V3/A2/A1/M1/c1 ),
    .A2(\V2/V3/A2/A1/M1/c2 ),
    .ZN(\V2/V3/A2/A1/c1 ));
 AND2_X1 \V2/V3/A2/A1/M2/M1/_0_  (.A1(\V2/V3/s1 [1]),
    .A2(\V2/V3/v1 [5]),
    .ZN(\V2/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M2/M1/_1_  (.A(\V2/V3/s1 [1]),
    .B(\V2/V3/v1 [5]),
    .Z(\V2/V3/A2/A1/M2/s1 ));
 AND2_X1 \V2/V3/A2/A1/M2/M2/_0_  (.A1(\V2/V3/A2/A1/M2/s1 ),
    .A2(\V2/V3/A2/A1/c1 ),
    .ZN(\V2/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M2/M2/_1_  (.A(\V2/V3/A2/A1/M2/s1 ),
    .B(\V2/V3/A2/A1/c1 ),
    .Z(\V2/v3 [5]));
 OR2_X1 \V2/V3/A2/A1/M2/_0_  (.A1(\V2/V3/A2/A1/M2/c1 ),
    .A2(\V2/V3/A2/A1/M2/c2 ),
    .ZN(\V2/V3/A2/A1/c2 ));
 AND2_X1 \V2/V3/A2/A1/M3/M1/_0_  (.A1(\V2/V3/s1 [2]),
    .A2(\V2/V3/v1 [6]),
    .ZN(\V2/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M3/M1/_1_  (.A(\V2/V3/s1 [2]),
    .B(\V2/V3/v1 [6]),
    .Z(\V2/V3/A2/A1/M3/s1 ));
 AND2_X1 \V2/V3/A2/A1/M3/M2/_0_  (.A1(\V2/V3/A2/A1/M3/s1 ),
    .A2(\V2/V3/A2/A1/c2 ),
    .ZN(\V2/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M3/M2/_1_  (.A(\V2/V3/A2/A1/M3/s1 ),
    .B(\V2/V3/A2/A1/c2 ),
    .Z(\V2/v3 [6]));
 OR2_X1 \V2/V3/A2/A1/M3/_0_  (.A1(\V2/V3/A2/A1/M3/c1 ),
    .A2(\V2/V3/A2/A1/M3/c2 ),
    .ZN(\V2/V3/A2/A1/c3 ));
 AND2_X1 \V2/V3/A2/A1/M4/M1/_0_  (.A1(\V2/V3/s1 [3]),
    .A2(\V2/V3/v1 [7]),
    .ZN(\V2/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A2/A1/M4/M1/_1_  (.A(\V2/V3/s1 [3]),
    .B(\V2/V3/v1 [7]),
    .Z(\V2/V3/A2/A1/M4/s1 ));
 AND2_X1 \V2/V3/A2/A1/M4/M2/_0_  (.A1(\V2/V3/A2/A1/M4/s1 ),
    .A2(\V2/V3/A2/A1/c3 ),
    .ZN(\V2/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A2/A1/M4/M2/_1_  (.A(\V2/V3/A2/A1/M4/s1 ),
    .B(\V2/V3/A2/A1/c3 ),
    .Z(\V2/v3 [7]));
 OR2_X1 \V2/V3/A2/A1/M4/_0_  (.A1(\V2/V3/A2/A1/M4/c1 ),
    .A2(\V2/V3/A2/A1/M4/c2 ),
    .ZN(\V2/V3/A2/c1 ));
 AND2_X1 \V2/V3/A2/A2/M1/M1/_0_  (.A1(\V2/V3/s1 [4]),
    .A2(net7),
    .ZN(\V2/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M1/M1/_1_  (.A(\V2/V3/s1 [4]),
    .B(net7),
    .Z(\V2/V3/A2/A2/M1/s1 ));
 AND2_X1 \V2/V3/A2/A2/M1/M2/_0_  (.A1(\V2/V3/A2/A2/M1/s1 ),
    .A2(\V2/V3/A2/c1 ),
    .ZN(\V2/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M1/M2/_1_  (.A(\V2/V3/A2/A2/M1/s1 ),
    .B(\V2/V3/A2/c1 ),
    .Z(\V2/V3/s2 [4]));
 OR2_X1 \V2/V3/A2/A2/M1/_0_  (.A1(\V2/V3/A2/A2/M1/c1 ),
    .A2(\V2/V3/A2/A2/M1/c2 ),
    .ZN(\V2/V3/A2/A2/c1 ));
 AND2_X1 \V2/V3/A2/A2/M2/M1/_0_  (.A1(\V2/V3/s1 [5]),
    .A2(net6),
    .ZN(\V2/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M2/M1/_1_  (.A(\V2/V3/s1 [5]),
    .B(net6),
    .Z(\V2/V3/A2/A2/M2/s1 ));
 AND2_X1 \V2/V3/A2/A2/M2/M2/_0_  (.A1(\V2/V3/A2/A2/M2/s1 ),
    .A2(\V2/V3/A2/A2/c1 ),
    .ZN(\V2/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M2/M2/_1_  (.A(\V2/V3/A2/A2/M2/s1 ),
    .B(\V2/V3/A2/A2/c1 ),
    .Z(\V2/V3/s2 [5]));
 OR2_X1 \V2/V3/A2/A2/M2/_0_  (.A1(\V2/V3/A2/A2/M2/c1 ),
    .A2(\V2/V3/A2/A2/M2/c2 ),
    .ZN(\V2/V3/A2/A2/c2 ));
 AND2_X1 \V2/V3/A2/A2/M3/M1/_0_  (.A1(\V2/V3/s1 [6]),
    .A2(net6),
    .ZN(\V2/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M3/M1/_1_  (.A(\V2/V3/s1 [6]),
    .B(net6),
    .Z(\V2/V3/A2/A2/M3/s1 ));
 AND2_X1 \V2/V3/A2/A2/M3/M2/_0_  (.A1(\V2/V3/A2/A2/M3/s1 ),
    .A2(\V2/V3/A2/A2/c2 ),
    .ZN(\V2/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M3/M2/_1_  (.A(\V2/V3/A2/A2/M3/s1 ),
    .B(\V2/V3/A2/A2/c2 ),
    .Z(\V2/V3/s2 [6]));
 OR2_X1 \V2/V3/A2/A2/M3/_0_  (.A1(\V2/V3/A2/A2/M3/c1 ),
    .A2(\V2/V3/A2/A2/M3/c2 ),
    .ZN(\V2/V3/A2/A2/c3 ));
 AND2_X1 \V2/V3/A2/A2/M4/M1/_0_  (.A1(\V2/V3/s1 [7]),
    .A2(net6),
    .ZN(\V2/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A2/A2/M4/M1/_1_  (.A(\V2/V3/s1 [7]),
    .B(net6),
    .Z(\V2/V3/A2/A2/M4/s1 ));
 AND2_X1 \V2/V3/A2/A2/M4/M2/_0_  (.A1(\V2/V3/A2/A2/M4/s1 ),
    .A2(\V2/V3/A2/A2/c3 ),
    .ZN(\V2/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A2/A2/M4/M2/_1_  (.A(\V2/V3/A2/A2/M4/s1 ),
    .B(\V2/V3/A2/A2/c3 ),
    .Z(\V2/V3/s2 [7]));
 OR2_X1 \V2/V3/A2/A2/M4/_0_  (.A1(\V2/V3/A2/A2/M4/c1 ),
    .A2(\V2/V3/A2/A2/M4/c2 ),
    .ZN(\V2/V3/c2 ));
 AND2_X1 \V2/V3/A3/A1/M1/M1/_0_  (.A1(\V2/V3/v4 [0]),
    .A2(\V2/V3/s2 [4]),
    .ZN(\V2/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M1/M1/_1_  (.A(\V2/V3/v4 [0]),
    .B(\V2/V3/s2 [4]),
    .Z(\V2/V3/A3/A1/M1/s1 ));
 AND2_X1 \V2/V3/A3/A1/M1/M2/_0_  (.A1(\V2/V3/A3/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M1/M2/_1_  (.A(\V2/V3/A3/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/v3 [8]));
 OR2_X1 \V2/V3/A3/A1/M1/_0_  (.A1(\V2/V3/A3/A1/M1/c1 ),
    .A2(\V2/V3/A3/A1/M1/c2 ),
    .ZN(\V2/V3/A3/A1/c1 ));
 AND2_X1 \V2/V3/A3/A1/M2/M1/_0_  (.A1(\V2/V3/v4 [1]),
    .A2(\V2/V3/s2 [5]),
    .ZN(\V2/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M2/M1/_1_  (.A(\V2/V3/v4 [1]),
    .B(\V2/V3/s2 [5]),
    .Z(\V2/V3/A3/A1/M2/s1 ));
 AND2_X1 \V2/V3/A3/A1/M2/M2/_0_  (.A1(\V2/V3/A3/A1/M2/s1 ),
    .A2(\V2/V3/A3/A1/c1 ),
    .ZN(\V2/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M2/M2/_1_  (.A(\V2/V3/A3/A1/M2/s1 ),
    .B(\V2/V3/A3/A1/c1 ),
    .Z(\V2/v3 [9]));
 OR2_X1 \V2/V3/A3/A1/M2/_0_  (.A1(\V2/V3/A3/A1/M2/c1 ),
    .A2(\V2/V3/A3/A1/M2/c2 ),
    .ZN(\V2/V3/A3/A1/c2 ));
 AND2_X1 \V2/V3/A3/A1/M3/M1/_0_  (.A1(\V2/V3/v4 [2]),
    .A2(\V2/V3/s2 [6]),
    .ZN(\V2/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M3/M1/_1_  (.A(\V2/V3/v4 [2]),
    .B(\V2/V3/s2 [6]),
    .Z(\V2/V3/A3/A1/M3/s1 ));
 AND2_X1 \V2/V3/A3/A1/M3/M2/_0_  (.A1(\V2/V3/A3/A1/M3/s1 ),
    .A2(\V2/V3/A3/A1/c2 ),
    .ZN(\V2/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M3/M2/_1_  (.A(\V2/V3/A3/A1/M3/s1 ),
    .B(\V2/V3/A3/A1/c2 ),
    .Z(\V2/v3 [10]));
 OR2_X1 \V2/V3/A3/A1/M3/_0_  (.A1(\V2/V3/A3/A1/M3/c1 ),
    .A2(\V2/V3/A3/A1/M3/c2 ),
    .ZN(\V2/V3/A3/A1/c3 ));
 AND2_X1 \V2/V3/A3/A1/M4/M1/_0_  (.A1(\V2/V3/v4 [3]),
    .A2(\V2/V3/s2 [7]),
    .ZN(\V2/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V3/A3/A1/M4/M1/_1_  (.A(\V2/V3/v4 [3]),
    .B(\V2/V3/s2 [7]),
    .Z(\V2/V3/A3/A1/M4/s1 ));
 AND2_X1 \V2/V3/A3/A1/M4/M2/_0_  (.A1(\V2/V3/A3/A1/M4/s1 ),
    .A2(\V2/V3/A3/A1/c3 ),
    .ZN(\V2/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V3/A3/A1/M4/M2/_1_  (.A(\V2/V3/A3/A1/M4/s1 ),
    .B(\V2/V3/A3/A1/c3 ),
    .Z(\V2/v3 [11]));
 OR2_X1 \V2/V3/A3/A1/M4/_0_  (.A1(\V2/V3/A3/A1/M4/c1 ),
    .A2(\V2/V3/A3/A1/M4/c2 ),
    .ZN(\V2/V3/A3/c1 ));
 AND2_X1 \V2/V3/A3/A2/M1/M1/_0_  (.A1(\V2/V3/v4 [4]),
    .A2(\V2/V3/c3 ),
    .ZN(\V2/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M1/M1/_1_  (.A(\V2/V3/v4 [4]),
    .B(\V2/V3/c3 ),
    .Z(\V2/V3/A3/A2/M1/s1 ));
 AND2_X1 \V2/V3/A3/A2/M1/M2/_0_  (.A1(\V2/V3/A3/A2/M1/s1 ),
    .A2(\V2/V3/A3/c1 ),
    .ZN(\V2/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M1/M2/_1_  (.A(\V2/V3/A3/A2/M1/s1 ),
    .B(\V2/V3/A3/c1 ),
    .Z(\V2/v3 [12]));
 OR2_X1 \V2/V3/A3/A2/M1/_0_  (.A1(\V2/V3/A3/A2/M1/c1 ),
    .A2(\V2/V3/A3/A2/M1/c2 ),
    .ZN(\V2/V3/A3/A2/c1 ));
 AND2_X1 \V2/V3/A3/A2/M2/M1/_0_  (.A1(\V2/V3/v4 [5]),
    .A2(net7),
    .ZN(\V2/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M2/M1/_1_  (.A(\V2/V3/v4 [5]),
    .B(net7),
    .Z(\V2/V3/A3/A2/M2/s1 ));
 AND2_X1 \V2/V3/A3/A2/M2/M2/_0_  (.A1(\V2/V3/A3/A2/M2/s1 ),
    .A2(\V2/V3/A3/A2/c1 ),
    .ZN(\V2/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M2/M2/_1_  (.A(\V2/V3/A3/A2/M2/s1 ),
    .B(\V2/V3/A3/A2/c1 ),
    .Z(\V2/v3 [13]));
 OR2_X1 \V2/V3/A3/A2/M2/_0_  (.A1(\V2/V3/A3/A2/M2/c1 ),
    .A2(\V2/V3/A3/A2/M2/c2 ),
    .ZN(\V2/V3/A3/A2/c2 ));
 AND2_X1 \V2/V3/A3/A2/M3/M1/_0_  (.A1(\V2/V3/v4 [6]),
    .A2(net7),
    .ZN(\V2/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M3/M1/_1_  (.A(\V2/V3/v4 [6]),
    .B(net7),
    .Z(\V2/V3/A3/A2/M3/s1 ));
 AND2_X1 \V2/V3/A3/A2/M3/M2/_0_  (.A1(\V2/V3/A3/A2/M3/s1 ),
    .A2(\V2/V3/A3/A2/c2 ),
    .ZN(\V2/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M3/M2/_1_  (.A(\V2/V3/A3/A2/M3/s1 ),
    .B(\V2/V3/A3/A2/c2 ),
    .Z(\V2/v3 [14]));
 OR2_X1 \V2/V3/A3/A2/M3/_0_  (.A1(\V2/V3/A3/A2/M3/c1 ),
    .A2(\V2/V3/A3/A2/M3/c2 ),
    .ZN(\V2/V3/A3/A2/c3 ));
 AND2_X1 \V2/V3/A3/A2/M4/M1/_0_  (.A1(\V2/V3/v4 [7]),
    .A2(net7),
    .ZN(\V2/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V3/A3/A2/M4/M1/_1_  (.A(\V2/V3/v4 [7]),
    .B(net7),
    .Z(\V2/V3/A3/A2/M4/s1 ));
 AND2_X1 \V2/V3/A3/A2/M4/M2/_0_  (.A1(\V2/V3/A3/A2/M4/s1 ),
    .A2(\V2/V3/A3/A2/c3 ),
    .ZN(\V2/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V3/A3/A2/M4/M2/_1_  (.A(\V2/V3/A3/A2/M4/s1 ),
    .B(\V2/V3/A3/A2/c3 ),
    .Z(\V2/v3 [15]));
 OR2_X1 \V2/V3/A3/A2/M4/_0_  (.A1(\V2/V3/A3/A2/M4/c1 ),
    .A2(\V2/V3/A3/A2/M4/c2 ),
    .ZN(\V2/V3/overflow ));
 AND2_X1 \V2/V3/V1/A1/M1/M1/_0_  (.A1(\V2/V3/V1/v2 [0]),
    .A2(\V2/V3/V1/v3 [0]),
    .ZN(\V2/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M1/M1/_1_  (.A(\V2/V3/V1/v2 [0]),
    .B(\V2/V3/V1/v3 [0]),
    .Z(\V2/V3/V1/A1/M1/s1 ));
 AND2_X1 \V2/V3/V1/A1/M1/M2/_0_  (.A1(\V2/V3/V1/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M1/M2/_1_  (.A(\V2/V3/V1/A1/M1/s1 ),
    .B(net2),
    .Z(\V2/V3/V1/s1 [0]));
 OR2_X1 \V2/V3/V1/A1/M1/_0_  (.A1(\V2/V3/V1/A1/M1/c1 ),
    .A2(\V2/V3/V1/A1/M1/c2 ),
    .ZN(\V2/V3/V1/A1/c1 ));
 AND2_X1 \V2/V3/V1/A1/M2/M1/_0_  (.A1(\V2/V3/V1/v2 [1]),
    .A2(\V2/V3/V1/v3 [1]),
    .ZN(\V2/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M2/M1/_1_  (.A(\V2/V3/V1/v2 [1]),
    .B(\V2/V3/V1/v3 [1]),
    .Z(\V2/V3/V1/A1/M2/s1 ));
 AND2_X1 \V2/V3/V1/A1/M2/M2/_0_  (.A1(\V2/V3/V1/A1/M2/s1 ),
    .A2(\V2/V3/V1/A1/c1 ),
    .ZN(\V2/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M2/M2/_1_  (.A(\V2/V3/V1/A1/M2/s1 ),
    .B(\V2/V3/V1/A1/c1 ),
    .Z(\V2/V3/V1/s1 [1]));
 OR2_X1 \V2/V3/V1/A1/M2/_0_  (.A1(\V2/V3/V1/A1/M2/c1 ),
    .A2(\V2/V3/V1/A1/M2/c2 ),
    .ZN(\V2/V3/V1/A1/c2 ));
 AND2_X1 \V2/V3/V1/A1/M3/M1/_0_  (.A1(\V2/V3/V1/v2 [2]),
    .A2(\V2/V3/V1/v3 [2]),
    .ZN(\V2/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M3/M1/_1_  (.A(\V2/V3/V1/v2 [2]),
    .B(\V2/V3/V1/v3 [2]),
    .Z(\V2/V3/V1/A1/M3/s1 ));
 AND2_X1 \V2/V3/V1/A1/M3/M2/_0_  (.A1(\V2/V3/V1/A1/M3/s1 ),
    .A2(\V2/V3/V1/A1/c2 ),
    .ZN(\V2/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M3/M2/_1_  (.A(\V2/V3/V1/A1/M3/s1 ),
    .B(\V2/V3/V1/A1/c2 ),
    .Z(\V2/V3/V1/s1 [2]));
 OR2_X1 \V2/V3/V1/A1/M3/_0_  (.A1(\V2/V3/V1/A1/M3/c1 ),
    .A2(\V2/V3/V1/A1/M3/c2 ),
    .ZN(\V2/V3/V1/A1/c3 ));
 AND2_X1 \V2/V3/V1/A1/M4/M1/_0_  (.A1(\V2/V3/V1/v2 [3]),
    .A2(\V2/V3/V1/v3 [3]),
    .ZN(\V2/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A1/M4/M1/_1_  (.A(\V2/V3/V1/v2 [3]),
    .B(\V2/V3/V1/v3 [3]),
    .Z(\V2/V3/V1/A1/M4/s1 ));
 AND2_X1 \V2/V3/V1/A1/M4/M2/_0_  (.A1(\V2/V3/V1/A1/M4/s1 ),
    .A2(\V2/V3/V1/A1/c3 ),
    .ZN(\V2/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A1/M4/M2/_1_  (.A(\V2/V3/V1/A1/M4/s1 ),
    .B(\V2/V3/V1/A1/c3 ),
    .Z(\V2/V3/V1/s1 [3]));
 OR2_X1 \V2/V3/V1/A1/M4/_0_  (.A1(\V2/V3/V1/A1/M4/c1 ),
    .A2(\V2/V3/V1/A1/M4/c2 ),
    .ZN(\V2/V3/V1/c1 ));
 AND2_X1 \V2/V3/V1/A2/M1/M1/_0_  (.A1(\V2/V3/V1/s1 [0]),
    .A2(\V2/V3/V1/v1 [2]),
    .ZN(\V2/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M1/M1/_1_  (.A(\V2/V3/V1/s1 [0]),
    .B(\V2/V3/V1/v1 [2]),
    .Z(\V2/V3/V1/A2/M1/s1 ));
 AND2_X1 \V2/V3/V1/A2/M1/M2/_0_  (.A1(\V2/V3/V1/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M1/M2/_1_  (.A(\V2/V3/V1/A2/M1/s1 ),
    .B(net2),
    .Z(\V2/v3 [2]));
 OR2_X1 \V2/V3/V1/A2/M1/_0_  (.A1(\V2/V3/V1/A2/M1/c1 ),
    .A2(\V2/V3/V1/A2/M1/c2 ),
    .ZN(\V2/V3/V1/A2/c1 ));
 AND2_X1 \V2/V3/V1/A2/M2/M1/_0_  (.A1(\V2/V3/V1/s1 [1]),
    .A2(\V2/V3/V1/v1 [3]),
    .ZN(\V2/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M2/M1/_1_  (.A(\V2/V3/V1/s1 [1]),
    .B(\V2/V3/V1/v1 [3]),
    .Z(\V2/V3/V1/A2/M2/s1 ));
 AND2_X1 \V2/V3/V1/A2/M2/M2/_0_  (.A1(\V2/V3/V1/A2/M2/s1 ),
    .A2(\V2/V3/V1/A2/c1 ),
    .ZN(\V2/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M2/M2/_1_  (.A(\V2/V3/V1/A2/M2/s1 ),
    .B(\V2/V3/V1/A2/c1 ),
    .Z(\V2/v3 [3]));
 OR2_X1 \V2/V3/V1/A2/M2/_0_  (.A1(\V2/V3/V1/A2/M2/c1 ),
    .A2(\V2/V3/V1/A2/M2/c2 ),
    .ZN(\V2/V3/V1/A2/c2 ));
 AND2_X1 \V2/V3/V1/A2/M3/M1/_0_  (.A1(\V2/V3/V1/s1 [2]),
    .A2(net2),
    .ZN(\V2/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M3/M1/_1_  (.A(\V2/V3/V1/s1 [2]),
    .B(net2),
    .Z(\V2/V3/V1/A2/M3/s1 ));
 AND2_X1 \V2/V3/V1/A2/M3/M2/_0_  (.A1(\V2/V3/V1/A2/M3/s1 ),
    .A2(\V2/V3/V1/A2/c2 ),
    .ZN(\V2/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M3/M2/_1_  (.A(\V2/V3/V1/A2/M3/s1 ),
    .B(\V2/V3/V1/A2/c2 ),
    .Z(\V2/V3/V1/s2 [2]));
 OR2_X1 \V2/V3/V1/A2/M3/_0_  (.A1(\V2/V3/V1/A2/M3/c1 ),
    .A2(\V2/V3/V1/A2/M3/c2 ),
    .ZN(\V2/V3/V1/A2/c3 ));
 AND2_X1 \V2/V3/V1/A2/M4/M1/_0_  (.A1(\V2/V3/V1/s1 [3]),
    .A2(net2),
    .ZN(\V2/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A2/M4/M1/_1_  (.A(\V2/V3/V1/s1 [3]),
    .B(net2),
    .Z(\V2/V3/V1/A2/M4/s1 ));
 AND2_X1 \V2/V3/V1/A2/M4/M2/_0_  (.A1(\V2/V3/V1/A2/M4/s1 ),
    .A2(\V2/V3/V1/A2/c3 ),
    .ZN(\V2/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A2/M4/M2/_1_  (.A(\V2/V3/V1/A2/M4/s1 ),
    .B(\V2/V3/V1/A2/c3 ),
    .Z(\V2/V3/V1/s2 [3]));
 OR2_X1 \V2/V3/V1/A2/M4/_0_  (.A1(\V2/V3/V1/A2/M4/c1 ),
    .A2(\V2/V3/V1/A2/M4/c2 ),
    .ZN(\V2/V3/V1/c2 ));
 AND2_X1 \V2/V3/V1/A3/M1/M1/_0_  (.A1(\V2/V3/V1/v4 [0]),
    .A2(\V2/V3/V1/s2 [2]),
    .ZN(\V2/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M1/M1/_1_  (.A(\V2/V3/V1/v4 [0]),
    .B(\V2/V3/V1/s2 [2]),
    .Z(\V2/V3/V1/A3/M1/s1 ));
 AND2_X1 \V2/V3/V1/A3/M1/M2/_0_  (.A1(\V2/V3/V1/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V2/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M1/M2/_1_  (.A(\V2/V3/V1/A3/M1/s1 ),
    .B(net2),
    .Z(\V2/V3/v1 [4]));
 OR2_X1 \V2/V3/V1/A3/M1/_0_  (.A1(\V2/V3/V1/A3/M1/c1 ),
    .A2(\V2/V3/V1/A3/M1/c2 ),
    .ZN(\V2/V3/V1/A3/c1 ));
 AND2_X1 \V2/V3/V1/A3/M2/M1/_0_  (.A1(\V2/V3/V1/v4 [1]),
    .A2(\V2/V3/V1/s2 [3]),
    .ZN(\V2/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M2/M1/_1_  (.A(\V2/V3/V1/v4 [1]),
    .B(\V2/V3/V1/s2 [3]),
    .Z(\V2/V3/V1/A3/M2/s1 ));
 AND2_X1 \V2/V3/V1/A3/M2/M2/_0_  (.A1(\V2/V3/V1/A3/M2/s1 ),
    .A2(\V2/V3/V1/A3/c1 ),
    .ZN(\V2/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M2/M2/_1_  (.A(\V2/V3/V1/A3/M2/s1 ),
    .B(\V2/V3/V1/A3/c1 ),
    .Z(\V2/V3/v1 [5]));
 OR2_X1 \V2/V3/V1/A3/M2/_0_  (.A1(\V2/V3/V1/A3/M2/c1 ),
    .A2(\V2/V3/V1/A3/M2/c2 ),
    .ZN(\V2/V3/V1/A3/c2 ));
 AND2_X1 \V2/V3/V1/A3/M3/M1/_0_  (.A1(\V2/V3/V1/v4 [2]),
    .A2(\V2/V3/V1/c3 ),
    .ZN(\V2/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M3/M1/_1_  (.A(\V2/V3/V1/v4 [2]),
    .B(\V2/V3/V1/c3 ),
    .Z(\V2/V3/V1/A3/M3/s1 ));
 AND2_X1 \V2/V3/V1/A3/M3/M2/_0_  (.A1(\V2/V3/V1/A3/M3/s1 ),
    .A2(\V2/V3/V1/A3/c2 ),
    .ZN(\V2/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M3/M2/_1_  (.A(\V2/V3/V1/A3/M3/s1 ),
    .B(\V2/V3/V1/A3/c2 ),
    .Z(\V2/V3/v1 [6]));
 OR2_X1 \V2/V3/V1/A3/M3/_0_  (.A1(\V2/V3/V1/A3/M3/c1 ),
    .A2(\V2/V3/V1/A3/M3/c2 ),
    .ZN(\V2/V3/V1/A3/c3 ));
 AND2_X1 \V2/V3/V1/A3/M4/M1/_0_  (.A1(\V2/V3/V1/v4 [3]),
    .A2(net7),
    .ZN(\V2/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V1/A3/M4/M1/_1_  (.A(\V2/V3/V1/v4 [3]),
    .B(net7),
    .Z(\V2/V3/V1/A3/M4/s1 ));
 AND2_X1 \V2/V3/V1/A3/M4/M2/_0_  (.A1(\V2/V3/V1/A3/M4/s1 ),
    .A2(\V2/V3/V1/A3/c3 ),
    .ZN(\V2/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V1/A3/M4/M2/_1_  (.A(\V2/V3/V1/A3/M4/s1 ),
    .B(\V2/V3/V1/A3/c3 ),
    .Z(\V2/V3/v1 [7]));
 OR2_X1 \V2/V3/V1/A3/M4/_0_  (.A1(\V2/V3/V1/A3/M4/c1 ),
    .A2(\V2/V3/V1/A3/M4/c2 ),
    .ZN(\V2/V3/V1/overflow ));
 AND2_X1 \V2/V3/V1/V1/HA1/_0_  (.A1(\V2/V3/V1/V1/w2 ),
    .A2(\V2/V3/V1/V1/w1 ),
    .ZN(\V2/V3/V1/V1/w4 ));
 XOR2_X2 \V2/V3/V1/V1/HA1/_1_  (.A(\V2/V3/V1/V1/w2 ),
    .B(\V2/V3/V1/V1/w1 ),
    .Z(\V2/v3 [1]));
 AND2_X1 \V2/V3/V1/V1/HA2/_0_  (.A1(\V2/V3/V1/V1/w4 ),
    .A2(\V2/V3/V1/V1/w3 ),
    .ZN(\V2/V3/V1/v1 [3]));
 XOR2_X2 \V2/V3/V1/V1/HA2/_1_  (.A(\V2/V3/V1/V1/w4 ),
    .B(\V2/V3/V1/V1/w3 ),
    .Z(\V2/V3/V1/v1 [2]));
 AND2_X1 \V2/V3/V1/V1/_0_  (.A1(net41),
    .A2(net12),
    .ZN(\V2/v3 [0]));
 AND2_X1 \V2/V3/V1/V1/_1_  (.A1(net41),
    .A2(net11),
    .ZN(\V2/V3/V1/V1/w1 ));
 AND2_X1 \V2/V3/V1/V1/_2_  (.A1(net12),
    .A2(net40),
    .ZN(\V2/V3/V1/V1/w2 ));
 AND2_X1 \V2/V3/V1/V1/_3_  (.A1(net11),
    .A2(net40),
    .ZN(\V2/V3/V1/V1/w3 ));
 AND2_X1 \V2/V3/V1/V2/HA1/_0_  (.A1(\V2/V3/V1/V2/w2 ),
    .A2(\V2/V3/V1/V2/w1 ),
    .ZN(\V2/V3/V1/V2/w4 ));
 XOR2_X2 \V2/V3/V1/V2/HA1/_1_  (.A(\V2/V3/V1/V2/w2 ),
    .B(\V2/V3/V1/V2/w1 ),
    .Z(\V2/V3/V1/v2 [1]));
 AND2_X1 \V2/V3/V1/V2/HA2/_0_  (.A1(\V2/V3/V1/V2/w4 ),
    .A2(\V2/V3/V1/V2/w3 ),
    .ZN(\V2/V3/V1/v2 [3]));
 XOR2_X2 \V2/V3/V1/V2/HA2/_1_  (.A(\V2/V3/V1/V2/w4 ),
    .B(\V2/V3/V1/V2/w3 ),
    .Z(\V2/V3/V1/v2 [2]));
 AND2_X1 \V2/V3/V1/V2/_0_  (.A1(net39),
    .A2(net12),
    .ZN(\V2/V3/V1/v2 [0]));
 AND2_X1 \V2/V3/V1/V2/_1_  (.A1(net39),
    .A2(net11),
    .ZN(\V2/V3/V1/V2/w1 ));
 AND2_X1 \V2/V3/V1/V2/_2_  (.A1(net12),
    .A2(net38),
    .ZN(\V2/V3/V1/V2/w2 ));
 AND2_X1 \V2/V3/V1/V2/_3_  (.A1(net11),
    .A2(net38),
    .ZN(\V2/V3/V1/V2/w3 ));
 AND2_X1 \V2/V3/V1/V3/HA1/_0_  (.A1(\V2/V3/V1/V3/w2 ),
    .A2(\V2/V3/V1/V3/w1 ),
    .ZN(\V2/V3/V1/V3/w4 ));
 XOR2_X2 \V2/V3/V1/V3/HA1/_1_  (.A(\V2/V3/V1/V3/w2 ),
    .B(\V2/V3/V1/V3/w1 ),
    .Z(\V2/V3/V1/v3 [1]));
 AND2_X1 \V2/V3/V1/V3/HA2/_0_  (.A1(\V2/V3/V1/V3/w4 ),
    .A2(\V2/V3/V1/V3/w3 ),
    .ZN(\V2/V3/V1/v3 [3]));
 XOR2_X2 \V2/V3/V1/V3/HA2/_1_  (.A(\V2/V3/V1/V3/w4 ),
    .B(\V2/V3/V1/V3/w3 ),
    .Z(\V2/V3/V1/v3 [2]));
 AND2_X1 \V2/V3/V1/V3/_0_  (.A1(net41),
    .A2(B[10]),
    .ZN(\V2/V3/V1/v3 [0]));
 AND2_X1 \V2/V3/V1/V3/_1_  (.A1(net41),
    .A2(B[11]),
    .ZN(\V2/V3/V1/V3/w1 ));
 AND2_X1 \V2/V3/V1/V3/_2_  (.A1(B[10]),
    .A2(net40),
    .ZN(\V2/V3/V1/V3/w2 ));
 AND2_X1 \V2/V3/V1/V3/_3_  (.A1(B[11]),
    .A2(net40),
    .ZN(\V2/V3/V1/V3/w3 ));
 AND2_X1 \V2/V3/V1/V4/HA1/_0_  (.A1(\V2/V3/V1/V4/w2 ),
    .A2(\V2/V3/V1/V4/w1 ),
    .ZN(\V2/V3/V1/V4/w4 ));
 XOR2_X2 \V2/V3/V1/V4/HA1/_1_  (.A(\V2/V3/V1/V4/w2 ),
    .B(\V2/V3/V1/V4/w1 ),
    .Z(\V2/V3/V1/v4 [1]));
 AND2_X1 \V2/V3/V1/V4/HA2/_0_  (.A1(\V2/V3/V1/V4/w4 ),
    .A2(\V2/V3/V1/V4/w3 ),
    .ZN(\V2/V3/V1/v4 [3]));
 XOR2_X2 \V2/V3/V1/V4/HA2/_1_  (.A(\V2/V3/V1/V4/w4 ),
    .B(\V2/V3/V1/V4/w3 ),
    .Z(\V2/V3/V1/v4 [2]));
 AND2_X1 \V2/V3/V1/V4/_0_  (.A1(net39),
    .A2(B[10]),
    .ZN(\V2/V3/V1/v4 [0]));
 AND2_X1 \V2/V3/V1/V4/_1_  (.A1(net39),
    .A2(B[11]),
    .ZN(\V2/V3/V1/V4/w1 ));
 AND2_X1 \V2/V3/V1/V4/_2_  (.A1(B[10]),
    .A2(net38),
    .ZN(\V2/V3/V1/V4/w2 ));
 AND2_X1 \V2/V3/V1/V4/_3_  (.A1(B[11]),
    .A2(net38),
    .ZN(\V2/V3/V1/V4/w3 ));
 OR2_X1 \V2/V3/V1/_0_  (.A1(\V2/V3/V1/c1 ),
    .A2(\V2/V3/V1/c2 ),
    .ZN(\V2/V3/V1/c3 ));
 AND2_X1 \V2/V3/V2/A1/M1/M1/_0_  (.A1(\V2/V3/V2/v2 [0]),
    .A2(\V2/V3/V2/v3 [0]),
    .ZN(\V2/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M1/M1/_1_  (.A(\V2/V3/V2/v2 [0]),
    .B(\V2/V3/V2/v3 [0]),
    .Z(\V2/V3/V2/A1/M1/s1 ));
 AND2_X1 \V2/V3/V2/A1/M1/M2/_0_  (.A1(\V2/V3/V2/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M1/M2/_1_  (.A(\V2/V3/V2/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/V2/s1 [0]));
 OR2_X1 \V2/V3/V2/A1/M1/_0_  (.A1(\V2/V3/V2/A1/M1/c1 ),
    .A2(\V2/V3/V2/A1/M1/c2 ),
    .ZN(\V2/V3/V2/A1/c1 ));
 AND2_X1 \V2/V3/V2/A1/M2/M1/_0_  (.A1(\V2/V3/V2/v2 [1]),
    .A2(\V2/V3/V2/v3 [1]),
    .ZN(\V2/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M2/M1/_1_  (.A(\V2/V3/V2/v2 [1]),
    .B(\V2/V3/V2/v3 [1]),
    .Z(\V2/V3/V2/A1/M2/s1 ));
 AND2_X1 \V2/V3/V2/A1/M2/M2/_0_  (.A1(\V2/V3/V2/A1/M2/s1 ),
    .A2(\V2/V3/V2/A1/c1 ),
    .ZN(\V2/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M2/M2/_1_  (.A(\V2/V3/V2/A1/M2/s1 ),
    .B(\V2/V3/V2/A1/c1 ),
    .Z(\V2/V3/V2/s1 [1]));
 OR2_X1 \V2/V3/V2/A1/M2/_0_  (.A1(\V2/V3/V2/A1/M2/c1 ),
    .A2(\V2/V3/V2/A1/M2/c2 ),
    .ZN(\V2/V3/V2/A1/c2 ));
 AND2_X1 \V2/V3/V2/A1/M3/M1/_0_  (.A1(\V2/V3/V2/v2 [2]),
    .A2(\V2/V3/V2/v3 [2]),
    .ZN(\V2/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M3/M1/_1_  (.A(\V2/V3/V2/v2 [2]),
    .B(\V2/V3/V2/v3 [2]),
    .Z(\V2/V3/V2/A1/M3/s1 ));
 AND2_X1 \V2/V3/V2/A1/M3/M2/_0_  (.A1(\V2/V3/V2/A1/M3/s1 ),
    .A2(\V2/V3/V2/A1/c2 ),
    .ZN(\V2/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M3/M2/_1_  (.A(\V2/V3/V2/A1/M3/s1 ),
    .B(\V2/V3/V2/A1/c2 ),
    .Z(\V2/V3/V2/s1 [2]));
 OR2_X1 \V2/V3/V2/A1/M3/_0_  (.A1(\V2/V3/V2/A1/M3/c1 ),
    .A2(\V2/V3/V2/A1/M3/c2 ),
    .ZN(\V2/V3/V2/A1/c3 ));
 AND2_X1 \V2/V3/V2/A1/M4/M1/_0_  (.A1(\V2/V3/V2/v2 [3]),
    .A2(\V2/V3/V2/v3 [3]),
    .ZN(\V2/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A1/M4/M1/_1_  (.A(\V2/V3/V2/v2 [3]),
    .B(\V2/V3/V2/v3 [3]),
    .Z(\V2/V3/V2/A1/M4/s1 ));
 AND2_X1 \V2/V3/V2/A1/M4/M2/_0_  (.A1(\V2/V3/V2/A1/M4/s1 ),
    .A2(\V2/V3/V2/A1/c3 ),
    .ZN(\V2/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A1/M4/M2/_1_  (.A(\V2/V3/V2/A1/M4/s1 ),
    .B(\V2/V3/V2/A1/c3 ),
    .Z(\V2/V3/V2/s1 [3]));
 OR2_X1 \V2/V3/V2/A1/M4/_0_  (.A1(\V2/V3/V2/A1/M4/c1 ),
    .A2(\V2/V3/V2/A1/M4/c2 ),
    .ZN(\V2/V3/V2/c1 ));
 AND2_X1 \V2/V3/V2/A2/M1/M1/_0_  (.A1(\V2/V3/V2/s1 [0]),
    .A2(\V2/V3/V2/v1 [2]),
    .ZN(\V2/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M1/M1/_1_  (.A(\V2/V3/V2/s1 [0]),
    .B(\V2/V3/V2/v1 [2]),
    .Z(\V2/V3/V2/A2/M1/s1 ));
 AND2_X1 \V2/V3/V2/A2/M1/M2/_0_  (.A1(\V2/V3/V2/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M1/M2/_1_  (.A(\V2/V3/V2/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/v2 [2]));
 OR2_X1 \V2/V3/V2/A2/M1/_0_  (.A1(\V2/V3/V2/A2/M1/c1 ),
    .A2(\V2/V3/V2/A2/M1/c2 ),
    .ZN(\V2/V3/V2/A2/c1 ));
 AND2_X1 \V2/V3/V2/A2/M2/M1/_0_  (.A1(\V2/V3/V2/s1 [1]),
    .A2(\V2/V3/V2/v1 [3]),
    .ZN(\V2/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M2/M1/_1_  (.A(\V2/V3/V2/s1 [1]),
    .B(\V2/V3/V2/v1 [3]),
    .Z(\V2/V3/V2/A2/M2/s1 ));
 AND2_X1 \V2/V3/V2/A2/M2/M2/_0_  (.A1(\V2/V3/V2/A2/M2/s1 ),
    .A2(\V2/V3/V2/A2/c1 ),
    .ZN(\V2/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M2/M2/_1_  (.A(\V2/V3/V2/A2/M2/s1 ),
    .B(\V2/V3/V2/A2/c1 ),
    .Z(\V2/V3/v2 [3]));
 OR2_X1 \V2/V3/V2/A2/M2/_0_  (.A1(\V2/V3/V2/A2/M2/c1 ),
    .A2(\V2/V3/V2/A2/M2/c2 ),
    .ZN(\V2/V3/V2/A2/c2 ));
 AND2_X1 \V2/V3/V2/A2/M3/M1/_0_  (.A1(\V2/V3/V2/s1 [2]),
    .A2(net6),
    .ZN(\V2/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M3/M1/_1_  (.A(\V2/V3/V2/s1 [2]),
    .B(net6),
    .Z(\V2/V3/V2/A2/M3/s1 ));
 AND2_X1 \V2/V3/V2/A2/M3/M2/_0_  (.A1(\V2/V3/V2/A2/M3/s1 ),
    .A2(\V2/V3/V2/A2/c2 ),
    .ZN(\V2/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M3/M2/_1_  (.A(\V2/V3/V2/A2/M3/s1 ),
    .B(\V2/V3/V2/A2/c2 ),
    .Z(\V2/V3/V2/s2 [2]));
 OR2_X1 \V2/V3/V2/A2/M3/_0_  (.A1(\V2/V3/V2/A2/M3/c1 ),
    .A2(\V2/V3/V2/A2/M3/c2 ),
    .ZN(\V2/V3/V2/A2/c3 ));
 AND2_X1 \V2/V3/V2/A2/M4/M1/_0_  (.A1(\V2/V3/V2/s1 [3]),
    .A2(net6),
    .ZN(\V2/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A2/M4/M1/_1_  (.A(\V2/V3/V2/s1 [3]),
    .B(net6),
    .Z(\V2/V3/V2/A2/M4/s1 ));
 AND2_X1 \V2/V3/V2/A2/M4/M2/_0_  (.A1(\V2/V3/V2/A2/M4/s1 ),
    .A2(\V2/V3/V2/A2/c3 ),
    .ZN(\V2/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A2/M4/M2/_1_  (.A(\V2/V3/V2/A2/M4/s1 ),
    .B(\V2/V3/V2/A2/c3 ),
    .Z(\V2/V3/V2/s2 [3]));
 OR2_X1 \V2/V3/V2/A2/M4/_0_  (.A1(\V2/V3/V2/A2/M4/c1 ),
    .A2(\V2/V3/V2/A2/M4/c2 ),
    .ZN(\V2/V3/V2/c2 ));
 AND2_X1 \V2/V3/V2/A3/M1/M1/_0_  (.A1(\V2/V3/V2/v4 [0]),
    .A2(\V2/V3/V2/s2 [2]),
    .ZN(\V2/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M1/M1/_1_  (.A(\V2/V3/V2/v4 [0]),
    .B(\V2/V3/V2/s2 [2]),
    .Z(\V2/V3/V2/A3/M1/s1 ));
 AND2_X1 \V2/V3/V2/A3/M1/M2/_0_  (.A1(\V2/V3/V2/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V2/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M1/M2/_1_  (.A(\V2/V3/V2/A3/M1/s1 ),
    .B(net6),
    .Z(\V2/V3/v2 [4]));
 OR2_X1 \V2/V3/V2/A3/M1/_0_  (.A1(\V2/V3/V2/A3/M1/c1 ),
    .A2(\V2/V3/V2/A3/M1/c2 ),
    .ZN(\V2/V3/V2/A3/c1 ));
 AND2_X1 \V2/V3/V2/A3/M2/M1/_0_  (.A1(\V2/V3/V2/v4 [1]),
    .A2(\V2/V3/V2/s2 [3]),
    .ZN(\V2/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M2/M1/_1_  (.A(\V2/V3/V2/v4 [1]),
    .B(\V2/V3/V2/s2 [3]),
    .Z(\V2/V3/V2/A3/M2/s1 ));
 AND2_X1 \V2/V3/V2/A3/M2/M2/_0_  (.A1(\V2/V3/V2/A3/M2/s1 ),
    .A2(\V2/V3/V2/A3/c1 ),
    .ZN(\V2/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M2/M2/_1_  (.A(\V2/V3/V2/A3/M2/s1 ),
    .B(\V2/V3/V2/A3/c1 ),
    .Z(\V2/V3/v2 [5]));
 OR2_X1 \V2/V3/V2/A3/M2/_0_  (.A1(\V2/V3/V2/A3/M2/c1 ),
    .A2(\V2/V3/V2/A3/M2/c2 ),
    .ZN(\V2/V3/V2/A3/c2 ));
 AND2_X1 \V2/V3/V2/A3/M3/M1/_0_  (.A1(\V2/V3/V2/v4 [2]),
    .A2(\V2/V3/V2/c3 ),
    .ZN(\V2/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M3/M1/_1_  (.A(\V2/V3/V2/v4 [2]),
    .B(\V2/V3/V2/c3 ),
    .Z(\V2/V3/V2/A3/M3/s1 ));
 AND2_X1 \V2/V3/V2/A3/M3/M2/_0_  (.A1(\V2/V3/V2/A3/M3/s1 ),
    .A2(\V2/V3/V2/A3/c2 ),
    .ZN(\V2/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M3/M2/_1_  (.A(\V2/V3/V2/A3/M3/s1 ),
    .B(\V2/V3/V2/A3/c2 ),
    .Z(\V2/V3/v2 [6]));
 OR2_X1 \V2/V3/V2/A3/M3/_0_  (.A1(\V2/V3/V2/A3/M3/c1 ),
    .A2(\V2/V3/V2/A3/M3/c2 ),
    .ZN(\V2/V3/V2/A3/c3 ));
 AND2_X1 \V2/V3/V2/A3/M4/M1/_0_  (.A1(\V2/V3/V2/v4 [3]),
    .A2(net6),
    .ZN(\V2/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V2/A3/M4/M1/_1_  (.A(\V2/V3/V2/v4 [3]),
    .B(net6),
    .Z(\V2/V3/V2/A3/M4/s1 ));
 AND2_X1 \V2/V3/V2/A3/M4/M2/_0_  (.A1(\V2/V3/V2/A3/M4/s1 ),
    .A2(\V2/V3/V2/A3/c3 ),
    .ZN(\V2/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V2/A3/M4/M2/_1_  (.A(\V2/V3/V2/A3/M4/s1 ),
    .B(\V2/V3/V2/A3/c3 ),
    .Z(\V2/V3/v2 [7]));
 OR2_X1 \V2/V3/V2/A3/M4/_0_  (.A1(\V2/V3/V2/A3/M4/c1 ),
    .A2(\V2/V3/V2/A3/M4/c2 ),
    .ZN(\V2/V3/V2/overflow ));
 AND2_X1 \V2/V3/V2/V1/HA1/_0_  (.A1(\V2/V3/V2/V1/w2 ),
    .A2(\V2/V3/V2/V1/w1 ),
    .ZN(\V2/V3/V2/V1/w4 ));
 XOR2_X2 \V2/V3/V2/V1/HA1/_1_  (.A(\V2/V3/V2/V1/w2 ),
    .B(\V2/V3/V2/V1/w1 ),
    .Z(\V2/V3/v2 [1]));
 AND2_X1 \V2/V3/V2/V1/HA2/_0_  (.A1(\V2/V3/V2/V1/w4 ),
    .A2(\V2/V3/V2/V1/w3 ),
    .ZN(\V2/V3/V2/v1 [3]));
 XOR2_X2 \V2/V3/V2/V1/HA2/_1_  (.A(\V2/V3/V2/V1/w4 ),
    .B(\V2/V3/V2/V1/w3 ),
    .Z(\V2/V3/V2/v1 [2]));
 AND2_X1 \V2/V3/V2/V1/_0_  (.A1(net37),
    .A2(net12),
    .ZN(\V2/V3/v2 [0]));
 AND2_X1 \V2/V3/V2/V1/_1_  (.A1(net37),
    .A2(net11),
    .ZN(\V2/V3/V2/V1/w1 ));
 AND2_X1 \V2/V3/V2/V1/_2_  (.A1(net12),
    .A2(net36),
    .ZN(\V2/V3/V2/V1/w2 ));
 AND2_X1 \V2/V3/V2/V1/_3_  (.A1(net11),
    .A2(net36),
    .ZN(\V2/V3/V2/V1/w3 ));
 AND2_X1 \V2/V3/V2/V2/HA1/_0_  (.A1(\V2/V3/V2/V2/w2 ),
    .A2(\V2/V3/V2/V2/w1 ),
    .ZN(\V2/V3/V2/V2/w4 ));
 XOR2_X2 \V2/V3/V2/V2/HA1/_1_  (.A(\V2/V3/V2/V2/w2 ),
    .B(\V2/V3/V2/V2/w1 ),
    .Z(\V2/V3/V2/v2 [1]));
 AND2_X1 \V2/V3/V2/V2/HA2/_0_  (.A1(\V2/V3/V2/V2/w4 ),
    .A2(\V2/V3/V2/V2/w3 ),
    .ZN(\V2/V3/V2/v2 [3]));
 XOR2_X2 \V2/V3/V2/V2/HA2/_1_  (.A(\V2/V3/V2/V2/w4 ),
    .B(\V2/V3/V2/V2/w3 ),
    .Z(\V2/V3/V2/v2 [2]));
 AND2_X1 \V2/V3/V2/V2/_0_  (.A1(net35),
    .A2(net12),
    .ZN(\V2/V3/V2/v2 [0]));
 AND2_X1 \V2/V3/V2/V2/_1_  (.A1(net35),
    .A2(net11),
    .ZN(\V2/V3/V2/V2/w1 ));
 AND2_X1 \V2/V3/V2/V2/_2_  (.A1(net12),
    .A2(net34),
    .ZN(\V2/V3/V2/V2/w2 ));
 AND2_X1 \V2/V3/V2/V2/_3_  (.A1(net11),
    .A2(net34),
    .ZN(\V2/V3/V2/V2/w3 ));
 AND2_X1 \V2/V3/V2/V3/HA1/_0_  (.A1(\V2/V3/V2/V3/w2 ),
    .A2(\V2/V3/V2/V3/w1 ),
    .ZN(\V2/V3/V2/V3/w4 ));
 XOR2_X2 \V2/V3/V2/V3/HA1/_1_  (.A(\V2/V3/V2/V3/w2 ),
    .B(\V2/V3/V2/V3/w1 ),
    .Z(\V2/V3/V2/v3 [1]));
 AND2_X1 \V2/V3/V2/V3/HA2/_0_  (.A1(\V2/V3/V2/V3/w4 ),
    .A2(\V2/V3/V2/V3/w3 ),
    .ZN(\V2/V3/V2/v3 [3]));
 XOR2_X2 \V2/V3/V2/V3/HA2/_1_  (.A(\V2/V3/V2/V3/w4 ),
    .B(\V2/V3/V2/V3/w3 ),
    .Z(\V2/V3/V2/v3 [2]));
 AND2_X1 \V2/V3/V2/V3/_0_  (.A1(net37),
    .A2(B[10]),
    .ZN(\V2/V3/V2/v3 [0]));
 AND2_X1 \V2/V3/V2/V3/_1_  (.A1(net37),
    .A2(B[11]),
    .ZN(\V2/V3/V2/V3/w1 ));
 AND2_X1 \V2/V3/V2/V3/_2_  (.A1(B[10]),
    .A2(net36),
    .ZN(\V2/V3/V2/V3/w2 ));
 AND2_X1 \V2/V3/V2/V3/_3_  (.A1(B[11]),
    .A2(net36),
    .ZN(\V2/V3/V2/V3/w3 ));
 AND2_X1 \V2/V3/V2/V4/HA1/_0_  (.A1(\V2/V3/V2/V4/w2 ),
    .A2(\V2/V3/V2/V4/w1 ),
    .ZN(\V2/V3/V2/V4/w4 ));
 XOR2_X2 \V2/V3/V2/V4/HA1/_1_  (.A(\V2/V3/V2/V4/w2 ),
    .B(\V2/V3/V2/V4/w1 ),
    .Z(\V2/V3/V2/v4 [1]));
 AND2_X1 \V2/V3/V2/V4/HA2/_0_  (.A1(\V2/V3/V2/V4/w4 ),
    .A2(\V2/V3/V2/V4/w3 ),
    .ZN(\V2/V3/V2/v4 [3]));
 XOR2_X2 \V2/V3/V2/V4/HA2/_1_  (.A(\V2/V3/V2/V4/w4 ),
    .B(\V2/V3/V2/V4/w3 ),
    .Z(\V2/V3/V2/v4 [2]));
 AND2_X1 \V2/V3/V2/V4/_0_  (.A1(net35),
    .A2(B[10]),
    .ZN(\V2/V3/V2/v4 [0]));
 AND2_X1 \V2/V3/V2/V4/_1_  (.A1(net35),
    .A2(B[11]),
    .ZN(\V2/V3/V2/V4/w1 ));
 AND2_X1 \V2/V3/V2/V4/_2_  (.A1(B[10]),
    .A2(net34),
    .ZN(\V2/V3/V2/V4/w2 ));
 AND2_X1 \V2/V3/V2/V4/_3_  (.A1(B[11]),
    .A2(net34),
    .ZN(\V2/V3/V2/V4/w3 ));
 OR2_X1 \V2/V3/V2/_0_  (.A1(\V2/V3/V2/c1 ),
    .A2(\V2/V3/V2/c2 ),
    .ZN(\V2/V3/V2/c3 ));
 AND2_X1 \V2/V3/V3/A1/M1/M1/_0_  (.A1(\V2/V3/V3/v2 [0]),
    .A2(\V2/V3/V3/v3 [0]),
    .ZN(\V2/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M1/M1/_1_  (.A(\V2/V3/V3/v2 [0]),
    .B(\V2/V3/V3/v3 [0]),
    .Z(\V2/V3/V3/A1/M1/s1 ));
 AND2_X1 \V2/V3/V3/A1/M1/M2/_0_  (.A1(\V2/V3/V3/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M1/M2/_1_  (.A(\V2/V3/V3/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/V3/s1 [0]));
 OR2_X1 \V2/V3/V3/A1/M1/_0_  (.A1(\V2/V3/V3/A1/M1/c1 ),
    .A2(\V2/V3/V3/A1/M1/c2 ),
    .ZN(\V2/V3/V3/A1/c1 ));
 AND2_X1 \V2/V3/V3/A1/M2/M1/_0_  (.A1(\V2/V3/V3/v2 [1]),
    .A2(\V2/V3/V3/v3 [1]),
    .ZN(\V2/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M2/M1/_1_  (.A(\V2/V3/V3/v2 [1]),
    .B(\V2/V3/V3/v3 [1]),
    .Z(\V2/V3/V3/A1/M2/s1 ));
 AND2_X1 \V2/V3/V3/A1/M2/M2/_0_  (.A1(\V2/V3/V3/A1/M2/s1 ),
    .A2(\V2/V3/V3/A1/c1 ),
    .ZN(\V2/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M2/M2/_1_  (.A(\V2/V3/V3/A1/M2/s1 ),
    .B(\V2/V3/V3/A1/c1 ),
    .Z(\V2/V3/V3/s1 [1]));
 OR2_X1 \V2/V3/V3/A1/M2/_0_  (.A1(\V2/V3/V3/A1/M2/c1 ),
    .A2(\V2/V3/V3/A1/M2/c2 ),
    .ZN(\V2/V3/V3/A1/c2 ));
 AND2_X1 \V2/V3/V3/A1/M3/M1/_0_  (.A1(\V2/V3/V3/v2 [2]),
    .A2(\V2/V3/V3/v3 [2]),
    .ZN(\V2/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M3/M1/_1_  (.A(\V2/V3/V3/v2 [2]),
    .B(\V2/V3/V3/v3 [2]),
    .Z(\V2/V3/V3/A1/M3/s1 ));
 AND2_X1 \V2/V3/V3/A1/M3/M2/_0_  (.A1(\V2/V3/V3/A1/M3/s1 ),
    .A2(\V2/V3/V3/A1/c2 ),
    .ZN(\V2/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M3/M2/_1_  (.A(\V2/V3/V3/A1/M3/s1 ),
    .B(\V2/V3/V3/A1/c2 ),
    .Z(\V2/V3/V3/s1 [2]));
 OR2_X1 \V2/V3/V3/A1/M3/_0_  (.A1(\V2/V3/V3/A1/M3/c1 ),
    .A2(\V2/V3/V3/A1/M3/c2 ),
    .ZN(\V2/V3/V3/A1/c3 ));
 AND2_X1 \V2/V3/V3/A1/M4/M1/_0_  (.A1(\V2/V3/V3/v2 [3]),
    .A2(\V2/V3/V3/v3 [3]),
    .ZN(\V2/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A1/M4/M1/_1_  (.A(\V2/V3/V3/v2 [3]),
    .B(\V2/V3/V3/v3 [3]),
    .Z(\V2/V3/V3/A1/M4/s1 ));
 AND2_X1 \V2/V3/V3/A1/M4/M2/_0_  (.A1(\V2/V3/V3/A1/M4/s1 ),
    .A2(\V2/V3/V3/A1/c3 ),
    .ZN(\V2/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A1/M4/M2/_1_  (.A(\V2/V3/V3/A1/M4/s1 ),
    .B(\V2/V3/V3/A1/c3 ),
    .Z(\V2/V3/V3/s1 [3]));
 OR2_X1 \V2/V3/V3/A1/M4/_0_  (.A1(\V2/V3/V3/A1/M4/c1 ),
    .A2(\V2/V3/V3/A1/M4/c2 ),
    .ZN(\V2/V3/V3/c1 ));
 AND2_X1 \V2/V3/V3/A2/M1/M1/_0_  (.A1(\V2/V3/V3/s1 [0]),
    .A2(\V2/V3/V3/v1 [2]),
    .ZN(\V2/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M1/M1/_1_  (.A(\V2/V3/V3/s1 [0]),
    .B(\V2/V3/V3/v1 [2]),
    .Z(\V2/V3/V3/A2/M1/s1 ));
 AND2_X1 \V2/V3/V3/A2/M1/M2/_0_  (.A1(\V2/V3/V3/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M1/M2/_1_  (.A(\V2/V3/V3/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/v3 [2]));
 OR2_X1 \V2/V3/V3/A2/M1/_0_  (.A1(\V2/V3/V3/A2/M1/c1 ),
    .A2(\V2/V3/V3/A2/M1/c2 ),
    .ZN(\V2/V3/V3/A2/c1 ));
 AND2_X1 \V2/V3/V3/A2/M2/M1/_0_  (.A1(\V2/V3/V3/s1 [1]),
    .A2(\V2/V3/V3/v1 [3]),
    .ZN(\V2/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M2/M1/_1_  (.A(\V2/V3/V3/s1 [1]),
    .B(\V2/V3/V3/v1 [3]),
    .Z(\V2/V3/V3/A2/M2/s1 ));
 AND2_X1 \V2/V3/V3/A2/M2/M2/_0_  (.A1(\V2/V3/V3/A2/M2/s1 ),
    .A2(\V2/V3/V3/A2/c1 ),
    .ZN(\V2/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M2/M2/_1_  (.A(\V2/V3/V3/A2/M2/s1 ),
    .B(\V2/V3/V3/A2/c1 ),
    .Z(\V2/V3/v3 [3]));
 OR2_X1 \V2/V3/V3/A2/M2/_0_  (.A1(\V2/V3/V3/A2/M2/c1 ),
    .A2(\V2/V3/V3/A2/M2/c2 ),
    .ZN(\V2/V3/V3/A2/c2 ));
 AND2_X1 \V2/V3/V3/A2/M3/M1/_0_  (.A1(\V2/V3/V3/s1 [2]),
    .A2(net6),
    .ZN(\V2/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M3/M1/_1_  (.A(\V2/V3/V3/s1 [2]),
    .B(net6),
    .Z(\V2/V3/V3/A2/M3/s1 ));
 AND2_X1 \V2/V3/V3/A2/M3/M2/_0_  (.A1(\V2/V3/V3/A2/M3/s1 ),
    .A2(\V2/V3/V3/A2/c2 ),
    .ZN(\V2/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M3/M2/_1_  (.A(\V2/V3/V3/A2/M3/s1 ),
    .B(\V2/V3/V3/A2/c2 ),
    .Z(\V2/V3/V3/s2 [2]));
 OR2_X1 \V2/V3/V3/A2/M3/_0_  (.A1(\V2/V3/V3/A2/M3/c1 ),
    .A2(\V2/V3/V3/A2/M3/c2 ),
    .ZN(\V2/V3/V3/A2/c3 ));
 AND2_X1 \V2/V3/V3/A2/M4/M1/_0_  (.A1(\V2/V3/V3/s1 [3]),
    .A2(net6),
    .ZN(\V2/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A2/M4/M1/_1_  (.A(\V2/V3/V3/s1 [3]),
    .B(net6),
    .Z(\V2/V3/V3/A2/M4/s1 ));
 AND2_X1 \V2/V3/V3/A2/M4/M2/_0_  (.A1(\V2/V3/V3/A2/M4/s1 ),
    .A2(\V2/V3/V3/A2/c3 ),
    .ZN(\V2/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A2/M4/M2/_1_  (.A(\V2/V3/V3/A2/M4/s1 ),
    .B(\V2/V3/V3/A2/c3 ),
    .Z(\V2/V3/V3/s2 [3]));
 OR2_X1 \V2/V3/V3/A2/M4/_0_  (.A1(\V2/V3/V3/A2/M4/c1 ),
    .A2(\V2/V3/V3/A2/M4/c2 ),
    .ZN(\V2/V3/V3/c2 ));
 AND2_X1 \V2/V3/V3/A3/M1/M1/_0_  (.A1(\V2/V3/V3/v4 [0]),
    .A2(\V2/V3/V3/s2 [2]),
    .ZN(\V2/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M1/M1/_1_  (.A(\V2/V3/V3/v4 [0]),
    .B(\V2/V3/V3/s2 [2]),
    .Z(\V2/V3/V3/A3/M1/s1 ));
 AND2_X1 \V2/V3/V3/A3/M1/M2/_0_  (.A1(\V2/V3/V3/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V2/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M1/M2/_1_  (.A(\V2/V3/V3/A3/M1/s1 ),
    .B(net6),
    .Z(\V2/V3/v3 [4]));
 OR2_X1 \V2/V3/V3/A3/M1/_0_  (.A1(\V2/V3/V3/A3/M1/c1 ),
    .A2(\V2/V3/V3/A3/M1/c2 ),
    .ZN(\V2/V3/V3/A3/c1 ));
 AND2_X1 \V2/V3/V3/A3/M2/M1/_0_  (.A1(\V2/V3/V3/v4 [1]),
    .A2(\V2/V3/V3/s2 [3]),
    .ZN(\V2/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M2/M1/_1_  (.A(\V2/V3/V3/v4 [1]),
    .B(\V2/V3/V3/s2 [3]),
    .Z(\V2/V3/V3/A3/M2/s1 ));
 AND2_X1 \V2/V3/V3/A3/M2/M2/_0_  (.A1(\V2/V3/V3/A3/M2/s1 ),
    .A2(\V2/V3/V3/A3/c1 ),
    .ZN(\V2/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M2/M2/_1_  (.A(\V2/V3/V3/A3/M2/s1 ),
    .B(\V2/V3/V3/A3/c1 ),
    .Z(\V2/V3/v3 [5]));
 OR2_X1 \V2/V3/V3/A3/M2/_0_  (.A1(\V2/V3/V3/A3/M2/c1 ),
    .A2(\V2/V3/V3/A3/M2/c2 ),
    .ZN(\V2/V3/V3/A3/c2 ));
 AND2_X1 \V2/V3/V3/A3/M3/M1/_0_  (.A1(\V2/V3/V3/v4 [2]),
    .A2(\V2/V3/V3/c3 ),
    .ZN(\V2/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M3/M1/_1_  (.A(\V2/V3/V3/v4 [2]),
    .B(\V2/V3/V3/c3 ),
    .Z(\V2/V3/V3/A3/M3/s1 ));
 AND2_X1 \V2/V3/V3/A3/M3/M2/_0_  (.A1(\V2/V3/V3/A3/M3/s1 ),
    .A2(\V2/V3/V3/A3/c2 ),
    .ZN(\V2/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M3/M2/_1_  (.A(\V2/V3/V3/A3/M3/s1 ),
    .B(\V2/V3/V3/A3/c2 ),
    .Z(\V2/V3/v3 [6]));
 OR2_X1 \V2/V3/V3/A3/M3/_0_  (.A1(\V2/V3/V3/A3/M3/c1 ),
    .A2(\V2/V3/V3/A3/M3/c2 ),
    .ZN(\V2/V3/V3/A3/c3 ));
 AND2_X1 \V2/V3/V3/A3/M4/M1/_0_  (.A1(\V2/V3/V3/v4 [3]),
    .A2(net6),
    .ZN(\V2/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V3/A3/M4/M1/_1_  (.A(\V2/V3/V3/v4 [3]),
    .B(net6),
    .Z(\V2/V3/V3/A3/M4/s1 ));
 AND2_X1 \V2/V3/V3/A3/M4/M2/_0_  (.A1(\V2/V3/V3/A3/M4/s1 ),
    .A2(\V2/V3/V3/A3/c3 ),
    .ZN(\V2/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V3/A3/M4/M2/_1_  (.A(\V2/V3/V3/A3/M4/s1 ),
    .B(\V2/V3/V3/A3/c3 ),
    .Z(\V2/V3/v3 [7]));
 OR2_X1 \V2/V3/V3/A3/M4/_0_  (.A1(\V2/V3/V3/A3/M4/c1 ),
    .A2(\V2/V3/V3/A3/M4/c2 ),
    .ZN(\V2/V3/V3/overflow ));
 AND2_X1 \V2/V3/V3/V1/HA1/_0_  (.A1(\V2/V3/V3/V1/w2 ),
    .A2(\V2/V3/V3/V1/w1 ),
    .ZN(\V2/V3/V3/V1/w4 ));
 XOR2_X2 \V2/V3/V3/V1/HA1/_1_  (.A(\V2/V3/V3/V1/w2 ),
    .B(\V2/V3/V3/V1/w1 ),
    .Z(\V2/V3/v3 [1]));
 AND2_X1 \V2/V3/V3/V1/HA2/_0_  (.A1(\V2/V3/V3/V1/w4 ),
    .A2(\V2/V3/V3/V1/w3 ),
    .ZN(\V2/V3/V3/v1 [3]));
 XOR2_X2 \V2/V3/V3/V1/HA2/_1_  (.A(\V2/V3/V3/V1/w4 ),
    .B(\V2/V3/V3/V1/w3 ),
    .Z(\V2/V3/V3/v1 [2]));
 AND2_X1 \V2/V3/V3/V1/_0_  (.A1(net41),
    .A2(B[12]),
    .ZN(\V2/V3/v3 [0]));
 AND2_X1 \V2/V3/V3/V1/_1_  (.A1(net41),
    .A2(B[13]),
    .ZN(\V2/V3/V3/V1/w1 ));
 AND2_X1 \V2/V3/V3/V1/_2_  (.A1(B[12]),
    .A2(net40),
    .ZN(\V2/V3/V3/V1/w2 ));
 AND2_X1 \V2/V3/V3/V1/_3_  (.A1(B[13]),
    .A2(net40),
    .ZN(\V2/V3/V3/V1/w3 ));
 AND2_X1 \V2/V3/V3/V2/HA1/_0_  (.A1(\V2/V3/V3/V2/w2 ),
    .A2(\V2/V3/V3/V2/w1 ),
    .ZN(\V2/V3/V3/V2/w4 ));
 XOR2_X2 \V2/V3/V3/V2/HA1/_1_  (.A(\V2/V3/V3/V2/w2 ),
    .B(\V2/V3/V3/V2/w1 ),
    .Z(\V2/V3/V3/v2 [1]));
 AND2_X1 \V2/V3/V3/V2/HA2/_0_  (.A1(\V2/V3/V3/V2/w4 ),
    .A2(\V2/V3/V3/V2/w3 ),
    .ZN(\V2/V3/V3/v2 [3]));
 XOR2_X2 \V2/V3/V3/V2/HA2/_1_  (.A(\V2/V3/V3/V2/w4 ),
    .B(\V2/V3/V3/V2/w3 ),
    .Z(\V2/V3/V3/v2 [2]));
 AND2_X1 \V2/V3/V3/V2/_0_  (.A1(net39),
    .A2(B[12]),
    .ZN(\V2/V3/V3/v2 [0]));
 AND2_X1 \V2/V3/V3/V2/_1_  (.A1(net39),
    .A2(B[13]),
    .ZN(\V2/V3/V3/V2/w1 ));
 AND2_X1 \V2/V3/V3/V2/_2_  (.A1(B[12]),
    .A2(net38),
    .ZN(\V2/V3/V3/V2/w2 ));
 AND2_X1 \V2/V3/V3/V2/_3_  (.A1(B[13]),
    .A2(net38),
    .ZN(\V2/V3/V3/V2/w3 ));
 AND2_X1 \V2/V3/V3/V3/HA1/_0_  (.A1(\V2/V3/V3/V3/w2 ),
    .A2(\V2/V3/V3/V3/w1 ),
    .ZN(\V2/V3/V3/V3/w4 ));
 XOR2_X2 \V2/V3/V3/V3/HA1/_1_  (.A(\V2/V3/V3/V3/w2 ),
    .B(\V2/V3/V3/V3/w1 ),
    .Z(\V2/V3/V3/v3 [1]));
 AND2_X1 \V2/V3/V3/V3/HA2/_0_  (.A1(\V2/V3/V3/V3/w4 ),
    .A2(\V2/V3/V3/V3/w3 ),
    .ZN(\V2/V3/V3/v3 [3]));
 XOR2_X2 \V2/V3/V3/V3/HA2/_1_  (.A(\V2/V3/V3/V3/w4 ),
    .B(\V2/V3/V3/V3/w3 ),
    .Z(\V2/V3/V3/v3 [2]));
 AND2_X1 \V2/V3/V3/V3/_0_  (.A1(net41),
    .A2(B[14]),
    .ZN(\V2/V3/V3/v3 [0]));
 AND2_X1 \V2/V3/V3/V3/_1_  (.A1(net41),
    .A2(B[15]),
    .ZN(\V2/V3/V3/V3/w1 ));
 AND2_X1 \V2/V3/V3/V3/_2_  (.A1(B[14]),
    .A2(net40),
    .ZN(\V2/V3/V3/V3/w2 ));
 AND2_X1 \V2/V3/V3/V3/_3_  (.A1(B[15]),
    .A2(net40),
    .ZN(\V2/V3/V3/V3/w3 ));
 AND2_X1 \V2/V3/V3/V4/HA1/_0_  (.A1(\V2/V3/V3/V4/w2 ),
    .A2(\V2/V3/V3/V4/w1 ),
    .ZN(\V2/V3/V3/V4/w4 ));
 XOR2_X2 \V2/V3/V3/V4/HA1/_1_  (.A(\V2/V3/V3/V4/w2 ),
    .B(\V2/V3/V3/V4/w1 ),
    .Z(\V2/V3/V3/v4 [1]));
 AND2_X1 \V2/V3/V3/V4/HA2/_0_  (.A1(\V2/V3/V3/V4/w4 ),
    .A2(\V2/V3/V3/V4/w3 ),
    .ZN(\V2/V3/V3/v4 [3]));
 XOR2_X2 \V2/V3/V3/V4/HA2/_1_  (.A(\V2/V3/V3/V4/w4 ),
    .B(\V2/V3/V3/V4/w3 ),
    .Z(\V2/V3/V3/v4 [2]));
 AND2_X1 \V2/V3/V3/V4/_0_  (.A1(net39),
    .A2(B[14]),
    .ZN(\V2/V3/V3/v4 [0]));
 AND2_X1 \V2/V3/V3/V4/_1_  (.A1(net39),
    .A2(B[15]),
    .ZN(\V2/V3/V3/V4/w1 ));
 AND2_X1 \V2/V3/V3/V4/_2_  (.A1(B[14]),
    .A2(net38),
    .ZN(\V2/V3/V3/V4/w2 ));
 AND2_X1 \V2/V3/V3/V4/_3_  (.A1(B[15]),
    .A2(net38),
    .ZN(\V2/V3/V3/V4/w3 ));
 OR2_X1 \V2/V3/V3/_0_  (.A1(\V2/V3/V3/c1 ),
    .A2(\V2/V3/V3/c2 ),
    .ZN(\V2/V3/V3/c3 ));
 AND2_X1 \V2/V3/V4/A1/M1/M1/_0_  (.A1(\V2/V3/V4/v2 [0]),
    .A2(\V2/V3/V4/v3 [0]),
    .ZN(\V2/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M1/M1/_1_  (.A(\V2/V3/V4/v2 [0]),
    .B(\V2/V3/V4/v3 [0]),
    .Z(\V2/V3/V4/A1/M1/s1 ));
 AND2_X1 \V2/V3/V4/A1/M1/M2/_0_  (.A1(\V2/V3/V4/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V2/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M1/M2/_1_  (.A(\V2/V3/V4/A1/M1/s1 ),
    .B(net6),
    .Z(\V2/V3/V4/s1 [0]));
 OR2_X1 \V2/V3/V4/A1/M1/_0_  (.A1(\V2/V3/V4/A1/M1/c1 ),
    .A2(\V2/V3/V4/A1/M1/c2 ),
    .ZN(\V2/V3/V4/A1/c1 ));
 AND2_X1 \V2/V3/V4/A1/M2/M1/_0_  (.A1(\V2/V3/V4/v2 [1]),
    .A2(\V2/V3/V4/v3 [1]),
    .ZN(\V2/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M2/M1/_1_  (.A(\V2/V3/V4/v2 [1]),
    .B(\V2/V3/V4/v3 [1]),
    .Z(\V2/V3/V4/A1/M2/s1 ));
 AND2_X1 \V2/V3/V4/A1/M2/M2/_0_  (.A1(\V2/V3/V4/A1/M2/s1 ),
    .A2(\V2/V3/V4/A1/c1 ),
    .ZN(\V2/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M2/M2/_1_  (.A(\V2/V3/V4/A1/M2/s1 ),
    .B(\V2/V3/V4/A1/c1 ),
    .Z(\V2/V3/V4/s1 [1]));
 OR2_X1 \V2/V3/V4/A1/M2/_0_  (.A1(\V2/V3/V4/A1/M2/c1 ),
    .A2(\V2/V3/V4/A1/M2/c2 ),
    .ZN(\V2/V3/V4/A1/c2 ));
 AND2_X1 \V2/V3/V4/A1/M3/M1/_0_  (.A1(\V2/V3/V4/v2 [2]),
    .A2(\V2/V3/V4/v3 [2]),
    .ZN(\V2/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M3/M1/_1_  (.A(\V2/V3/V4/v2 [2]),
    .B(\V2/V3/V4/v3 [2]),
    .Z(\V2/V3/V4/A1/M3/s1 ));
 AND2_X1 \V2/V3/V4/A1/M3/M2/_0_  (.A1(\V2/V3/V4/A1/M3/s1 ),
    .A2(\V2/V3/V4/A1/c2 ),
    .ZN(\V2/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M3/M2/_1_  (.A(\V2/V3/V4/A1/M3/s1 ),
    .B(\V2/V3/V4/A1/c2 ),
    .Z(\V2/V3/V4/s1 [2]));
 OR2_X1 \V2/V3/V4/A1/M3/_0_  (.A1(\V2/V3/V4/A1/M3/c1 ),
    .A2(\V2/V3/V4/A1/M3/c2 ),
    .ZN(\V2/V3/V4/A1/c3 ));
 AND2_X1 \V2/V3/V4/A1/M4/M1/_0_  (.A1(\V2/V3/V4/v2 [3]),
    .A2(\V2/V3/V4/v3 [3]),
    .ZN(\V2/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A1/M4/M1/_1_  (.A(\V2/V3/V4/v2 [3]),
    .B(\V2/V3/V4/v3 [3]),
    .Z(\V2/V3/V4/A1/M4/s1 ));
 AND2_X1 \V2/V3/V4/A1/M4/M2/_0_  (.A1(\V2/V3/V4/A1/M4/s1 ),
    .A2(\V2/V3/V4/A1/c3 ),
    .ZN(\V2/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A1/M4/M2/_1_  (.A(\V2/V3/V4/A1/M4/s1 ),
    .B(\V2/V3/V4/A1/c3 ),
    .Z(\V2/V3/V4/s1 [3]));
 OR2_X1 \V2/V3/V4/A1/M4/_0_  (.A1(\V2/V3/V4/A1/M4/c1 ),
    .A2(\V2/V3/V4/A1/M4/c2 ),
    .ZN(\V2/V3/V4/c1 ));
 AND2_X1 \V2/V3/V4/A2/M1/M1/_0_  (.A1(\V2/V3/V4/s1 [0]),
    .A2(\V2/V3/V4/v1 [2]),
    .ZN(\V2/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M1/M1/_1_  (.A(\V2/V3/V4/s1 [0]),
    .B(\V2/V3/V4/v1 [2]),
    .Z(\V2/V3/V4/A2/M1/s1 ));
 AND2_X1 \V2/V3/V4/A2/M1/M2/_0_  (.A1(\V2/V3/V4/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M1/M2/_1_  (.A(\V2/V3/V4/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/v4 [2]));
 OR2_X1 \V2/V3/V4/A2/M1/_0_  (.A1(\V2/V3/V4/A2/M1/c1 ),
    .A2(\V2/V3/V4/A2/M1/c2 ),
    .ZN(\V2/V3/V4/A2/c1 ));
 AND2_X1 \V2/V3/V4/A2/M2/M1/_0_  (.A1(\V2/V3/V4/s1 [1]),
    .A2(\V2/V3/V4/v1 [3]),
    .ZN(\V2/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M2/M1/_1_  (.A(\V2/V3/V4/s1 [1]),
    .B(\V2/V3/V4/v1 [3]),
    .Z(\V2/V3/V4/A2/M2/s1 ));
 AND2_X1 \V2/V3/V4/A2/M2/M2/_0_  (.A1(\V2/V3/V4/A2/M2/s1 ),
    .A2(\V2/V3/V4/A2/c1 ),
    .ZN(\V2/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M2/M2/_1_  (.A(\V2/V3/V4/A2/M2/s1 ),
    .B(\V2/V3/V4/A2/c1 ),
    .Z(\V2/V3/v4 [3]));
 OR2_X1 \V2/V3/V4/A2/M2/_0_  (.A1(\V2/V3/V4/A2/M2/c1 ),
    .A2(\V2/V3/V4/A2/M2/c2 ),
    .ZN(\V2/V3/V4/A2/c2 ));
 AND2_X1 \V2/V3/V4/A2/M3/M1/_0_  (.A1(\V2/V3/V4/s1 [2]),
    .A2(net6),
    .ZN(\V2/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M3/M1/_1_  (.A(\V2/V3/V4/s1 [2]),
    .B(net6),
    .Z(\V2/V3/V4/A2/M3/s1 ));
 AND2_X1 \V2/V3/V4/A2/M3/M2/_0_  (.A1(\V2/V3/V4/A2/M3/s1 ),
    .A2(\V2/V3/V4/A2/c2 ),
    .ZN(\V2/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M3/M2/_1_  (.A(\V2/V3/V4/A2/M3/s1 ),
    .B(\V2/V3/V4/A2/c2 ),
    .Z(\V2/V3/V4/s2 [2]));
 OR2_X1 \V2/V3/V4/A2/M3/_0_  (.A1(\V2/V3/V4/A2/M3/c1 ),
    .A2(\V2/V3/V4/A2/M3/c2 ),
    .ZN(\V2/V3/V4/A2/c3 ));
 AND2_X1 \V2/V3/V4/A2/M4/M1/_0_  (.A1(\V2/V3/V4/s1 [3]),
    .A2(net6),
    .ZN(\V2/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A2/M4/M1/_1_  (.A(\V2/V3/V4/s1 [3]),
    .B(net6),
    .Z(\V2/V3/V4/A2/M4/s1 ));
 AND2_X1 \V2/V3/V4/A2/M4/M2/_0_  (.A1(\V2/V3/V4/A2/M4/s1 ),
    .A2(\V2/V3/V4/A2/c3 ),
    .ZN(\V2/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A2/M4/M2/_1_  (.A(\V2/V3/V4/A2/M4/s1 ),
    .B(\V2/V3/V4/A2/c3 ),
    .Z(\V2/V3/V4/s2 [3]));
 OR2_X1 \V2/V3/V4/A2/M4/_0_  (.A1(\V2/V3/V4/A2/M4/c1 ),
    .A2(\V2/V3/V4/A2/M4/c2 ),
    .ZN(\V2/V3/V4/c2 ));
 AND2_X1 \V2/V3/V4/A3/M1/M1/_0_  (.A1(\V2/V3/V4/v4 [0]),
    .A2(\V2/V3/V4/s2 [2]),
    .ZN(\V2/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M1/M1/_1_  (.A(\V2/V3/V4/v4 [0]),
    .B(\V2/V3/V4/s2 [2]),
    .Z(\V2/V3/V4/A3/M1/s1 ));
 AND2_X1 \V2/V3/V4/A3/M1/M2/_0_  (.A1(\V2/V3/V4/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M1/M2/_1_  (.A(\V2/V3/V4/A3/M1/s1 ),
    .B(net7),
    .Z(\V2/V3/v4 [4]));
 OR2_X1 \V2/V3/V4/A3/M1/_0_  (.A1(\V2/V3/V4/A3/M1/c1 ),
    .A2(\V2/V3/V4/A3/M1/c2 ),
    .ZN(\V2/V3/V4/A3/c1 ));
 AND2_X1 \V2/V3/V4/A3/M2/M1/_0_  (.A1(\V2/V3/V4/v4 [1]),
    .A2(\V2/V3/V4/s2 [3]),
    .ZN(\V2/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M2/M1/_1_  (.A(\V2/V3/V4/v4 [1]),
    .B(\V2/V3/V4/s2 [3]),
    .Z(\V2/V3/V4/A3/M2/s1 ));
 AND2_X1 \V2/V3/V4/A3/M2/M2/_0_  (.A1(\V2/V3/V4/A3/M2/s1 ),
    .A2(\V2/V3/V4/A3/c1 ),
    .ZN(\V2/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M2/M2/_1_  (.A(\V2/V3/V4/A3/M2/s1 ),
    .B(\V2/V3/V4/A3/c1 ),
    .Z(\V2/V3/v4 [5]));
 OR2_X1 \V2/V3/V4/A3/M2/_0_  (.A1(\V2/V3/V4/A3/M2/c1 ),
    .A2(\V2/V3/V4/A3/M2/c2 ),
    .ZN(\V2/V3/V4/A3/c2 ));
 AND2_X1 \V2/V3/V4/A3/M3/M1/_0_  (.A1(\V2/V3/V4/v4 [2]),
    .A2(\V2/V3/V4/c3 ),
    .ZN(\V2/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M3/M1/_1_  (.A(\V2/V3/V4/v4 [2]),
    .B(\V2/V3/V4/c3 ),
    .Z(\V2/V3/V4/A3/M3/s1 ));
 AND2_X1 \V2/V3/V4/A3/M3/M2/_0_  (.A1(\V2/V3/V4/A3/M3/s1 ),
    .A2(\V2/V3/V4/A3/c2 ),
    .ZN(\V2/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M3/M2/_1_  (.A(\V2/V3/V4/A3/M3/s1 ),
    .B(\V2/V3/V4/A3/c2 ),
    .Z(\V2/V3/v4 [6]));
 OR2_X1 \V2/V3/V4/A3/M3/_0_  (.A1(\V2/V3/V4/A3/M3/c1 ),
    .A2(\V2/V3/V4/A3/M3/c2 ),
    .ZN(\V2/V3/V4/A3/c3 ));
 AND2_X1 \V2/V3/V4/A3/M4/M1/_0_  (.A1(\V2/V3/V4/v4 [3]),
    .A2(net7),
    .ZN(\V2/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V3/V4/A3/M4/M1/_1_  (.A(\V2/V3/V4/v4 [3]),
    .B(net7),
    .Z(\V2/V3/V4/A3/M4/s1 ));
 AND2_X1 \V2/V3/V4/A3/M4/M2/_0_  (.A1(\V2/V3/V4/A3/M4/s1 ),
    .A2(\V2/V3/V4/A3/c3 ),
    .ZN(\V2/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V3/V4/A3/M4/M2/_1_  (.A(\V2/V3/V4/A3/M4/s1 ),
    .B(\V2/V3/V4/A3/c3 ),
    .Z(\V2/V3/v4 [7]));
 OR2_X1 \V2/V3/V4/A3/M4/_0_  (.A1(\V2/V3/V4/A3/M4/c1 ),
    .A2(\V2/V3/V4/A3/M4/c2 ),
    .ZN(\V2/V3/V4/overflow ));
 AND2_X1 \V2/V3/V4/V1/HA1/_0_  (.A1(\V2/V3/V4/V1/w2 ),
    .A2(\V2/V3/V4/V1/w1 ),
    .ZN(\V2/V3/V4/V1/w4 ));
 XOR2_X2 \V2/V3/V4/V1/HA1/_1_  (.A(\V2/V3/V4/V1/w2 ),
    .B(\V2/V3/V4/V1/w1 ),
    .Z(\V2/V3/v4 [1]));
 AND2_X1 \V2/V3/V4/V1/HA2/_0_  (.A1(\V2/V3/V4/V1/w4 ),
    .A2(\V2/V3/V4/V1/w3 ),
    .ZN(\V2/V3/V4/v1 [3]));
 XOR2_X2 \V2/V3/V4/V1/HA2/_1_  (.A(\V2/V3/V4/V1/w4 ),
    .B(\V2/V3/V4/V1/w3 ),
    .Z(\V2/V3/V4/v1 [2]));
 AND2_X1 \V2/V3/V4/V1/_0_  (.A1(net37),
    .A2(B[12]),
    .ZN(\V2/V3/v4 [0]));
 AND2_X1 \V2/V3/V4/V1/_1_  (.A1(net37),
    .A2(B[13]),
    .ZN(\V2/V3/V4/V1/w1 ));
 AND2_X1 \V2/V3/V4/V1/_2_  (.A1(B[12]),
    .A2(net36),
    .ZN(\V2/V3/V4/V1/w2 ));
 AND2_X1 \V2/V3/V4/V1/_3_  (.A1(B[13]),
    .A2(net36),
    .ZN(\V2/V3/V4/V1/w3 ));
 AND2_X1 \V2/V3/V4/V2/HA1/_0_  (.A1(\V2/V3/V4/V2/w2 ),
    .A2(\V2/V3/V4/V2/w1 ),
    .ZN(\V2/V3/V4/V2/w4 ));
 XOR2_X2 \V2/V3/V4/V2/HA1/_1_  (.A(\V2/V3/V4/V2/w2 ),
    .B(\V2/V3/V4/V2/w1 ),
    .Z(\V2/V3/V4/v2 [1]));
 AND2_X1 \V2/V3/V4/V2/HA2/_0_  (.A1(\V2/V3/V4/V2/w4 ),
    .A2(\V2/V3/V4/V2/w3 ),
    .ZN(\V2/V3/V4/v2 [3]));
 XOR2_X2 \V2/V3/V4/V2/HA2/_1_  (.A(\V2/V3/V4/V2/w4 ),
    .B(\V2/V3/V4/V2/w3 ),
    .Z(\V2/V3/V4/v2 [2]));
 AND2_X1 \V2/V3/V4/V2/_0_  (.A1(net35),
    .A2(B[12]),
    .ZN(\V2/V3/V4/v2 [0]));
 AND2_X1 \V2/V3/V4/V2/_1_  (.A1(net35),
    .A2(B[13]),
    .ZN(\V2/V3/V4/V2/w1 ));
 AND2_X1 \V2/V3/V4/V2/_2_  (.A1(B[12]),
    .A2(net34),
    .ZN(\V2/V3/V4/V2/w2 ));
 AND2_X1 \V2/V3/V4/V2/_3_  (.A1(B[13]),
    .A2(net34),
    .ZN(\V2/V3/V4/V2/w3 ));
 AND2_X1 \V2/V3/V4/V3/HA1/_0_  (.A1(\V2/V3/V4/V3/w2 ),
    .A2(\V2/V3/V4/V3/w1 ),
    .ZN(\V2/V3/V4/V3/w4 ));
 XOR2_X2 \V2/V3/V4/V3/HA1/_1_  (.A(\V2/V3/V4/V3/w2 ),
    .B(\V2/V3/V4/V3/w1 ),
    .Z(\V2/V3/V4/v3 [1]));
 AND2_X1 \V2/V3/V4/V3/HA2/_0_  (.A1(\V2/V3/V4/V3/w4 ),
    .A2(\V2/V3/V4/V3/w3 ),
    .ZN(\V2/V3/V4/v3 [3]));
 XOR2_X2 \V2/V3/V4/V3/HA2/_1_  (.A(\V2/V3/V4/V3/w4 ),
    .B(\V2/V3/V4/V3/w3 ),
    .Z(\V2/V3/V4/v3 [2]));
 AND2_X1 \V2/V3/V4/V3/_0_  (.A1(net37),
    .A2(B[14]),
    .ZN(\V2/V3/V4/v3 [0]));
 AND2_X1 \V2/V3/V4/V3/_1_  (.A1(net37),
    .A2(B[15]),
    .ZN(\V2/V3/V4/V3/w1 ));
 AND2_X1 \V2/V3/V4/V3/_2_  (.A1(B[14]),
    .A2(net36),
    .ZN(\V2/V3/V4/V3/w2 ));
 AND2_X1 \V2/V3/V4/V3/_3_  (.A1(B[15]),
    .A2(net36),
    .ZN(\V2/V3/V4/V3/w3 ));
 AND2_X1 \V2/V3/V4/V4/HA1/_0_  (.A1(\V2/V3/V4/V4/w2 ),
    .A2(\V2/V3/V4/V4/w1 ),
    .ZN(\V2/V3/V4/V4/w4 ));
 XOR2_X2 \V2/V3/V4/V4/HA1/_1_  (.A(\V2/V3/V4/V4/w2 ),
    .B(\V2/V3/V4/V4/w1 ),
    .Z(\V2/V3/V4/v4 [1]));
 AND2_X1 \V2/V3/V4/V4/HA2/_0_  (.A1(\V2/V3/V4/V4/w4 ),
    .A2(\V2/V3/V4/V4/w3 ),
    .ZN(\V2/V3/V4/v4 [3]));
 XOR2_X2 \V2/V3/V4/V4/HA2/_1_  (.A(\V2/V3/V4/V4/w4 ),
    .B(\V2/V3/V4/V4/w3 ),
    .Z(\V2/V3/V4/v4 [2]));
 AND2_X1 \V2/V3/V4/V4/_0_  (.A1(net35),
    .A2(B[14]),
    .ZN(\V2/V3/V4/v4 [0]));
 AND2_X1 \V2/V3/V4/V4/_1_  (.A1(net35),
    .A2(B[15]),
    .ZN(\V2/V3/V4/V4/w1 ));
 AND2_X1 \V2/V3/V4/V4/_2_  (.A1(B[14]),
    .A2(net34),
    .ZN(\V2/V3/V4/V4/w2 ));
 AND2_X1 \V2/V3/V4/V4/_3_  (.A1(B[15]),
    .A2(net34),
    .ZN(\V2/V3/V4/V4/w3 ));
 OR2_X1 \V2/V3/V4/_0_  (.A1(\V2/V3/V4/c1 ),
    .A2(\V2/V3/V4/c2 ),
    .ZN(\V2/V3/V4/c3 ));
 OR2_X1 \V2/V3/_0_  (.A1(\V2/V3/c1 ),
    .A2(\V2/V3/c2 ),
    .ZN(\V2/V3/c3 ));
 AND2_X1 \V2/V4/A1/A1/M1/M1/_0_  (.A1(\V2/V4/v2 [0]),
    .A2(\V2/V4/v3 [0]),
    .ZN(\V2/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M1/M1/_1_  (.A(\V2/V4/v2 [0]),
    .B(\V2/V4/v3 [0]),
    .Z(\V2/V4/A1/A1/M1/s1 ));
 AND2_X1 \V2/V4/A1/A1/M1/M2/_0_  (.A1(\V2/V4/A1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M1/M2/_1_  (.A(\V2/V4/A1/A1/M1/s1 ),
    .B(net9),
    .Z(\V2/V4/s1 [0]));
 OR2_X1 \V2/V4/A1/A1/M1/_0_  (.A1(\V2/V4/A1/A1/M1/c1 ),
    .A2(\V2/V4/A1/A1/M1/c2 ),
    .ZN(\V2/V4/A1/A1/c1 ));
 AND2_X1 \V2/V4/A1/A1/M2/M1/_0_  (.A1(\V2/V4/v2 [1]),
    .A2(\V2/V4/v3 [1]),
    .ZN(\V2/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M2/M1/_1_  (.A(\V2/V4/v2 [1]),
    .B(\V2/V4/v3 [1]),
    .Z(\V2/V4/A1/A1/M2/s1 ));
 AND2_X1 \V2/V4/A1/A1/M2/M2/_0_  (.A1(\V2/V4/A1/A1/M2/s1 ),
    .A2(\V2/V4/A1/A1/c1 ),
    .ZN(\V2/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M2/M2/_1_  (.A(\V2/V4/A1/A1/M2/s1 ),
    .B(\V2/V4/A1/A1/c1 ),
    .Z(\V2/V4/s1 [1]));
 OR2_X1 \V2/V4/A1/A1/M2/_0_  (.A1(\V2/V4/A1/A1/M2/c1 ),
    .A2(\V2/V4/A1/A1/M2/c2 ),
    .ZN(\V2/V4/A1/A1/c2 ));
 AND2_X1 \V2/V4/A1/A1/M3/M1/_0_  (.A1(\V2/V4/v2 [2]),
    .A2(\V2/V4/v3 [2]),
    .ZN(\V2/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M3/M1/_1_  (.A(\V2/V4/v2 [2]),
    .B(\V2/V4/v3 [2]),
    .Z(\V2/V4/A1/A1/M3/s1 ));
 AND2_X1 \V2/V4/A1/A1/M3/M2/_0_  (.A1(\V2/V4/A1/A1/M3/s1 ),
    .A2(\V2/V4/A1/A1/c2 ),
    .ZN(\V2/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M3/M2/_1_  (.A(\V2/V4/A1/A1/M3/s1 ),
    .B(\V2/V4/A1/A1/c2 ),
    .Z(\V2/V4/s1 [2]));
 OR2_X1 \V2/V4/A1/A1/M3/_0_  (.A1(\V2/V4/A1/A1/M3/c1 ),
    .A2(\V2/V4/A1/A1/M3/c2 ),
    .ZN(\V2/V4/A1/A1/c3 ));
 AND2_X1 \V2/V4/A1/A1/M4/M1/_0_  (.A1(\V2/V4/v2 [3]),
    .A2(\V2/V4/v3 [3]),
    .ZN(\V2/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A1/A1/M4/M1/_1_  (.A(\V2/V4/v2 [3]),
    .B(\V2/V4/v3 [3]),
    .Z(\V2/V4/A1/A1/M4/s1 ));
 AND2_X1 \V2/V4/A1/A1/M4/M2/_0_  (.A1(\V2/V4/A1/A1/M4/s1 ),
    .A2(\V2/V4/A1/A1/c3 ),
    .ZN(\V2/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A1/A1/M4/M2/_1_  (.A(\V2/V4/A1/A1/M4/s1 ),
    .B(\V2/V4/A1/A1/c3 ),
    .Z(\V2/V4/s1 [3]));
 OR2_X1 \V2/V4/A1/A1/M4/_0_  (.A1(\V2/V4/A1/A1/M4/c1 ),
    .A2(\V2/V4/A1/A1/M4/c2 ),
    .ZN(\V2/V4/A1/c1 ));
 AND2_X1 \V2/V4/A1/A2/M1/M1/_0_  (.A1(\V2/V4/v2 [4]),
    .A2(\V2/V4/v3 [4]),
    .ZN(\V2/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M1/M1/_1_  (.A(\V2/V4/v2 [4]),
    .B(\V2/V4/v3 [4]),
    .Z(\V2/V4/A1/A2/M1/s1 ));
 AND2_X1 \V2/V4/A1/A2/M1/M2/_0_  (.A1(\V2/V4/A1/A2/M1/s1 ),
    .A2(\V2/V4/A1/c1 ),
    .ZN(\V2/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M1/M2/_1_  (.A(\V2/V4/A1/A2/M1/s1 ),
    .B(\V2/V4/A1/c1 ),
    .Z(\V2/V4/s1 [4]));
 OR2_X1 \V2/V4/A1/A2/M1/_0_  (.A1(\V2/V4/A1/A2/M1/c1 ),
    .A2(\V2/V4/A1/A2/M1/c2 ),
    .ZN(\V2/V4/A1/A2/c1 ));
 AND2_X1 \V2/V4/A1/A2/M2/M1/_0_  (.A1(\V2/V4/v2 [5]),
    .A2(\V2/V4/v3 [5]),
    .ZN(\V2/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M2/M1/_1_  (.A(\V2/V4/v2 [5]),
    .B(\V2/V4/v3 [5]),
    .Z(\V2/V4/A1/A2/M2/s1 ));
 AND2_X1 \V2/V4/A1/A2/M2/M2/_0_  (.A1(\V2/V4/A1/A2/M2/s1 ),
    .A2(\V2/V4/A1/A2/c1 ),
    .ZN(\V2/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M2/M2/_1_  (.A(\V2/V4/A1/A2/M2/s1 ),
    .B(\V2/V4/A1/A2/c1 ),
    .Z(\V2/V4/s1 [5]));
 OR2_X1 \V2/V4/A1/A2/M2/_0_  (.A1(\V2/V4/A1/A2/M2/c1 ),
    .A2(\V2/V4/A1/A2/M2/c2 ),
    .ZN(\V2/V4/A1/A2/c2 ));
 AND2_X1 \V2/V4/A1/A2/M3/M1/_0_  (.A1(\V2/V4/v2 [6]),
    .A2(\V2/V4/v3 [6]),
    .ZN(\V2/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M3/M1/_1_  (.A(\V2/V4/v2 [6]),
    .B(\V2/V4/v3 [6]),
    .Z(\V2/V4/A1/A2/M3/s1 ));
 AND2_X1 \V2/V4/A1/A2/M3/M2/_0_  (.A1(\V2/V4/A1/A2/M3/s1 ),
    .A2(\V2/V4/A1/A2/c2 ),
    .ZN(\V2/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M3/M2/_1_  (.A(\V2/V4/A1/A2/M3/s1 ),
    .B(\V2/V4/A1/A2/c2 ),
    .Z(\V2/V4/s1 [6]));
 OR2_X1 \V2/V4/A1/A2/M3/_0_  (.A1(\V2/V4/A1/A2/M3/c1 ),
    .A2(\V2/V4/A1/A2/M3/c2 ),
    .ZN(\V2/V4/A1/A2/c3 ));
 AND2_X1 \V2/V4/A1/A2/M4/M1/_0_  (.A1(\V2/V4/v2 [7]),
    .A2(\V2/V4/v3 [7]),
    .ZN(\V2/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A1/A2/M4/M1/_1_  (.A(\V2/V4/v2 [7]),
    .B(\V2/V4/v3 [7]),
    .Z(\V2/V4/A1/A2/M4/s1 ));
 AND2_X1 \V2/V4/A1/A2/M4/M2/_0_  (.A1(\V2/V4/A1/A2/M4/s1 ),
    .A2(\V2/V4/A1/A2/c3 ),
    .ZN(\V2/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A1/A2/M4/M2/_1_  (.A(\V2/V4/A1/A2/M4/s1 ),
    .B(\V2/V4/A1/A2/c3 ),
    .Z(\V2/V4/s1 [7]));
 OR2_X1 \V2/V4/A1/A2/M4/_0_  (.A1(\V2/V4/A1/A2/M4/c1 ),
    .A2(\V2/V4/A1/A2/M4/c2 ),
    .ZN(\V2/V4/c1 ));
 AND2_X1 \V2/V4/A2/A1/M1/M1/_0_  (.A1(\V2/V4/s1 [0]),
    .A2(\V2/V4/v1 [4]),
    .ZN(\V2/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M1/M1/_1_  (.A(\V2/V4/s1 [0]),
    .B(\V2/V4/v1 [4]),
    .Z(\V2/V4/A2/A1/M1/s1 ));
 AND2_X1 \V2/V4/A2/A1/M1/M2/_0_  (.A1(\V2/V4/A2/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M1/M2/_1_  (.A(\V2/V4/A2/A1/M1/s1 ),
    .B(net9),
    .Z(\V2/v4 [4]));
 OR2_X1 \V2/V4/A2/A1/M1/_0_  (.A1(\V2/V4/A2/A1/M1/c1 ),
    .A2(\V2/V4/A2/A1/M1/c2 ),
    .ZN(\V2/V4/A2/A1/c1 ));
 AND2_X1 \V2/V4/A2/A1/M2/M1/_0_  (.A1(\V2/V4/s1 [1]),
    .A2(\V2/V4/v1 [5]),
    .ZN(\V2/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M2/M1/_1_  (.A(\V2/V4/s1 [1]),
    .B(\V2/V4/v1 [5]),
    .Z(\V2/V4/A2/A1/M2/s1 ));
 AND2_X1 \V2/V4/A2/A1/M2/M2/_0_  (.A1(\V2/V4/A2/A1/M2/s1 ),
    .A2(\V2/V4/A2/A1/c1 ),
    .ZN(\V2/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M2/M2/_1_  (.A(\V2/V4/A2/A1/M2/s1 ),
    .B(\V2/V4/A2/A1/c1 ),
    .Z(\V2/v4 [5]));
 OR2_X1 \V2/V4/A2/A1/M2/_0_  (.A1(\V2/V4/A2/A1/M2/c1 ),
    .A2(\V2/V4/A2/A1/M2/c2 ),
    .ZN(\V2/V4/A2/A1/c2 ));
 AND2_X1 \V2/V4/A2/A1/M3/M1/_0_  (.A1(\V2/V4/s1 [2]),
    .A2(\V2/V4/v1 [6]),
    .ZN(\V2/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M3/M1/_1_  (.A(\V2/V4/s1 [2]),
    .B(\V2/V4/v1 [6]),
    .Z(\V2/V4/A2/A1/M3/s1 ));
 AND2_X1 \V2/V4/A2/A1/M3/M2/_0_  (.A1(\V2/V4/A2/A1/M3/s1 ),
    .A2(\V2/V4/A2/A1/c2 ),
    .ZN(\V2/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M3/M2/_1_  (.A(\V2/V4/A2/A1/M3/s1 ),
    .B(\V2/V4/A2/A1/c2 ),
    .Z(\V2/v4 [6]));
 OR2_X1 \V2/V4/A2/A1/M3/_0_  (.A1(\V2/V4/A2/A1/M3/c1 ),
    .A2(\V2/V4/A2/A1/M3/c2 ),
    .ZN(\V2/V4/A2/A1/c3 ));
 AND2_X1 \V2/V4/A2/A1/M4/M1/_0_  (.A1(\V2/V4/s1 [3]),
    .A2(\V2/V4/v1 [7]),
    .ZN(\V2/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A2/A1/M4/M1/_1_  (.A(\V2/V4/s1 [3]),
    .B(\V2/V4/v1 [7]),
    .Z(\V2/V4/A2/A1/M4/s1 ));
 AND2_X1 \V2/V4/A2/A1/M4/M2/_0_  (.A1(\V2/V4/A2/A1/M4/s1 ),
    .A2(\V2/V4/A2/A1/c3 ),
    .ZN(\V2/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A2/A1/M4/M2/_1_  (.A(\V2/V4/A2/A1/M4/s1 ),
    .B(\V2/V4/A2/A1/c3 ),
    .Z(\V2/v4 [7]));
 OR2_X1 \V2/V4/A2/A1/M4/_0_  (.A1(\V2/V4/A2/A1/M4/c1 ),
    .A2(\V2/V4/A2/A1/M4/c2 ),
    .ZN(\V2/V4/A2/c1 ));
 AND2_X1 \V2/V4/A2/A2/M1/M1/_0_  (.A1(\V2/V4/s1 [4]),
    .A2(net7),
    .ZN(\V2/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M1/M1/_1_  (.A(\V2/V4/s1 [4]),
    .B(net7),
    .Z(\V2/V4/A2/A2/M1/s1 ));
 AND2_X1 \V2/V4/A2/A2/M1/M2/_0_  (.A1(\V2/V4/A2/A2/M1/s1 ),
    .A2(\V2/V4/A2/c1 ),
    .ZN(\V2/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M1/M2/_1_  (.A(\V2/V4/A2/A2/M1/s1 ),
    .B(\V2/V4/A2/c1 ),
    .Z(\V2/V4/s2 [4]));
 OR2_X1 \V2/V4/A2/A2/M1/_0_  (.A1(\V2/V4/A2/A2/M1/c1 ),
    .A2(\V2/V4/A2/A2/M1/c2 ),
    .ZN(\V2/V4/A2/A2/c1 ));
 AND2_X1 \V2/V4/A2/A2/M2/M1/_0_  (.A1(\V2/V4/s1 [5]),
    .A2(net7),
    .ZN(\V2/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M2/M1/_1_  (.A(\V2/V4/s1 [5]),
    .B(net7),
    .Z(\V2/V4/A2/A2/M2/s1 ));
 AND2_X1 \V2/V4/A2/A2/M2/M2/_0_  (.A1(\V2/V4/A2/A2/M2/s1 ),
    .A2(\V2/V4/A2/A2/c1 ),
    .ZN(\V2/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M2/M2/_1_  (.A(\V2/V4/A2/A2/M2/s1 ),
    .B(\V2/V4/A2/A2/c1 ),
    .Z(\V2/V4/s2 [5]));
 OR2_X1 \V2/V4/A2/A2/M2/_0_  (.A1(\V2/V4/A2/A2/M2/c1 ),
    .A2(\V2/V4/A2/A2/M2/c2 ),
    .ZN(\V2/V4/A2/A2/c2 ));
 AND2_X1 \V2/V4/A2/A2/M3/M1/_0_  (.A1(\V2/V4/s1 [6]),
    .A2(net7),
    .ZN(\V2/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M3/M1/_1_  (.A(\V2/V4/s1 [6]),
    .B(net7),
    .Z(\V2/V4/A2/A2/M3/s1 ));
 AND2_X1 \V2/V4/A2/A2/M3/M2/_0_  (.A1(\V2/V4/A2/A2/M3/s1 ),
    .A2(\V2/V4/A2/A2/c2 ),
    .ZN(\V2/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M3/M2/_1_  (.A(\V2/V4/A2/A2/M3/s1 ),
    .B(\V2/V4/A2/A2/c2 ),
    .Z(\V2/V4/s2 [6]));
 OR2_X1 \V2/V4/A2/A2/M3/_0_  (.A1(\V2/V4/A2/A2/M3/c1 ),
    .A2(\V2/V4/A2/A2/M3/c2 ),
    .ZN(\V2/V4/A2/A2/c3 ));
 AND2_X1 \V2/V4/A2/A2/M4/M1/_0_  (.A1(\V2/V4/s1 [7]),
    .A2(net7),
    .ZN(\V2/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A2/A2/M4/M1/_1_  (.A(\V2/V4/s1 [7]),
    .B(net7),
    .Z(\V2/V4/A2/A2/M4/s1 ));
 AND2_X1 \V2/V4/A2/A2/M4/M2/_0_  (.A1(\V2/V4/A2/A2/M4/s1 ),
    .A2(\V2/V4/A2/A2/c3 ),
    .ZN(\V2/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A2/A2/M4/M2/_1_  (.A(\V2/V4/A2/A2/M4/s1 ),
    .B(\V2/V4/A2/A2/c3 ),
    .Z(\V2/V4/s2 [7]));
 OR2_X1 \V2/V4/A2/A2/M4/_0_  (.A1(\V2/V4/A2/A2/M4/c1 ),
    .A2(\V2/V4/A2/A2/M4/c2 ),
    .ZN(\V2/V4/c2 ));
 AND2_X1 \V2/V4/A3/A1/M1/M1/_0_  (.A1(\V2/V4/v4 [0]),
    .A2(\V2/V4/s2 [4]),
    .ZN(\V2/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M1/M1/_1_  (.A(\V2/V4/v4 [0]),
    .B(\V2/V4/s2 [4]),
    .Z(\V2/V4/A3/A1/M1/s1 ));
 AND2_X1 \V2/V4/A3/A1/M1/M2/_0_  (.A1(\V2/V4/A3/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M1/M2/_1_  (.A(\V2/V4/A3/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/v4 [8]));
 OR2_X1 \V2/V4/A3/A1/M1/_0_  (.A1(\V2/V4/A3/A1/M1/c1 ),
    .A2(\V2/V4/A3/A1/M1/c2 ),
    .ZN(\V2/V4/A3/A1/c1 ));
 AND2_X1 \V2/V4/A3/A1/M2/M1/_0_  (.A1(\V2/V4/v4 [1]),
    .A2(\V2/V4/s2 [5]),
    .ZN(\V2/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M2/M1/_1_  (.A(\V2/V4/v4 [1]),
    .B(\V2/V4/s2 [5]),
    .Z(\V2/V4/A3/A1/M2/s1 ));
 AND2_X1 \V2/V4/A3/A1/M2/M2/_0_  (.A1(\V2/V4/A3/A1/M2/s1 ),
    .A2(\V2/V4/A3/A1/c1 ),
    .ZN(\V2/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M2/M2/_1_  (.A(\V2/V4/A3/A1/M2/s1 ),
    .B(\V2/V4/A3/A1/c1 ),
    .Z(\V2/v4 [9]));
 OR2_X1 \V2/V4/A3/A1/M2/_0_  (.A1(\V2/V4/A3/A1/M2/c1 ),
    .A2(\V2/V4/A3/A1/M2/c2 ),
    .ZN(\V2/V4/A3/A1/c2 ));
 AND2_X1 \V2/V4/A3/A1/M3/M1/_0_  (.A1(\V2/V4/v4 [2]),
    .A2(\V2/V4/s2 [6]),
    .ZN(\V2/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M3/M1/_1_  (.A(\V2/V4/v4 [2]),
    .B(\V2/V4/s2 [6]),
    .Z(\V2/V4/A3/A1/M3/s1 ));
 AND2_X1 \V2/V4/A3/A1/M3/M2/_0_  (.A1(\V2/V4/A3/A1/M3/s1 ),
    .A2(\V2/V4/A3/A1/c2 ),
    .ZN(\V2/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M3/M2/_1_  (.A(\V2/V4/A3/A1/M3/s1 ),
    .B(\V2/V4/A3/A1/c2 ),
    .Z(\V2/v4 [10]));
 OR2_X1 \V2/V4/A3/A1/M3/_0_  (.A1(\V2/V4/A3/A1/M3/c1 ),
    .A2(\V2/V4/A3/A1/M3/c2 ),
    .ZN(\V2/V4/A3/A1/c3 ));
 AND2_X1 \V2/V4/A3/A1/M4/M1/_0_  (.A1(\V2/V4/v4 [3]),
    .A2(\V2/V4/s2 [7]),
    .ZN(\V2/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V2/V4/A3/A1/M4/M1/_1_  (.A(\V2/V4/v4 [3]),
    .B(\V2/V4/s2 [7]),
    .Z(\V2/V4/A3/A1/M4/s1 ));
 AND2_X1 \V2/V4/A3/A1/M4/M2/_0_  (.A1(\V2/V4/A3/A1/M4/s1 ),
    .A2(\V2/V4/A3/A1/c3 ),
    .ZN(\V2/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V2/V4/A3/A1/M4/M2/_1_  (.A(\V2/V4/A3/A1/M4/s1 ),
    .B(\V2/V4/A3/A1/c3 ),
    .Z(\V2/v4 [11]));
 OR2_X1 \V2/V4/A3/A1/M4/_0_  (.A1(\V2/V4/A3/A1/M4/c1 ),
    .A2(\V2/V4/A3/A1/M4/c2 ),
    .ZN(\V2/V4/A3/c1 ));
 AND2_X1 \V2/V4/A3/A2/M1/M1/_0_  (.A1(\V2/V4/v4 [4]),
    .A2(\V2/V4/c3 ),
    .ZN(\V2/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M1/M1/_1_  (.A(\V2/V4/v4 [4]),
    .B(\V2/V4/c3 ),
    .Z(\V2/V4/A3/A2/M1/s1 ));
 AND2_X1 \V2/V4/A3/A2/M1/M2/_0_  (.A1(\V2/V4/A3/A2/M1/s1 ),
    .A2(\V2/V4/A3/c1 ),
    .ZN(\V2/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M1/M2/_1_  (.A(\V2/V4/A3/A2/M1/s1 ),
    .B(\V2/V4/A3/c1 ),
    .Z(\V2/v4 [12]));
 OR2_X1 \V2/V4/A3/A2/M1/_0_  (.A1(\V2/V4/A3/A2/M1/c1 ),
    .A2(\V2/V4/A3/A2/M1/c2 ),
    .ZN(\V2/V4/A3/A2/c1 ));
 AND2_X1 \V2/V4/A3/A2/M2/M1/_0_  (.A1(\V2/V4/v4 [5]),
    .A2(net6),
    .ZN(\V2/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M2/M1/_1_  (.A(\V2/V4/v4 [5]),
    .B(net6),
    .Z(\V2/V4/A3/A2/M2/s1 ));
 AND2_X1 \V2/V4/A3/A2/M2/M2/_0_  (.A1(\V2/V4/A3/A2/M2/s1 ),
    .A2(\V2/V4/A3/A2/c1 ),
    .ZN(\V2/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M2/M2/_1_  (.A(\V2/V4/A3/A2/M2/s1 ),
    .B(\V2/V4/A3/A2/c1 ),
    .Z(\V2/v4 [13]));
 OR2_X1 \V2/V4/A3/A2/M2/_0_  (.A1(\V2/V4/A3/A2/M2/c1 ),
    .A2(\V2/V4/A3/A2/M2/c2 ),
    .ZN(\V2/V4/A3/A2/c2 ));
 AND2_X1 \V2/V4/A3/A2/M3/M1/_0_  (.A1(\V2/V4/v4 [6]),
    .A2(net6),
    .ZN(\V2/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M3/M1/_1_  (.A(\V2/V4/v4 [6]),
    .B(net6),
    .Z(\V2/V4/A3/A2/M3/s1 ));
 AND2_X1 \V2/V4/A3/A2/M3/M2/_0_  (.A1(\V2/V4/A3/A2/M3/s1 ),
    .A2(\V2/V4/A3/A2/c2 ),
    .ZN(\V2/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M3/M2/_1_  (.A(\V2/V4/A3/A2/M3/s1 ),
    .B(\V2/V4/A3/A2/c2 ),
    .Z(\V2/v4 [14]));
 OR2_X1 \V2/V4/A3/A2/M3/_0_  (.A1(\V2/V4/A3/A2/M3/c1 ),
    .A2(\V2/V4/A3/A2/M3/c2 ),
    .ZN(\V2/V4/A3/A2/c3 ));
 AND2_X1 \V2/V4/A3/A2/M4/M1/_0_  (.A1(\V2/V4/v4 [7]),
    .A2(net6),
    .ZN(\V2/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V2/V4/A3/A2/M4/M1/_1_  (.A(\V2/V4/v4 [7]),
    .B(net6),
    .Z(\V2/V4/A3/A2/M4/s1 ));
 AND2_X1 \V2/V4/A3/A2/M4/M2/_0_  (.A1(\V2/V4/A3/A2/M4/s1 ),
    .A2(\V2/V4/A3/A2/c3 ),
    .ZN(\V2/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V2/V4/A3/A2/M4/M2/_1_  (.A(\V2/V4/A3/A2/M4/s1 ),
    .B(\V2/V4/A3/A2/c3 ),
    .Z(\V2/v4 [15]));
 OR2_X1 \V2/V4/A3/A2/M4/_0_  (.A1(\V2/V4/A3/A2/M4/c1 ),
    .A2(\V2/V4/A3/A2/M4/c2 ),
    .ZN(\V2/V4/overflow ));
 AND2_X1 \V2/V4/V1/A1/M1/M1/_0_  (.A1(\V2/V4/V1/v2 [0]),
    .A2(\V2/V4/V1/v3 [0]),
    .ZN(\V2/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M1/M1/_1_  (.A(\V2/V4/V1/v2 [0]),
    .B(\V2/V4/V1/v3 [0]),
    .Z(\V2/V4/V1/A1/M1/s1 ));
 AND2_X1 \V2/V4/V1/A1/M1/M2/_0_  (.A1(\V2/V4/V1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M1/M2/_1_  (.A(\V2/V4/V1/A1/M1/s1 ),
    .B(net9),
    .Z(\V2/V4/V1/s1 [0]));
 OR2_X1 \V2/V4/V1/A1/M1/_0_  (.A1(\V2/V4/V1/A1/M1/c1 ),
    .A2(\V2/V4/V1/A1/M1/c2 ),
    .ZN(\V2/V4/V1/A1/c1 ));
 AND2_X1 \V2/V4/V1/A1/M2/M1/_0_  (.A1(\V2/V4/V1/v2 [1]),
    .A2(\V2/V4/V1/v3 [1]),
    .ZN(\V2/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M2/M1/_1_  (.A(\V2/V4/V1/v2 [1]),
    .B(\V2/V4/V1/v3 [1]),
    .Z(\V2/V4/V1/A1/M2/s1 ));
 AND2_X1 \V2/V4/V1/A1/M2/M2/_0_  (.A1(\V2/V4/V1/A1/M2/s1 ),
    .A2(\V2/V4/V1/A1/c1 ),
    .ZN(\V2/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M2/M2/_1_  (.A(\V2/V4/V1/A1/M2/s1 ),
    .B(\V2/V4/V1/A1/c1 ),
    .Z(\V2/V4/V1/s1 [1]));
 OR2_X1 \V2/V4/V1/A1/M2/_0_  (.A1(\V2/V4/V1/A1/M2/c1 ),
    .A2(\V2/V4/V1/A1/M2/c2 ),
    .ZN(\V2/V4/V1/A1/c2 ));
 AND2_X1 \V2/V4/V1/A1/M3/M1/_0_  (.A1(\V2/V4/V1/v2 [2]),
    .A2(\V2/V4/V1/v3 [2]),
    .ZN(\V2/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M3/M1/_1_  (.A(\V2/V4/V1/v2 [2]),
    .B(\V2/V4/V1/v3 [2]),
    .Z(\V2/V4/V1/A1/M3/s1 ));
 AND2_X1 \V2/V4/V1/A1/M3/M2/_0_  (.A1(\V2/V4/V1/A1/M3/s1 ),
    .A2(\V2/V4/V1/A1/c2 ),
    .ZN(\V2/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M3/M2/_1_  (.A(\V2/V4/V1/A1/M3/s1 ),
    .B(\V2/V4/V1/A1/c2 ),
    .Z(\V2/V4/V1/s1 [2]));
 OR2_X1 \V2/V4/V1/A1/M3/_0_  (.A1(\V2/V4/V1/A1/M3/c1 ),
    .A2(\V2/V4/V1/A1/M3/c2 ),
    .ZN(\V2/V4/V1/A1/c3 ));
 AND2_X1 \V2/V4/V1/A1/M4/M1/_0_  (.A1(\V2/V4/V1/v2 [3]),
    .A2(\V2/V4/V1/v3 [3]),
    .ZN(\V2/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A1/M4/M1/_1_  (.A(\V2/V4/V1/v2 [3]),
    .B(\V2/V4/V1/v3 [3]),
    .Z(\V2/V4/V1/A1/M4/s1 ));
 AND2_X1 \V2/V4/V1/A1/M4/M2/_0_  (.A1(\V2/V4/V1/A1/M4/s1 ),
    .A2(\V2/V4/V1/A1/c3 ),
    .ZN(\V2/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A1/M4/M2/_1_  (.A(\V2/V4/V1/A1/M4/s1 ),
    .B(\V2/V4/V1/A1/c3 ),
    .Z(\V2/V4/V1/s1 [3]));
 OR2_X1 \V2/V4/V1/A1/M4/_0_  (.A1(\V2/V4/V1/A1/M4/c1 ),
    .A2(\V2/V4/V1/A1/M4/c2 ),
    .ZN(\V2/V4/V1/c1 ));
 AND2_X1 \V2/V4/V1/A2/M1/M1/_0_  (.A1(\V2/V4/V1/s1 [0]),
    .A2(\V2/V4/V1/v1 [2]),
    .ZN(\V2/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M1/M1/_1_  (.A(\V2/V4/V1/s1 [0]),
    .B(\V2/V4/V1/v1 [2]),
    .Z(\V2/V4/V1/A2/M1/s1 ));
 AND2_X1 \V2/V4/V1/A2/M1/M2/_0_  (.A1(\V2/V4/V1/A2/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M1/M2/_1_  (.A(\V2/V4/V1/A2/M1/s1 ),
    .B(net9),
    .Z(\V2/v4 [2]));
 OR2_X1 \V2/V4/V1/A2/M1/_0_  (.A1(\V2/V4/V1/A2/M1/c1 ),
    .A2(\V2/V4/V1/A2/M1/c2 ),
    .ZN(\V2/V4/V1/A2/c1 ));
 AND2_X1 \V2/V4/V1/A2/M2/M1/_0_  (.A1(\V2/V4/V1/s1 [1]),
    .A2(\V2/V4/V1/v1 [3]),
    .ZN(\V2/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M2/M1/_1_  (.A(\V2/V4/V1/s1 [1]),
    .B(\V2/V4/V1/v1 [3]),
    .Z(\V2/V4/V1/A2/M2/s1 ));
 AND2_X1 \V2/V4/V1/A2/M2/M2/_0_  (.A1(\V2/V4/V1/A2/M2/s1 ),
    .A2(\V2/V4/V1/A2/c1 ),
    .ZN(\V2/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M2/M2/_1_  (.A(\V2/V4/V1/A2/M2/s1 ),
    .B(\V2/V4/V1/A2/c1 ),
    .Z(\V2/v4 [3]));
 OR2_X1 \V2/V4/V1/A2/M2/_0_  (.A1(\V2/V4/V1/A2/M2/c1 ),
    .A2(\V2/V4/V1/A2/M2/c2 ),
    .ZN(\V2/V4/V1/A2/c2 ));
 AND2_X1 \V2/V4/V1/A2/M3/M1/_0_  (.A1(\V2/V4/V1/s1 [2]),
    .A2(net9),
    .ZN(\V2/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M3/M1/_1_  (.A(\V2/V4/V1/s1 [2]),
    .B(net9),
    .Z(\V2/V4/V1/A2/M3/s1 ));
 AND2_X1 \V2/V4/V1/A2/M3/M2/_0_  (.A1(\V2/V4/V1/A2/M3/s1 ),
    .A2(\V2/V4/V1/A2/c2 ),
    .ZN(\V2/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M3/M2/_1_  (.A(\V2/V4/V1/A2/M3/s1 ),
    .B(\V2/V4/V1/A2/c2 ),
    .Z(\V2/V4/V1/s2 [2]));
 OR2_X1 \V2/V4/V1/A2/M3/_0_  (.A1(\V2/V4/V1/A2/M3/c1 ),
    .A2(\V2/V4/V1/A2/M3/c2 ),
    .ZN(\V2/V4/V1/A2/c3 ));
 AND2_X1 \V2/V4/V1/A2/M4/M1/_0_  (.A1(\V2/V4/V1/s1 [3]),
    .A2(net9),
    .ZN(\V2/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A2/M4/M1/_1_  (.A(\V2/V4/V1/s1 [3]),
    .B(net9),
    .Z(\V2/V4/V1/A2/M4/s1 ));
 AND2_X1 \V2/V4/V1/A2/M4/M2/_0_  (.A1(\V2/V4/V1/A2/M4/s1 ),
    .A2(\V2/V4/V1/A2/c3 ),
    .ZN(\V2/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A2/M4/M2/_1_  (.A(\V2/V4/V1/A2/M4/s1 ),
    .B(\V2/V4/V1/A2/c3 ),
    .Z(\V2/V4/V1/s2 [3]));
 OR2_X1 \V2/V4/V1/A2/M4/_0_  (.A1(\V2/V4/V1/A2/M4/c1 ),
    .A2(\V2/V4/V1/A2/M4/c2 ),
    .ZN(\V2/V4/V1/c2 ));
 AND2_X1 \V2/V4/V1/A3/M1/M1/_0_  (.A1(\V2/V4/V1/v4 [0]),
    .A2(\V2/V4/V1/s2 [2]),
    .ZN(\V2/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M1/M1/_1_  (.A(\V2/V4/V1/v4 [0]),
    .B(\V2/V4/V1/s2 [2]),
    .Z(\V2/V4/V1/A3/M1/s1 ));
 AND2_X1 \V2/V4/V1/A3/M1/M2/_0_  (.A1(\V2/V4/V1/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M1/M2/_1_  (.A(\V2/V4/V1/A3/M1/s1 ),
    .B(net9),
    .Z(\V2/V4/v1 [4]));
 OR2_X1 \V2/V4/V1/A3/M1/_0_  (.A1(\V2/V4/V1/A3/M1/c1 ),
    .A2(\V2/V4/V1/A3/M1/c2 ),
    .ZN(\V2/V4/V1/A3/c1 ));
 AND2_X1 \V2/V4/V1/A3/M2/M1/_0_  (.A1(\V2/V4/V1/v4 [1]),
    .A2(\V2/V4/V1/s2 [3]),
    .ZN(\V2/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M2/M1/_1_  (.A(\V2/V4/V1/v4 [1]),
    .B(\V2/V4/V1/s2 [3]),
    .Z(\V2/V4/V1/A3/M2/s1 ));
 AND2_X1 \V2/V4/V1/A3/M2/M2/_0_  (.A1(\V2/V4/V1/A3/M2/s1 ),
    .A2(\V2/V4/V1/A3/c1 ),
    .ZN(\V2/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M2/M2/_1_  (.A(\V2/V4/V1/A3/M2/s1 ),
    .B(\V2/V4/V1/A3/c1 ),
    .Z(\V2/V4/v1 [5]));
 OR2_X1 \V2/V4/V1/A3/M2/_0_  (.A1(\V2/V4/V1/A3/M2/c1 ),
    .A2(\V2/V4/V1/A3/M2/c2 ),
    .ZN(\V2/V4/V1/A3/c2 ));
 AND2_X1 \V2/V4/V1/A3/M3/M1/_0_  (.A1(\V2/V4/V1/v4 [2]),
    .A2(\V2/V4/V1/c3 ),
    .ZN(\V2/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M3/M1/_1_  (.A(\V2/V4/V1/v4 [2]),
    .B(\V2/V4/V1/c3 ),
    .Z(\V2/V4/V1/A3/M3/s1 ));
 AND2_X1 \V2/V4/V1/A3/M3/M2/_0_  (.A1(\V2/V4/V1/A3/M3/s1 ),
    .A2(\V2/V4/V1/A3/c2 ),
    .ZN(\V2/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M3/M2/_1_  (.A(\V2/V4/V1/A3/M3/s1 ),
    .B(\V2/V4/V1/A3/c2 ),
    .Z(\V2/V4/v1 [6]));
 OR2_X1 \V2/V4/V1/A3/M3/_0_  (.A1(\V2/V4/V1/A3/M3/c1 ),
    .A2(\V2/V4/V1/A3/M3/c2 ),
    .ZN(\V2/V4/V1/A3/c3 ));
 AND2_X1 \V2/V4/V1/A3/M4/M1/_0_  (.A1(\V2/V4/V1/v4 [3]),
    .A2(net9),
    .ZN(\V2/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V1/A3/M4/M1/_1_  (.A(\V2/V4/V1/v4 [3]),
    .B(net9),
    .Z(\V2/V4/V1/A3/M4/s1 ));
 AND2_X1 \V2/V4/V1/A3/M4/M2/_0_  (.A1(\V2/V4/V1/A3/M4/s1 ),
    .A2(\V2/V4/V1/A3/c3 ),
    .ZN(\V2/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V1/A3/M4/M2/_1_  (.A(\V2/V4/V1/A3/M4/s1 ),
    .B(\V2/V4/V1/A3/c3 ),
    .Z(\V2/V4/v1 [7]));
 OR2_X1 \V2/V4/V1/A3/M4/_0_  (.A1(\V2/V4/V1/A3/M4/c1 ),
    .A2(\V2/V4/V1/A3/M4/c2 ),
    .ZN(\V2/V4/V1/overflow ));
 AND2_X1 \V2/V4/V1/V1/HA1/_0_  (.A1(\V2/V4/V1/V1/w2 ),
    .A2(\V2/V4/V1/V1/w1 ),
    .ZN(\V2/V4/V1/V1/w4 ));
 XOR2_X2 \V2/V4/V1/V1/HA1/_1_  (.A(\V2/V4/V1/V1/w2 ),
    .B(\V2/V4/V1/V1/w1 ),
    .Z(\V2/v4 [1]));
 AND2_X1 \V2/V4/V1/V1/HA2/_0_  (.A1(\V2/V4/V1/V1/w4 ),
    .A2(\V2/V4/V1/V1/w3 ),
    .ZN(\V2/V4/V1/v1 [3]));
 XOR2_X2 \V2/V4/V1/V1/HA2/_1_  (.A(\V2/V4/V1/V1/w4 ),
    .B(\V2/V4/V1/V1/w3 ),
    .Z(\V2/V4/V1/v1 [2]));
 AND2_X1 \V2/V4/V1/V1/_0_  (.A1(net33),
    .A2(net12),
    .ZN(\V2/v4 [0]));
 AND2_X1 \V2/V4/V1/V1/_1_  (.A1(net33),
    .A2(net11),
    .ZN(\V2/V4/V1/V1/w1 ));
 AND2_X1 \V2/V4/V1/V1/_2_  (.A1(net12),
    .A2(net32),
    .ZN(\V2/V4/V1/V1/w2 ));
 AND2_X1 \V2/V4/V1/V1/_3_  (.A1(net11),
    .A2(net32),
    .ZN(\V2/V4/V1/V1/w3 ));
 AND2_X1 \V2/V4/V1/V2/HA1/_0_  (.A1(\V2/V4/V1/V2/w2 ),
    .A2(\V2/V4/V1/V2/w1 ),
    .ZN(\V2/V4/V1/V2/w4 ));
 XOR2_X2 \V2/V4/V1/V2/HA1/_1_  (.A(\V2/V4/V1/V2/w2 ),
    .B(\V2/V4/V1/V2/w1 ),
    .Z(\V2/V4/V1/v2 [1]));
 AND2_X1 \V2/V4/V1/V2/HA2/_0_  (.A1(\V2/V4/V1/V2/w4 ),
    .A2(\V2/V4/V1/V2/w3 ),
    .ZN(\V2/V4/V1/v2 [3]));
 XOR2_X2 \V2/V4/V1/V2/HA2/_1_  (.A(\V2/V4/V1/V2/w4 ),
    .B(\V2/V4/V1/V2/w3 ),
    .Z(\V2/V4/V1/v2 [2]));
 AND2_X1 \V2/V4/V1/V2/_0_  (.A1(net31),
    .A2(net12),
    .ZN(\V2/V4/V1/v2 [0]));
 AND2_X1 \V2/V4/V1/V2/_1_  (.A1(net31),
    .A2(net11),
    .ZN(\V2/V4/V1/V2/w1 ));
 AND2_X1 \V2/V4/V1/V2/_2_  (.A1(net12),
    .A2(net30),
    .ZN(\V2/V4/V1/V2/w2 ));
 AND2_X1 \V2/V4/V1/V2/_3_  (.A1(net11),
    .A2(net30),
    .ZN(\V2/V4/V1/V2/w3 ));
 AND2_X1 \V2/V4/V1/V3/HA1/_0_  (.A1(\V2/V4/V1/V3/w2 ),
    .A2(\V2/V4/V1/V3/w1 ),
    .ZN(\V2/V4/V1/V3/w4 ));
 XOR2_X2 \V2/V4/V1/V3/HA1/_1_  (.A(\V2/V4/V1/V3/w2 ),
    .B(\V2/V4/V1/V3/w1 ),
    .Z(\V2/V4/V1/v3 [1]));
 AND2_X1 \V2/V4/V1/V3/HA2/_0_  (.A1(\V2/V4/V1/V3/w4 ),
    .A2(\V2/V4/V1/V3/w3 ),
    .ZN(\V2/V4/V1/v3 [3]));
 XOR2_X2 \V2/V4/V1/V3/HA2/_1_  (.A(\V2/V4/V1/V3/w4 ),
    .B(\V2/V4/V1/V3/w3 ),
    .Z(\V2/V4/V1/v3 [2]));
 AND2_X1 \V2/V4/V1/V3/_0_  (.A1(net33),
    .A2(B[10]),
    .ZN(\V2/V4/V1/v3 [0]));
 AND2_X1 \V2/V4/V1/V3/_1_  (.A1(net33),
    .A2(B[11]),
    .ZN(\V2/V4/V1/V3/w1 ));
 AND2_X1 \V2/V4/V1/V3/_2_  (.A1(B[10]),
    .A2(net32),
    .ZN(\V2/V4/V1/V3/w2 ));
 AND2_X1 \V2/V4/V1/V3/_3_  (.A1(B[11]),
    .A2(net32),
    .ZN(\V2/V4/V1/V3/w3 ));
 AND2_X1 \V2/V4/V1/V4/HA1/_0_  (.A1(\V2/V4/V1/V4/w2 ),
    .A2(\V2/V4/V1/V4/w1 ),
    .ZN(\V2/V4/V1/V4/w4 ));
 XOR2_X2 \V2/V4/V1/V4/HA1/_1_  (.A(\V2/V4/V1/V4/w2 ),
    .B(\V2/V4/V1/V4/w1 ),
    .Z(\V2/V4/V1/v4 [1]));
 AND2_X1 \V2/V4/V1/V4/HA2/_0_  (.A1(\V2/V4/V1/V4/w4 ),
    .A2(\V2/V4/V1/V4/w3 ),
    .ZN(\V2/V4/V1/v4 [3]));
 XOR2_X2 \V2/V4/V1/V4/HA2/_1_  (.A(\V2/V4/V1/V4/w4 ),
    .B(\V2/V4/V1/V4/w3 ),
    .Z(\V2/V4/V1/v4 [2]));
 AND2_X1 \V2/V4/V1/V4/_0_  (.A1(net31),
    .A2(B[10]),
    .ZN(\V2/V4/V1/v4 [0]));
 AND2_X1 \V2/V4/V1/V4/_1_  (.A1(net31),
    .A2(B[11]),
    .ZN(\V2/V4/V1/V4/w1 ));
 AND2_X1 \V2/V4/V1/V4/_2_  (.A1(B[10]),
    .A2(net30),
    .ZN(\V2/V4/V1/V4/w2 ));
 AND2_X1 \V2/V4/V1/V4/_3_  (.A1(B[11]),
    .A2(net30),
    .ZN(\V2/V4/V1/V4/w3 ));
 OR2_X1 \V2/V4/V1/_0_  (.A1(\V2/V4/V1/c1 ),
    .A2(\V2/V4/V1/c2 ),
    .ZN(\V2/V4/V1/c3 ));
 AND2_X1 \V2/V4/V2/A1/M1/M1/_0_  (.A1(\V2/V4/V2/v2 [0]),
    .A2(\V2/V4/V2/v3 [0]),
    .ZN(\V2/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M1/M1/_1_  (.A(\V2/V4/V2/v2 [0]),
    .B(\V2/V4/V2/v3 [0]),
    .Z(\V2/V4/V2/A1/M1/s1 ));
 AND2_X1 \V2/V4/V2/A1/M1/M2/_0_  (.A1(\V2/V4/V2/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M1/M2/_1_  (.A(\V2/V4/V2/A1/M1/s1 ),
    .B(net9),
    .Z(\V2/V4/V2/s1 [0]));
 OR2_X1 \V2/V4/V2/A1/M1/_0_  (.A1(\V2/V4/V2/A1/M1/c1 ),
    .A2(\V2/V4/V2/A1/M1/c2 ),
    .ZN(\V2/V4/V2/A1/c1 ));
 AND2_X1 \V2/V4/V2/A1/M2/M1/_0_  (.A1(\V2/V4/V2/v2 [1]),
    .A2(\V2/V4/V2/v3 [1]),
    .ZN(\V2/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M2/M1/_1_  (.A(\V2/V4/V2/v2 [1]),
    .B(\V2/V4/V2/v3 [1]),
    .Z(\V2/V4/V2/A1/M2/s1 ));
 AND2_X1 \V2/V4/V2/A1/M2/M2/_0_  (.A1(\V2/V4/V2/A1/M2/s1 ),
    .A2(\V2/V4/V2/A1/c1 ),
    .ZN(\V2/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M2/M2/_1_  (.A(\V2/V4/V2/A1/M2/s1 ),
    .B(\V2/V4/V2/A1/c1 ),
    .Z(\V2/V4/V2/s1 [1]));
 OR2_X1 \V2/V4/V2/A1/M2/_0_  (.A1(\V2/V4/V2/A1/M2/c1 ),
    .A2(\V2/V4/V2/A1/M2/c2 ),
    .ZN(\V2/V4/V2/A1/c2 ));
 AND2_X1 \V2/V4/V2/A1/M3/M1/_0_  (.A1(\V2/V4/V2/v2 [2]),
    .A2(\V2/V4/V2/v3 [2]),
    .ZN(\V2/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M3/M1/_1_  (.A(\V2/V4/V2/v2 [2]),
    .B(\V2/V4/V2/v3 [2]),
    .Z(\V2/V4/V2/A1/M3/s1 ));
 AND2_X1 \V2/V4/V2/A1/M3/M2/_0_  (.A1(\V2/V4/V2/A1/M3/s1 ),
    .A2(\V2/V4/V2/A1/c2 ),
    .ZN(\V2/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M3/M2/_1_  (.A(\V2/V4/V2/A1/M3/s1 ),
    .B(\V2/V4/V2/A1/c2 ),
    .Z(\V2/V4/V2/s1 [2]));
 OR2_X1 \V2/V4/V2/A1/M3/_0_  (.A1(\V2/V4/V2/A1/M3/c1 ),
    .A2(\V2/V4/V2/A1/M3/c2 ),
    .ZN(\V2/V4/V2/A1/c3 ));
 AND2_X1 \V2/V4/V2/A1/M4/M1/_0_  (.A1(\V2/V4/V2/v2 [3]),
    .A2(\V2/V4/V2/v3 [3]),
    .ZN(\V2/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A1/M4/M1/_1_  (.A(\V2/V4/V2/v2 [3]),
    .B(\V2/V4/V2/v3 [3]),
    .Z(\V2/V4/V2/A1/M4/s1 ));
 AND2_X1 \V2/V4/V2/A1/M4/M2/_0_  (.A1(\V2/V4/V2/A1/M4/s1 ),
    .A2(\V2/V4/V2/A1/c3 ),
    .ZN(\V2/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A1/M4/M2/_1_  (.A(\V2/V4/V2/A1/M4/s1 ),
    .B(\V2/V4/V2/A1/c3 ),
    .Z(\V2/V4/V2/s1 [3]));
 OR2_X1 \V2/V4/V2/A1/M4/_0_  (.A1(\V2/V4/V2/A1/M4/c1 ),
    .A2(\V2/V4/V2/A1/M4/c2 ),
    .ZN(\V2/V4/V2/c1 ));
 AND2_X1 \V2/V4/V2/A2/M1/M1/_0_  (.A1(\V2/V4/V2/s1 [0]),
    .A2(\V2/V4/V2/v1 [2]),
    .ZN(\V2/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M1/M1/_1_  (.A(\V2/V4/V2/s1 [0]),
    .B(\V2/V4/V2/v1 [2]),
    .Z(\V2/V4/V2/A2/M1/s1 ));
 AND2_X1 \V2/V4/V2/A2/M1/M2/_0_  (.A1(\V2/V4/V2/A2/M1/s1 ),
    .A2(net9),
    .ZN(\V2/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M1/M2/_1_  (.A(\V2/V4/V2/A2/M1/s1 ),
    .B(net9),
    .Z(\V2/V4/v2 [2]));
 OR2_X1 \V2/V4/V2/A2/M1/_0_  (.A1(\V2/V4/V2/A2/M1/c1 ),
    .A2(\V2/V4/V2/A2/M1/c2 ),
    .ZN(\V2/V4/V2/A2/c1 ));
 AND2_X1 \V2/V4/V2/A2/M2/M1/_0_  (.A1(\V2/V4/V2/s1 [1]),
    .A2(\V2/V4/V2/v1 [3]),
    .ZN(\V2/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M2/M1/_1_  (.A(\V2/V4/V2/s1 [1]),
    .B(\V2/V4/V2/v1 [3]),
    .Z(\V2/V4/V2/A2/M2/s1 ));
 AND2_X1 \V2/V4/V2/A2/M2/M2/_0_  (.A1(\V2/V4/V2/A2/M2/s1 ),
    .A2(\V2/V4/V2/A2/c1 ),
    .ZN(\V2/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M2/M2/_1_  (.A(\V2/V4/V2/A2/M2/s1 ),
    .B(\V2/V4/V2/A2/c1 ),
    .Z(\V2/V4/v2 [3]));
 OR2_X1 \V2/V4/V2/A2/M2/_0_  (.A1(\V2/V4/V2/A2/M2/c1 ),
    .A2(\V2/V4/V2/A2/M2/c2 ),
    .ZN(\V2/V4/V2/A2/c2 ));
 AND2_X1 \V2/V4/V2/A2/M3/M1/_0_  (.A1(\V2/V4/V2/s1 [2]),
    .A2(net9),
    .ZN(\V2/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M3/M1/_1_  (.A(\V2/V4/V2/s1 [2]),
    .B(net9),
    .Z(\V2/V4/V2/A2/M3/s1 ));
 AND2_X1 \V2/V4/V2/A2/M3/M2/_0_  (.A1(\V2/V4/V2/A2/M3/s1 ),
    .A2(\V2/V4/V2/A2/c2 ),
    .ZN(\V2/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M3/M2/_1_  (.A(\V2/V4/V2/A2/M3/s1 ),
    .B(\V2/V4/V2/A2/c2 ),
    .Z(\V2/V4/V2/s2 [2]));
 OR2_X1 \V2/V4/V2/A2/M3/_0_  (.A1(\V2/V4/V2/A2/M3/c1 ),
    .A2(\V2/V4/V2/A2/M3/c2 ),
    .ZN(\V2/V4/V2/A2/c3 ));
 AND2_X1 \V2/V4/V2/A2/M4/M1/_0_  (.A1(\V2/V4/V2/s1 [3]),
    .A2(net9),
    .ZN(\V2/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A2/M4/M1/_1_  (.A(\V2/V4/V2/s1 [3]),
    .B(net9),
    .Z(\V2/V4/V2/A2/M4/s1 ));
 AND2_X1 \V2/V4/V2/A2/M4/M2/_0_  (.A1(\V2/V4/V2/A2/M4/s1 ),
    .A2(\V2/V4/V2/A2/c3 ),
    .ZN(\V2/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A2/M4/M2/_1_  (.A(\V2/V4/V2/A2/M4/s1 ),
    .B(\V2/V4/V2/A2/c3 ),
    .Z(\V2/V4/V2/s2 [3]));
 OR2_X1 \V2/V4/V2/A2/M4/_0_  (.A1(\V2/V4/V2/A2/M4/c1 ),
    .A2(\V2/V4/V2/A2/M4/c2 ),
    .ZN(\V2/V4/V2/c2 ));
 AND2_X1 \V2/V4/V2/A3/M1/M1/_0_  (.A1(\V2/V4/V2/v4 [0]),
    .A2(\V2/V4/V2/s2 [2]),
    .ZN(\V2/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M1/M1/_1_  (.A(\V2/V4/V2/v4 [0]),
    .B(\V2/V4/V2/s2 [2]),
    .Z(\V2/V4/V2/A3/M1/s1 ));
 AND2_X1 \V2/V4/V2/A3/M1/M2/_0_  (.A1(\V2/V4/V2/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M1/M2/_1_  (.A(\V2/V4/V2/A3/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/v2 [4]));
 OR2_X1 \V2/V4/V2/A3/M1/_0_  (.A1(\V2/V4/V2/A3/M1/c1 ),
    .A2(\V2/V4/V2/A3/M1/c2 ),
    .ZN(\V2/V4/V2/A3/c1 ));
 AND2_X1 \V2/V4/V2/A3/M2/M1/_0_  (.A1(\V2/V4/V2/v4 [1]),
    .A2(\V2/V4/V2/s2 [3]),
    .ZN(\V2/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M2/M1/_1_  (.A(\V2/V4/V2/v4 [1]),
    .B(\V2/V4/V2/s2 [3]),
    .Z(\V2/V4/V2/A3/M2/s1 ));
 AND2_X1 \V2/V4/V2/A3/M2/M2/_0_  (.A1(\V2/V4/V2/A3/M2/s1 ),
    .A2(\V2/V4/V2/A3/c1 ),
    .ZN(\V2/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M2/M2/_1_  (.A(\V2/V4/V2/A3/M2/s1 ),
    .B(\V2/V4/V2/A3/c1 ),
    .Z(\V2/V4/v2 [5]));
 OR2_X1 \V2/V4/V2/A3/M2/_0_  (.A1(\V2/V4/V2/A3/M2/c1 ),
    .A2(\V2/V4/V2/A3/M2/c2 ),
    .ZN(\V2/V4/V2/A3/c2 ));
 AND2_X1 \V2/V4/V2/A3/M3/M1/_0_  (.A1(\V2/V4/V2/v4 [2]),
    .A2(\V2/V4/V2/c3 ),
    .ZN(\V2/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M3/M1/_1_  (.A(\V2/V4/V2/v4 [2]),
    .B(\V2/V4/V2/c3 ),
    .Z(\V2/V4/V2/A3/M3/s1 ));
 AND2_X1 \V2/V4/V2/A3/M3/M2/_0_  (.A1(\V2/V4/V2/A3/M3/s1 ),
    .A2(\V2/V4/V2/A3/c2 ),
    .ZN(\V2/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M3/M2/_1_  (.A(\V2/V4/V2/A3/M3/s1 ),
    .B(\V2/V4/V2/A3/c2 ),
    .Z(\V2/V4/v2 [6]));
 OR2_X1 \V2/V4/V2/A3/M3/_0_  (.A1(\V2/V4/V2/A3/M3/c1 ),
    .A2(\V2/V4/V2/A3/M3/c2 ),
    .ZN(\V2/V4/V2/A3/c3 ));
 AND2_X1 \V2/V4/V2/A3/M4/M1/_0_  (.A1(\V2/V4/V2/v4 [3]),
    .A2(net9),
    .ZN(\V2/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V2/A3/M4/M1/_1_  (.A(\V2/V4/V2/v4 [3]),
    .B(net9),
    .Z(\V2/V4/V2/A3/M4/s1 ));
 AND2_X1 \V2/V4/V2/A3/M4/M2/_0_  (.A1(\V2/V4/V2/A3/M4/s1 ),
    .A2(\V2/V4/V2/A3/c3 ),
    .ZN(\V2/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V2/A3/M4/M2/_1_  (.A(\V2/V4/V2/A3/M4/s1 ),
    .B(\V2/V4/V2/A3/c3 ),
    .Z(\V2/V4/v2 [7]));
 OR2_X1 \V2/V4/V2/A3/M4/_0_  (.A1(\V2/V4/V2/A3/M4/c1 ),
    .A2(\V2/V4/V2/A3/M4/c2 ),
    .ZN(\V2/V4/V2/overflow ));
 AND2_X1 \V2/V4/V2/V1/HA1/_0_  (.A1(\V2/V4/V2/V1/w2 ),
    .A2(\V2/V4/V2/V1/w1 ),
    .ZN(\V2/V4/V2/V1/w4 ));
 XOR2_X2 \V2/V4/V2/V1/HA1/_1_  (.A(\V2/V4/V2/V1/w2 ),
    .B(\V2/V4/V2/V1/w1 ),
    .Z(\V2/V4/v2 [1]));
 AND2_X1 \V2/V4/V2/V1/HA2/_0_  (.A1(\V2/V4/V2/V1/w4 ),
    .A2(\V2/V4/V2/V1/w3 ),
    .ZN(\V2/V4/V2/v1 [3]));
 XOR2_X2 \V2/V4/V2/V1/HA2/_1_  (.A(\V2/V4/V2/V1/w4 ),
    .B(\V2/V4/V2/V1/w3 ),
    .Z(\V2/V4/V2/v1 [2]));
 AND2_X1 \V2/V4/V2/V1/_0_  (.A1(net29),
    .A2(net12),
    .ZN(\V2/V4/v2 [0]));
 AND2_X1 \V2/V4/V2/V1/_1_  (.A1(net29),
    .A2(net11),
    .ZN(\V2/V4/V2/V1/w1 ));
 AND2_X1 \V2/V4/V2/V1/_2_  (.A1(net12),
    .A2(net28),
    .ZN(\V2/V4/V2/V1/w2 ));
 AND2_X1 \V2/V4/V2/V1/_3_  (.A1(net11),
    .A2(net28),
    .ZN(\V2/V4/V2/V1/w3 ));
 AND2_X1 \V2/V4/V2/V2/HA1/_0_  (.A1(\V2/V4/V2/V2/w2 ),
    .A2(\V2/V4/V2/V2/w1 ),
    .ZN(\V2/V4/V2/V2/w4 ));
 XOR2_X2 \V2/V4/V2/V2/HA1/_1_  (.A(\V2/V4/V2/V2/w2 ),
    .B(\V2/V4/V2/V2/w1 ),
    .Z(\V2/V4/V2/v2 [1]));
 AND2_X1 \V2/V4/V2/V2/HA2/_0_  (.A1(\V2/V4/V2/V2/w4 ),
    .A2(\V2/V4/V2/V2/w3 ),
    .ZN(\V2/V4/V2/v2 [3]));
 XOR2_X2 \V2/V4/V2/V2/HA2/_1_  (.A(\V2/V4/V2/V2/w4 ),
    .B(\V2/V4/V2/V2/w3 ),
    .Z(\V2/V4/V2/v2 [2]));
 AND2_X1 \V2/V4/V2/V2/_0_  (.A1(net27),
    .A2(net12),
    .ZN(\V2/V4/V2/v2 [0]));
 AND2_X1 \V2/V4/V2/V2/_1_  (.A1(net27),
    .A2(net11),
    .ZN(\V2/V4/V2/V2/w1 ));
 AND2_X1 \V2/V4/V2/V2/_2_  (.A1(net12),
    .A2(net26),
    .ZN(\V2/V4/V2/V2/w2 ));
 AND2_X1 \V2/V4/V2/V2/_3_  (.A1(net11),
    .A2(net26),
    .ZN(\V2/V4/V2/V2/w3 ));
 AND2_X1 \V2/V4/V2/V3/HA1/_0_  (.A1(\V2/V4/V2/V3/w2 ),
    .A2(\V2/V4/V2/V3/w1 ),
    .ZN(\V2/V4/V2/V3/w4 ));
 XOR2_X2 \V2/V4/V2/V3/HA1/_1_  (.A(\V2/V4/V2/V3/w2 ),
    .B(\V2/V4/V2/V3/w1 ),
    .Z(\V2/V4/V2/v3 [1]));
 AND2_X1 \V2/V4/V2/V3/HA2/_0_  (.A1(\V2/V4/V2/V3/w4 ),
    .A2(\V2/V4/V2/V3/w3 ),
    .ZN(\V2/V4/V2/v3 [3]));
 XOR2_X2 \V2/V4/V2/V3/HA2/_1_  (.A(\V2/V4/V2/V3/w4 ),
    .B(\V2/V4/V2/V3/w3 ),
    .Z(\V2/V4/V2/v3 [2]));
 AND2_X1 \V2/V4/V2/V3/_0_  (.A1(net29),
    .A2(B[10]),
    .ZN(\V2/V4/V2/v3 [0]));
 AND2_X1 \V2/V4/V2/V3/_1_  (.A1(net29),
    .A2(B[11]),
    .ZN(\V2/V4/V2/V3/w1 ));
 AND2_X1 \V2/V4/V2/V3/_2_  (.A1(B[10]),
    .A2(net28),
    .ZN(\V2/V4/V2/V3/w2 ));
 AND2_X1 \V2/V4/V2/V3/_3_  (.A1(B[11]),
    .A2(net28),
    .ZN(\V2/V4/V2/V3/w3 ));
 AND2_X1 \V2/V4/V2/V4/HA1/_0_  (.A1(\V2/V4/V2/V4/w2 ),
    .A2(\V2/V4/V2/V4/w1 ),
    .ZN(\V2/V4/V2/V4/w4 ));
 XOR2_X2 \V2/V4/V2/V4/HA1/_1_  (.A(\V2/V4/V2/V4/w2 ),
    .B(\V2/V4/V2/V4/w1 ),
    .Z(\V2/V4/V2/v4 [1]));
 AND2_X1 \V2/V4/V2/V4/HA2/_0_  (.A1(\V2/V4/V2/V4/w4 ),
    .A2(\V2/V4/V2/V4/w3 ),
    .ZN(\V2/V4/V2/v4 [3]));
 XOR2_X2 \V2/V4/V2/V4/HA2/_1_  (.A(\V2/V4/V2/V4/w4 ),
    .B(\V2/V4/V2/V4/w3 ),
    .Z(\V2/V4/V2/v4 [2]));
 AND2_X1 \V2/V4/V2/V4/_0_  (.A1(net27),
    .A2(B[10]),
    .ZN(\V2/V4/V2/v4 [0]));
 AND2_X1 \V2/V4/V2/V4/_1_  (.A1(net27),
    .A2(B[11]),
    .ZN(\V2/V4/V2/V4/w1 ));
 AND2_X1 \V2/V4/V2/V4/_2_  (.A1(B[10]),
    .A2(net26),
    .ZN(\V2/V4/V2/V4/w2 ));
 AND2_X1 \V2/V4/V2/V4/_3_  (.A1(B[11]),
    .A2(net26),
    .ZN(\V2/V4/V2/V4/w3 ));
 OR2_X1 \V2/V4/V2/_0_  (.A1(\V2/V4/V2/c1 ),
    .A2(\V2/V4/V2/c2 ),
    .ZN(\V2/V4/V2/c3 ));
 AND2_X1 \V2/V4/V3/A1/M1/M1/_0_  (.A1(\V2/V4/V3/v2 [0]),
    .A2(\V2/V4/V3/v3 [0]),
    .ZN(\V2/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M1/M1/_1_  (.A(\V2/V4/V3/v2 [0]),
    .B(\V2/V4/V3/v3 [0]),
    .Z(\V2/V4/V3/A1/M1/s1 ));
 AND2_X1 \V2/V4/V3/A1/M1/M2/_0_  (.A1(\V2/V4/V3/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M1/M2/_1_  (.A(\V2/V4/V3/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/V3/s1 [0]));
 OR2_X1 \V2/V4/V3/A1/M1/_0_  (.A1(\V2/V4/V3/A1/M1/c1 ),
    .A2(\V2/V4/V3/A1/M1/c2 ),
    .ZN(\V2/V4/V3/A1/c1 ));
 AND2_X1 \V2/V4/V3/A1/M2/M1/_0_  (.A1(\V2/V4/V3/v2 [1]),
    .A2(\V2/V4/V3/v3 [1]),
    .ZN(\V2/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M2/M1/_1_  (.A(\V2/V4/V3/v2 [1]),
    .B(\V2/V4/V3/v3 [1]),
    .Z(\V2/V4/V3/A1/M2/s1 ));
 AND2_X1 \V2/V4/V3/A1/M2/M2/_0_  (.A1(\V2/V4/V3/A1/M2/s1 ),
    .A2(\V2/V4/V3/A1/c1 ),
    .ZN(\V2/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M2/M2/_1_  (.A(\V2/V4/V3/A1/M2/s1 ),
    .B(\V2/V4/V3/A1/c1 ),
    .Z(\V2/V4/V3/s1 [1]));
 OR2_X1 \V2/V4/V3/A1/M2/_0_  (.A1(\V2/V4/V3/A1/M2/c1 ),
    .A2(\V2/V4/V3/A1/M2/c2 ),
    .ZN(\V2/V4/V3/A1/c2 ));
 AND2_X1 \V2/V4/V3/A1/M3/M1/_0_  (.A1(\V2/V4/V3/v2 [2]),
    .A2(\V2/V4/V3/v3 [2]),
    .ZN(\V2/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M3/M1/_1_  (.A(\V2/V4/V3/v2 [2]),
    .B(\V2/V4/V3/v3 [2]),
    .Z(\V2/V4/V3/A1/M3/s1 ));
 AND2_X1 \V2/V4/V3/A1/M3/M2/_0_  (.A1(\V2/V4/V3/A1/M3/s1 ),
    .A2(\V2/V4/V3/A1/c2 ),
    .ZN(\V2/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M3/M2/_1_  (.A(\V2/V4/V3/A1/M3/s1 ),
    .B(\V2/V4/V3/A1/c2 ),
    .Z(\V2/V4/V3/s1 [2]));
 OR2_X1 \V2/V4/V3/A1/M3/_0_  (.A1(\V2/V4/V3/A1/M3/c1 ),
    .A2(\V2/V4/V3/A1/M3/c2 ),
    .ZN(\V2/V4/V3/A1/c3 ));
 AND2_X1 \V2/V4/V3/A1/M4/M1/_0_  (.A1(\V2/V4/V3/v2 [3]),
    .A2(\V2/V4/V3/v3 [3]),
    .ZN(\V2/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A1/M4/M1/_1_  (.A(\V2/V4/V3/v2 [3]),
    .B(\V2/V4/V3/v3 [3]),
    .Z(\V2/V4/V3/A1/M4/s1 ));
 AND2_X1 \V2/V4/V3/A1/M4/M2/_0_  (.A1(\V2/V4/V3/A1/M4/s1 ),
    .A2(\V2/V4/V3/A1/c3 ),
    .ZN(\V2/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A1/M4/M2/_1_  (.A(\V2/V4/V3/A1/M4/s1 ),
    .B(\V2/V4/V3/A1/c3 ),
    .Z(\V2/V4/V3/s1 [3]));
 OR2_X1 \V2/V4/V3/A1/M4/_0_  (.A1(\V2/V4/V3/A1/M4/c1 ),
    .A2(\V2/V4/V3/A1/M4/c2 ),
    .ZN(\V2/V4/V3/c1 ));
 AND2_X1 \V2/V4/V3/A2/M1/M1/_0_  (.A1(\V2/V4/V3/s1 [0]),
    .A2(\V2/V4/V3/v1 [2]),
    .ZN(\V2/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M1/M1/_1_  (.A(\V2/V4/V3/s1 [0]),
    .B(\V2/V4/V3/v1 [2]),
    .Z(\V2/V4/V3/A2/M1/s1 ));
 AND2_X1 \V2/V4/V3/A2/M1/M2/_0_  (.A1(\V2/V4/V3/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M1/M2/_1_  (.A(\V2/V4/V3/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/v3 [2]));
 OR2_X1 \V2/V4/V3/A2/M1/_0_  (.A1(\V2/V4/V3/A2/M1/c1 ),
    .A2(\V2/V4/V3/A2/M1/c2 ),
    .ZN(\V2/V4/V3/A2/c1 ));
 AND2_X1 \V2/V4/V3/A2/M2/M1/_0_  (.A1(\V2/V4/V3/s1 [1]),
    .A2(\V2/V4/V3/v1 [3]),
    .ZN(\V2/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M2/M1/_1_  (.A(\V2/V4/V3/s1 [1]),
    .B(\V2/V4/V3/v1 [3]),
    .Z(\V2/V4/V3/A2/M2/s1 ));
 AND2_X1 \V2/V4/V3/A2/M2/M2/_0_  (.A1(\V2/V4/V3/A2/M2/s1 ),
    .A2(\V2/V4/V3/A2/c1 ),
    .ZN(\V2/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M2/M2/_1_  (.A(\V2/V4/V3/A2/M2/s1 ),
    .B(\V2/V4/V3/A2/c1 ),
    .Z(\V2/V4/v3 [3]));
 OR2_X1 \V2/V4/V3/A2/M2/_0_  (.A1(\V2/V4/V3/A2/M2/c1 ),
    .A2(\V2/V4/V3/A2/M2/c2 ),
    .ZN(\V2/V4/V3/A2/c2 ));
 AND2_X1 \V2/V4/V3/A2/M3/M1/_0_  (.A1(\V2/V4/V3/s1 [2]),
    .A2(net7),
    .ZN(\V2/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M3/M1/_1_  (.A(\V2/V4/V3/s1 [2]),
    .B(net7),
    .Z(\V2/V4/V3/A2/M3/s1 ));
 AND2_X1 \V2/V4/V3/A2/M3/M2/_0_  (.A1(\V2/V4/V3/A2/M3/s1 ),
    .A2(\V2/V4/V3/A2/c2 ),
    .ZN(\V2/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M3/M2/_1_  (.A(\V2/V4/V3/A2/M3/s1 ),
    .B(\V2/V4/V3/A2/c2 ),
    .Z(\V2/V4/V3/s2 [2]));
 OR2_X1 \V2/V4/V3/A2/M3/_0_  (.A1(\V2/V4/V3/A2/M3/c1 ),
    .A2(\V2/V4/V3/A2/M3/c2 ),
    .ZN(\V2/V4/V3/A2/c3 ));
 AND2_X1 \V2/V4/V3/A2/M4/M1/_0_  (.A1(\V2/V4/V3/s1 [3]),
    .A2(net7),
    .ZN(\V2/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A2/M4/M1/_1_  (.A(\V2/V4/V3/s1 [3]),
    .B(net7),
    .Z(\V2/V4/V3/A2/M4/s1 ));
 AND2_X1 \V2/V4/V3/A2/M4/M2/_0_  (.A1(\V2/V4/V3/A2/M4/s1 ),
    .A2(\V2/V4/V3/A2/c3 ),
    .ZN(\V2/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A2/M4/M2/_1_  (.A(\V2/V4/V3/A2/M4/s1 ),
    .B(\V2/V4/V3/A2/c3 ),
    .Z(\V2/V4/V3/s2 [3]));
 OR2_X1 \V2/V4/V3/A2/M4/_0_  (.A1(\V2/V4/V3/A2/M4/c1 ),
    .A2(\V2/V4/V3/A2/M4/c2 ),
    .ZN(\V2/V4/V3/c2 ));
 AND2_X1 \V2/V4/V3/A3/M1/M1/_0_  (.A1(\V2/V4/V3/v4 [0]),
    .A2(\V2/V4/V3/s2 [2]),
    .ZN(\V2/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M1/M1/_1_  (.A(\V2/V4/V3/v4 [0]),
    .B(\V2/V4/V3/s2 [2]),
    .Z(\V2/V4/V3/A3/M1/s1 ));
 AND2_X1 \V2/V4/V3/A3/M1/M2/_0_  (.A1(\V2/V4/V3/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M1/M2/_1_  (.A(\V2/V4/V3/A3/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/v3 [4]));
 OR2_X1 \V2/V4/V3/A3/M1/_0_  (.A1(\V2/V4/V3/A3/M1/c1 ),
    .A2(\V2/V4/V3/A3/M1/c2 ),
    .ZN(\V2/V4/V3/A3/c1 ));
 AND2_X1 \V2/V4/V3/A3/M2/M1/_0_  (.A1(\V2/V4/V3/v4 [1]),
    .A2(\V2/V4/V3/s2 [3]),
    .ZN(\V2/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M2/M1/_1_  (.A(\V2/V4/V3/v4 [1]),
    .B(\V2/V4/V3/s2 [3]),
    .Z(\V2/V4/V3/A3/M2/s1 ));
 AND2_X1 \V2/V4/V3/A3/M2/M2/_0_  (.A1(\V2/V4/V3/A3/M2/s1 ),
    .A2(\V2/V4/V3/A3/c1 ),
    .ZN(\V2/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M2/M2/_1_  (.A(\V2/V4/V3/A3/M2/s1 ),
    .B(\V2/V4/V3/A3/c1 ),
    .Z(\V2/V4/v3 [5]));
 OR2_X1 \V2/V4/V3/A3/M2/_0_  (.A1(\V2/V4/V3/A3/M2/c1 ),
    .A2(\V2/V4/V3/A3/M2/c2 ),
    .ZN(\V2/V4/V3/A3/c2 ));
 AND2_X1 \V2/V4/V3/A3/M3/M1/_0_  (.A1(\V2/V4/V3/v4 [2]),
    .A2(\V2/V4/V3/c3 ),
    .ZN(\V2/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M3/M1/_1_  (.A(\V2/V4/V3/v4 [2]),
    .B(\V2/V4/V3/c3 ),
    .Z(\V2/V4/V3/A3/M3/s1 ));
 AND2_X1 \V2/V4/V3/A3/M3/M2/_0_  (.A1(\V2/V4/V3/A3/M3/s1 ),
    .A2(\V2/V4/V3/A3/c2 ),
    .ZN(\V2/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M3/M2/_1_  (.A(\V2/V4/V3/A3/M3/s1 ),
    .B(\V2/V4/V3/A3/c2 ),
    .Z(\V2/V4/v3 [6]));
 OR2_X1 \V2/V4/V3/A3/M3/_0_  (.A1(\V2/V4/V3/A3/M3/c1 ),
    .A2(\V2/V4/V3/A3/M3/c2 ),
    .ZN(\V2/V4/V3/A3/c3 ));
 AND2_X1 \V2/V4/V3/A3/M4/M1/_0_  (.A1(\V2/V4/V3/v4 [3]),
    .A2(net7),
    .ZN(\V2/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V3/A3/M4/M1/_1_  (.A(\V2/V4/V3/v4 [3]),
    .B(net7),
    .Z(\V2/V4/V3/A3/M4/s1 ));
 AND2_X1 \V2/V4/V3/A3/M4/M2/_0_  (.A1(\V2/V4/V3/A3/M4/s1 ),
    .A2(\V2/V4/V3/A3/c3 ),
    .ZN(\V2/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V3/A3/M4/M2/_1_  (.A(\V2/V4/V3/A3/M4/s1 ),
    .B(\V2/V4/V3/A3/c3 ),
    .Z(\V2/V4/v3 [7]));
 OR2_X1 \V2/V4/V3/A3/M4/_0_  (.A1(\V2/V4/V3/A3/M4/c1 ),
    .A2(\V2/V4/V3/A3/M4/c2 ),
    .ZN(\V2/V4/V3/overflow ));
 AND2_X1 \V2/V4/V3/V1/HA1/_0_  (.A1(\V2/V4/V3/V1/w2 ),
    .A2(\V2/V4/V3/V1/w1 ),
    .ZN(\V2/V4/V3/V1/w4 ));
 XOR2_X2 \V2/V4/V3/V1/HA1/_1_  (.A(\V2/V4/V3/V1/w2 ),
    .B(\V2/V4/V3/V1/w1 ),
    .Z(\V2/V4/v3 [1]));
 AND2_X1 \V2/V4/V3/V1/HA2/_0_  (.A1(\V2/V4/V3/V1/w4 ),
    .A2(\V2/V4/V3/V1/w3 ),
    .ZN(\V2/V4/V3/v1 [3]));
 XOR2_X2 \V2/V4/V3/V1/HA2/_1_  (.A(\V2/V4/V3/V1/w4 ),
    .B(\V2/V4/V3/V1/w3 ),
    .Z(\V2/V4/V3/v1 [2]));
 AND2_X1 \V2/V4/V3/V1/_0_  (.A1(net33),
    .A2(B[12]),
    .ZN(\V2/V4/v3 [0]));
 AND2_X1 \V2/V4/V3/V1/_1_  (.A1(net33),
    .A2(B[13]),
    .ZN(\V2/V4/V3/V1/w1 ));
 AND2_X1 \V2/V4/V3/V1/_2_  (.A1(B[12]),
    .A2(net32),
    .ZN(\V2/V4/V3/V1/w2 ));
 AND2_X1 \V2/V4/V3/V1/_3_  (.A1(B[13]),
    .A2(net32),
    .ZN(\V2/V4/V3/V1/w3 ));
 AND2_X1 \V2/V4/V3/V2/HA1/_0_  (.A1(\V2/V4/V3/V2/w2 ),
    .A2(\V2/V4/V3/V2/w1 ),
    .ZN(\V2/V4/V3/V2/w4 ));
 XOR2_X2 \V2/V4/V3/V2/HA1/_1_  (.A(\V2/V4/V3/V2/w2 ),
    .B(\V2/V4/V3/V2/w1 ),
    .Z(\V2/V4/V3/v2 [1]));
 AND2_X1 \V2/V4/V3/V2/HA2/_0_  (.A1(\V2/V4/V3/V2/w4 ),
    .A2(\V2/V4/V3/V2/w3 ),
    .ZN(\V2/V4/V3/v2 [3]));
 XOR2_X2 \V2/V4/V3/V2/HA2/_1_  (.A(\V2/V4/V3/V2/w4 ),
    .B(\V2/V4/V3/V2/w3 ),
    .Z(\V2/V4/V3/v2 [2]));
 AND2_X1 \V2/V4/V3/V2/_0_  (.A1(net31),
    .A2(B[12]),
    .ZN(\V2/V4/V3/v2 [0]));
 AND2_X1 \V2/V4/V3/V2/_1_  (.A1(net31),
    .A2(B[13]),
    .ZN(\V2/V4/V3/V2/w1 ));
 AND2_X1 \V2/V4/V3/V2/_2_  (.A1(B[12]),
    .A2(net30),
    .ZN(\V2/V4/V3/V2/w2 ));
 AND2_X1 \V2/V4/V3/V2/_3_  (.A1(B[13]),
    .A2(net30),
    .ZN(\V2/V4/V3/V2/w3 ));
 AND2_X1 \V2/V4/V3/V3/HA1/_0_  (.A1(\V2/V4/V3/V3/w2 ),
    .A2(\V2/V4/V3/V3/w1 ),
    .ZN(\V2/V4/V3/V3/w4 ));
 XOR2_X2 \V2/V4/V3/V3/HA1/_1_  (.A(\V2/V4/V3/V3/w2 ),
    .B(\V2/V4/V3/V3/w1 ),
    .Z(\V2/V4/V3/v3 [1]));
 AND2_X1 \V2/V4/V3/V3/HA2/_0_  (.A1(\V2/V4/V3/V3/w4 ),
    .A2(\V2/V4/V3/V3/w3 ),
    .ZN(\V2/V4/V3/v3 [3]));
 XOR2_X2 \V2/V4/V3/V3/HA2/_1_  (.A(\V2/V4/V3/V3/w4 ),
    .B(\V2/V4/V3/V3/w3 ),
    .Z(\V2/V4/V3/v3 [2]));
 AND2_X1 \V2/V4/V3/V3/_0_  (.A1(net33),
    .A2(B[14]),
    .ZN(\V2/V4/V3/v3 [0]));
 AND2_X1 \V2/V4/V3/V3/_1_  (.A1(net33),
    .A2(B[15]),
    .ZN(\V2/V4/V3/V3/w1 ));
 AND2_X1 \V2/V4/V3/V3/_2_  (.A1(B[14]),
    .A2(net32),
    .ZN(\V2/V4/V3/V3/w2 ));
 AND2_X1 \V2/V4/V3/V3/_3_  (.A1(B[15]),
    .A2(net32),
    .ZN(\V2/V4/V3/V3/w3 ));
 AND2_X1 \V2/V4/V3/V4/HA1/_0_  (.A1(\V2/V4/V3/V4/w2 ),
    .A2(\V2/V4/V3/V4/w1 ),
    .ZN(\V2/V4/V3/V4/w4 ));
 XOR2_X2 \V2/V4/V3/V4/HA1/_1_  (.A(\V2/V4/V3/V4/w2 ),
    .B(\V2/V4/V3/V4/w1 ),
    .Z(\V2/V4/V3/v4 [1]));
 AND2_X1 \V2/V4/V3/V4/HA2/_0_  (.A1(\V2/V4/V3/V4/w4 ),
    .A2(\V2/V4/V3/V4/w3 ),
    .ZN(\V2/V4/V3/v4 [3]));
 XOR2_X2 \V2/V4/V3/V4/HA2/_1_  (.A(\V2/V4/V3/V4/w4 ),
    .B(\V2/V4/V3/V4/w3 ),
    .Z(\V2/V4/V3/v4 [2]));
 AND2_X1 \V2/V4/V3/V4/_0_  (.A1(net31),
    .A2(B[14]),
    .ZN(\V2/V4/V3/v4 [0]));
 AND2_X1 \V2/V4/V3/V4/_1_  (.A1(net31),
    .A2(B[15]),
    .ZN(\V2/V4/V3/V4/w1 ));
 AND2_X1 \V2/V4/V3/V4/_2_  (.A1(B[14]),
    .A2(net30),
    .ZN(\V2/V4/V3/V4/w2 ));
 AND2_X1 \V2/V4/V3/V4/_3_  (.A1(B[15]),
    .A2(net30),
    .ZN(\V2/V4/V3/V4/w3 ));
 OR2_X1 \V2/V4/V3/_0_  (.A1(\V2/V4/V3/c1 ),
    .A2(\V2/V4/V3/c2 ),
    .ZN(\V2/V4/V3/c3 ));
 AND2_X1 \V2/V4/V4/A1/M1/M1/_0_  (.A1(\V2/V4/V4/v2 [0]),
    .A2(\V2/V4/V4/v3 [0]),
    .ZN(\V2/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M1/M1/_1_  (.A(\V2/V4/V4/v2 [0]),
    .B(\V2/V4/V4/v3 [0]),
    .Z(\V2/V4/V4/A1/M1/s1 ));
 AND2_X1 \V2/V4/V4/A1/M1/M2/_0_  (.A1(\V2/V4/V4/A1/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M1/M2/_1_  (.A(\V2/V4/V4/A1/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/V4/s1 [0]));
 OR2_X1 \V2/V4/V4/A1/M1/_0_  (.A1(\V2/V4/V4/A1/M1/c1 ),
    .A2(\V2/V4/V4/A1/M1/c2 ),
    .ZN(\V2/V4/V4/A1/c1 ));
 AND2_X1 \V2/V4/V4/A1/M2/M1/_0_  (.A1(\V2/V4/V4/v2 [1]),
    .A2(\V2/V4/V4/v3 [1]),
    .ZN(\V2/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M2/M1/_1_  (.A(\V2/V4/V4/v2 [1]),
    .B(\V2/V4/V4/v3 [1]),
    .Z(\V2/V4/V4/A1/M2/s1 ));
 AND2_X1 \V2/V4/V4/A1/M2/M2/_0_  (.A1(\V2/V4/V4/A1/M2/s1 ),
    .A2(\V2/V4/V4/A1/c1 ),
    .ZN(\V2/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M2/M2/_1_  (.A(\V2/V4/V4/A1/M2/s1 ),
    .B(\V2/V4/V4/A1/c1 ),
    .Z(\V2/V4/V4/s1 [1]));
 OR2_X1 \V2/V4/V4/A1/M2/_0_  (.A1(\V2/V4/V4/A1/M2/c1 ),
    .A2(\V2/V4/V4/A1/M2/c2 ),
    .ZN(\V2/V4/V4/A1/c2 ));
 AND2_X1 \V2/V4/V4/A1/M3/M1/_0_  (.A1(\V2/V4/V4/v2 [2]),
    .A2(\V2/V4/V4/v3 [2]),
    .ZN(\V2/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M3/M1/_1_  (.A(\V2/V4/V4/v2 [2]),
    .B(\V2/V4/V4/v3 [2]),
    .Z(\V2/V4/V4/A1/M3/s1 ));
 AND2_X1 \V2/V4/V4/A1/M3/M2/_0_  (.A1(\V2/V4/V4/A1/M3/s1 ),
    .A2(\V2/V4/V4/A1/c2 ),
    .ZN(\V2/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M3/M2/_1_  (.A(\V2/V4/V4/A1/M3/s1 ),
    .B(\V2/V4/V4/A1/c2 ),
    .Z(\V2/V4/V4/s1 [2]));
 OR2_X1 \V2/V4/V4/A1/M3/_0_  (.A1(\V2/V4/V4/A1/M3/c1 ),
    .A2(\V2/V4/V4/A1/M3/c2 ),
    .ZN(\V2/V4/V4/A1/c3 ));
 AND2_X1 \V2/V4/V4/A1/M4/M1/_0_  (.A1(\V2/V4/V4/v2 [3]),
    .A2(\V2/V4/V4/v3 [3]),
    .ZN(\V2/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A1/M4/M1/_1_  (.A(\V2/V4/V4/v2 [3]),
    .B(\V2/V4/V4/v3 [3]),
    .Z(\V2/V4/V4/A1/M4/s1 ));
 AND2_X1 \V2/V4/V4/A1/M4/M2/_0_  (.A1(\V2/V4/V4/A1/M4/s1 ),
    .A2(\V2/V4/V4/A1/c3 ),
    .ZN(\V2/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A1/M4/M2/_1_  (.A(\V2/V4/V4/A1/M4/s1 ),
    .B(\V2/V4/V4/A1/c3 ),
    .Z(\V2/V4/V4/s1 [3]));
 OR2_X1 \V2/V4/V4/A1/M4/_0_  (.A1(\V2/V4/V4/A1/M4/c1 ),
    .A2(\V2/V4/V4/A1/M4/c2 ),
    .ZN(\V2/V4/V4/c1 ));
 AND2_X1 \V2/V4/V4/A2/M1/M1/_0_  (.A1(\V2/V4/V4/s1 [0]),
    .A2(\V2/V4/V4/v1 [2]),
    .ZN(\V2/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M1/M1/_1_  (.A(\V2/V4/V4/s1 [0]),
    .B(\V2/V4/V4/v1 [2]),
    .Z(\V2/V4/V4/A2/M1/s1 ));
 AND2_X1 \V2/V4/V4/A2/M1/M2/_0_  (.A1(\V2/V4/V4/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V2/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M1/M2/_1_  (.A(\V2/V4/V4/A2/M1/s1 ),
    .B(net7),
    .Z(\V2/V4/v4 [2]));
 OR2_X1 \V2/V4/V4/A2/M1/_0_  (.A1(\V2/V4/V4/A2/M1/c1 ),
    .A2(\V2/V4/V4/A2/M1/c2 ),
    .ZN(\V2/V4/V4/A2/c1 ));
 AND2_X1 \V2/V4/V4/A2/M2/M1/_0_  (.A1(\V2/V4/V4/s1 [1]),
    .A2(\V2/V4/V4/v1 [3]),
    .ZN(\V2/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M2/M1/_1_  (.A(\V2/V4/V4/s1 [1]),
    .B(\V2/V4/V4/v1 [3]),
    .Z(\V2/V4/V4/A2/M2/s1 ));
 AND2_X1 \V2/V4/V4/A2/M2/M2/_0_  (.A1(\V2/V4/V4/A2/M2/s1 ),
    .A2(\V2/V4/V4/A2/c1 ),
    .ZN(\V2/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M2/M2/_1_  (.A(\V2/V4/V4/A2/M2/s1 ),
    .B(\V2/V4/V4/A2/c1 ),
    .Z(\V2/V4/v4 [3]));
 OR2_X1 \V2/V4/V4/A2/M2/_0_  (.A1(\V2/V4/V4/A2/M2/c1 ),
    .A2(\V2/V4/V4/A2/M2/c2 ),
    .ZN(\V2/V4/V4/A2/c2 ));
 AND2_X1 \V2/V4/V4/A2/M3/M1/_0_  (.A1(\V2/V4/V4/s1 [2]),
    .A2(net6),
    .ZN(\V2/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M3/M1/_1_  (.A(\V2/V4/V4/s1 [2]),
    .B(net6),
    .Z(\V2/V4/V4/A2/M3/s1 ));
 AND2_X1 \V2/V4/V4/A2/M3/M2/_0_  (.A1(\V2/V4/V4/A2/M3/s1 ),
    .A2(\V2/V4/V4/A2/c2 ),
    .ZN(\V2/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M3/M2/_1_  (.A(\V2/V4/V4/A2/M3/s1 ),
    .B(\V2/V4/V4/A2/c2 ),
    .Z(\V2/V4/V4/s2 [2]));
 OR2_X1 \V2/V4/V4/A2/M3/_0_  (.A1(\V2/V4/V4/A2/M3/c1 ),
    .A2(\V2/V4/V4/A2/M3/c2 ),
    .ZN(\V2/V4/V4/A2/c3 ));
 AND2_X1 \V2/V4/V4/A2/M4/M1/_0_  (.A1(\V2/V4/V4/s1 [3]),
    .A2(net6),
    .ZN(\V2/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A2/M4/M1/_1_  (.A(\V2/V4/V4/s1 [3]),
    .B(net6),
    .Z(\V2/V4/V4/A2/M4/s1 ));
 AND2_X1 \V2/V4/V4/A2/M4/M2/_0_  (.A1(\V2/V4/V4/A2/M4/s1 ),
    .A2(\V2/V4/V4/A2/c3 ),
    .ZN(\V2/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A2/M4/M2/_1_  (.A(\V2/V4/V4/A2/M4/s1 ),
    .B(\V2/V4/V4/A2/c3 ),
    .Z(\V2/V4/V4/s2 [3]));
 OR2_X1 \V2/V4/V4/A2/M4/_0_  (.A1(\V2/V4/V4/A2/M4/c1 ),
    .A2(\V2/V4/V4/A2/M4/c2 ),
    .ZN(\V2/V4/V4/c2 ));
 AND2_X1 \V2/V4/V4/A3/M1/M1/_0_  (.A1(\V2/V4/V4/v4 [0]),
    .A2(\V2/V4/V4/s2 [2]),
    .ZN(\V2/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M1/M1/_1_  (.A(\V2/V4/V4/v4 [0]),
    .B(\V2/V4/V4/s2 [2]),
    .Z(\V2/V4/V4/A3/M1/s1 ));
 AND2_X1 \V2/V4/V4/A3/M1/M2/_0_  (.A1(\V2/V4/V4/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V2/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M1/M2/_1_  (.A(\V2/V4/V4/A3/M1/s1 ),
    .B(net6),
    .Z(\V2/V4/v4 [4]));
 OR2_X1 \V2/V4/V4/A3/M1/_0_  (.A1(\V2/V4/V4/A3/M1/c1 ),
    .A2(\V2/V4/V4/A3/M1/c2 ),
    .ZN(\V2/V4/V4/A3/c1 ));
 AND2_X1 \V2/V4/V4/A3/M2/M1/_0_  (.A1(\V2/V4/V4/v4 [1]),
    .A2(\V2/V4/V4/s2 [3]),
    .ZN(\V2/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M2/M1/_1_  (.A(\V2/V4/V4/v4 [1]),
    .B(\V2/V4/V4/s2 [3]),
    .Z(\V2/V4/V4/A3/M2/s1 ));
 AND2_X1 \V2/V4/V4/A3/M2/M2/_0_  (.A1(\V2/V4/V4/A3/M2/s1 ),
    .A2(\V2/V4/V4/A3/c1 ),
    .ZN(\V2/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M2/M2/_1_  (.A(\V2/V4/V4/A3/M2/s1 ),
    .B(\V2/V4/V4/A3/c1 ),
    .Z(\V2/V4/v4 [5]));
 OR2_X1 \V2/V4/V4/A3/M2/_0_  (.A1(\V2/V4/V4/A3/M2/c1 ),
    .A2(\V2/V4/V4/A3/M2/c2 ),
    .ZN(\V2/V4/V4/A3/c2 ));
 AND2_X1 \V2/V4/V4/A3/M3/M1/_0_  (.A1(\V2/V4/V4/v4 [2]),
    .A2(\V2/V4/V4/c3 ),
    .ZN(\V2/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M3/M1/_1_  (.A(\V2/V4/V4/v4 [2]),
    .B(\V2/V4/V4/c3 ),
    .Z(\V2/V4/V4/A3/M3/s1 ));
 AND2_X1 \V2/V4/V4/A3/M3/M2/_0_  (.A1(\V2/V4/V4/A3/M3/s1 ),
    .A2(\V2/V4/V4/A3/c2 ),
    .ZN(\V2/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M3/M2/_1_  (.A(\V2/V4/V4/A3/M3/s1 ),
    .B(\V2/V4/V4/A3/c2 ),
    .Z(\V2/V4/v4 [6]));
 OR2_X1 \V2/V4/V4/A3/M3/_0_  (.A1(\V2/V4/V4/A3/M3/c1 ),
    .A2(\V2/V4/V4/A3/M3/c2 ),
    .ZN(\V2/V4/V4/A3/c3 ));
 AND2_X1 \V2/V4/V4/A3/M4/M1/_0_  (.A1(\V2/V4/V4/v4 [3]),
    .A2(net6),
    .ZN(\V2/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V2/V4/V4/A3/M4/M1/_1_  (.A(\V2/V4/V4/v4 [3]),
    .B(net6),
    .Z(\V2/V4/V4/A3/M4/s1 ));
 AND2_X1 \V2/V4/V4/A3/M4/M2/_0_  (.A1(\V2/V4/V4/A3/M4/s1 ),
    .A2(\V2/V4/V4/A3/c3 ),
    .ZN(\V2/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V2/V4/V4/A3/M4/M2/_1_  (.A(\V2/V4/V4/A3/M4/s1 ),
    .B(\V2/V4/V4/A3/c3 ),
    .Z(\V2/V4/v4 [7]));
 OR2_X1 \V2/V4/V4/A3/M4/_0_  (.A1(\V2/V4/V4/A3/M4/c1 ),
    .A2(\V2/V4/V4/A3/M4/c2 ),
    .ZN(\V2/V4/V4/overflow ));
 AND2_X1 \V2/V4/V4/V1/HA1/_0_  (.A1(\V2/V4/V4/V1/w2 ),
    .A2(\V2/V4/V4/V1/w1 ),
    .ZN(\V2/V4/V4/V1/w4 ));
 XOR2_X2 \V2/V4/V4/V1/HA1/_1_  (.A(\V2/V4/V4/V1/w2 ),
    .B(\V2/V4/V4/V1/w1 ),
    .Z(\V2/V4/v4 [1]));
 AND2_X1 \V2/V4/V4/V1/HA2/_0_  (.A1(\V2/V4/V4/V1/w4 ),
    .A2(\V2/V4/V4/V1/w3 ),
    .ZN(\V2/V4/V4/v1 [3]));
 XOR2_X2 \V2/V4/V4/V1/HA2/_1_  (.A(\V2/V4/V4/V1/w4 ),
    .B(\V2/V4/V4/V1/w3 ),
    .Z(\V2/V4/V4/v1 [2]));
 AND2_X1 \V2/V4/V4/V1/_0_  (.A1(net29),
    .A2(B[12]),
    .ZN(\V2/V4/v4 [0]));
 AND2_X1 \V2/V4/V4/V1/_1_  (.A1(net29),
    .A2(B[13]),
    .ZN(\V2/V4/V4/V1/w1 ));
 AND2_X1 \V2/V4/V4/V1/_2_  (.A1(B[12]),
    .A2(net28),
    .ZN(\V2/V4/V4/V1/w2 ));
 AND2_X1 \V2/V4/V4/V1/_3_  (.A1(B[13]),
    .A2(net28),
    .ZN(\V2/V4/V4/V1/w3 ));
 AND2_X1 \V2/V4/V4/V2/HA1/_0_  (.A1(\V2/V4/V4/V2/w2 ),
    .A2(\V2/V4/V4/V2/w1 ),
    .ZN(\V2/V4/V4/V2/w4 ));
 XOR2_X2 \V2/V4/V4/V2/HA1/_1_  (.A(\V2/V4/V4/V2/w2 ),
    .B(\V2/V4/V4/V2/w1 ),
    .Z(\V2/V4/V4/v2 [1]));
 AND2_X1 \V2/V4/V4/V2/HA2/_0_  (.A1(\V2/V4/V4/V2/w4 ),
    .A2(\V2/V4/V4/V2/w3 ),
    .ZN(\V2/V4/V4/v2 [3]));
 XOR2_X2 \V2/V4/V4/V2/HA2/_1_  (.A(\V2/V4/V4/V2/w4 ),
    .B(\V2/V4/V4/V2/w3 ),
    .Z(\V2/V4/V4/v2 [2]));
 AND2_X1 \V2/V4/V4/V2/_0_  (.A1(net27),
    .A2(B[12]),
    .ZN(\V2/V4/V4/v2 [0]));
 AND2_X1 \V2/V4/V4/V2/_1_  (.A1(net27),
    .A2(B[13]),
    .ZN(\V2/V4/V4/V2/w1 ));
 AND2_X1 \V2/V4/V4/V2/_2_  (.A1(B[12]),
    .A2(net26),
    .ZN(\V2/V4/V4/V2/w2 ));
 AND2_X1 \V2/V4/V4/V2/_3_  (.A1(B[13]),
    .A2(net26),
    .ZN(\V2/V4/V4/V2/w3 ));
 AND2_X1 \V2/V4/V4/V3/HA1/_0_  (.A1(\V2/V4/V4/V3/w2 ),
    .A2(\V2/V4/V4/V3/w1 ),
    .ZN(\V2/V4/V4/V3/w4 ));
 XOR2_X2 \V2/V4/V4/V3/HA1/_1_  (.A(\V2/V4/V4/V3/w2 ),
    .B(\V2/V4/V4/V3/w1 ),
    .Z(\V2/V4/V4/v3 [1]));
 AND2_X1 \V2/V4/V4/V3/HA2/_0_  (.A1(\V2/V4/V4/V3/w4 ),
    .A2(\V2/V4/V4/V3/w3 ),
    .ZN(\V2/V4/V4/v3 [3]));
 XOR2_X2 \V2/V4/V4/V3/HA2/_1_  (.A(\V2/V4/V4/V3/w4 ),
    .B(\V2/V4/V4/V3/w3 ),
    .Z(\V2/V4/V4/v3 [2]));
 AND2_X1 \V2/V4/V4/V3/_0_  (.A1(net29),
    .A2(B[14]),
    .ZN(\V2/V4/V4/v3 [0]));
 AND2_X1 \V2/V4/V4/V3/_1_  (.A1(net29),
    .A2(B[15]),
    .ZN(\V2/V4/V4/V3/w1 ));
 AND2_X1 \V2/V4/V4/V3/_2_  (.A1(B[14]),
    .A2(net28),
    .ZN(\V2/V4/V4/V3/w2 ));
 AND2_X1 \V2/V4/V4/V3/_3_  (.A1(B[15]),
    .A2(net28),
    .ZN(\V2/V4/V4/V3/w3 ));
 AND2_X1 \V2/V4/V4/V4/HA1/_0_  (.A1(\V2/V4/V4/V4/w2 ),
    .A2(\V2/V4/V4/V4/w1 ),
    .ZN(\V2/V4/V4/V4/w4 ));
 XOR2_X2 \V2/V4/V4/V4/HA1/_1_  (.A(\V2/V4/V4/V4/w2 ),
    .B(\V2/V4/V4/V4/w1 ),
    .Z(\V2/V4/V4/v4 [1]));
 AND2_X1 \V2/V4/V4/V4/HA2/_0_  (.A1(\V2/V4/V4/V4/w4 ),
    .A2(\V2/V4/V4/V4/w3 ),
    .ZN(\V2/V4/V4/v4 [3]));
 XOR2_X2 \V2/V4/V4/V4/HA2/_1_  (.A(\V2/V4/V4/V4/w4 ),
    .B(\V2/V4/V4/V4/w3 ),
    .Z(\V2/V4/V4/v4 [2]));
 AND2_X1 \V2/V4/V4/V4/_0_  (.A1(net27),
    .A2(B[14]),
    .ZN(\V2/V4/V4/v4 [0]));
 AND2_X1 \V2/V4/V4/V4/_1_  (.A1(net27),
    .A2(B[15]),
    .ZN(\V2/V4/V4/V4/w1 ));
 AND2_X1 \V2/V4/V4/V4/_2_  (.A1(B[14]),
    .A2(net26),
    .ZN(\V2/V4/V4/V4/w2 ));
 AND2_X1 \V2/V4/V4/V4/_3_  (.A1(B[15]),
    .A2(net26),
    .ZN(\V2/V4/V4/V4/w3 ));
 OR2_X1 \V2/V4/V4/_0_  (.A1(\V2/V4/V4/c1 ),
    .A2(\V2/V4/V4/c2 ),
    .ZN(\V2/V4/V4/c3 ));
 OR2_X1 \V2/V4/_0_  (.A1(\V2/V4/c1 ),
    .A2(\V2/V4/c2 ),
    .ZN(\V2/V4/c3 ));
 OR2_X1 \V2/_0_  (.A1(\V2/c1 ),
    .A2(\V2/c2 ),
    .ZN(\V2/c3 ));
 AND2_X1 \V3/A1/A1/A1/M1/M1/_0_  (.A1(\V3/v2 [0]),
    .A2(\V3/v3 [0]),
    .ZN(\V3/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M1/M1/_1_  (.A(\V3/v2 [0]),
    .B(\V3/v3 [0]),
    .Z(\V3/A1/A1/A1/M1/s1 ));
 AND2_X1 \V3/A1/A1/A1/M1/M2/_0_  (.A1(\V3/A1/A1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M1/M2/_1_  (.A(\V3/A1/A1/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/s1 [0]));
 OR2_X1 \V3/A1/A1/A1/M1/_0_  (.A1(\V3/A1/A1/A1/M1/c1 ),
    .A2(\V3/A1/A1/A1/M1/c2 ),
    .ZN(\V3/A1/A1/A1/c1 ));
 AND2_X1 \V3/A1/A1/A1/M2/M1/_0_  (.A1(\V3/v2 [1]),
    .A2(\V3/v3 [1]),
    .ZN(\V3/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M2/M1/_1_  (.A(\V3/v2 [1]),
    .B(\V3/v3 [1]),
    .Z(\V3/A1/A1/A1/M2/s1 ));
 AND2_X1 \V3/A1/A1/A1/M2/M2/_0_  (.A1(\V3/A1/A1/A1/M2/s1 ),
    .A2(\V3/A1/A1/A1/c1 ),
    .ZN(\V3/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M2/M2/_1_  (.A(\V3/A1/A1/A1/M2/s1 ),
    .B(\V3/A1/A1/A1/c1 ),
    .Z(\V3/s1 [1]));
 OR2_X1 \V3/A1/A1/A1/M2/_0_  (.A1(\V3/A1/A1/A1/M2/c1 ),
    .A2(\V3/A1/A1/A1/M2/c2 ),
    .ZN(\V3/A1/A1/A1/c2 ));
 AND2_X1 \V3/A1/A1/A1/M3/M1/_0_  (.A1(\V3/v2 [2]),
    .A2(\V3/v3 [2]),
    .ZN(\V3/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M3/M1/_1_  (.A(\V3/v2 [2]),
    .B(\V3/v3 [2]),
    .Z(\V3/A1/A1/A1/M3/s1 ));
 AND2_X1 \V3/A1/A1/A1/M3/M2/_0_  (.A1(\V3/A1/A1/A1/M3/s1 ),
    .A2(\V3/A1/A1/A1/c2 ),
    .ZN(\V3/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M3/M2/_1_  (.A(\V3/A1/A1/A1/M3/s1 ),
    .B(\V3/A1/A1/A1/c2 ),
    .Z(\V3/s1 [2]));
 OR2_X1 \V3/A1/A1/A1/M3/_0_  (.A1(\V3/A1/A1/A1/M3/c1 ),
    .A2(\V3/A1/A1/A1/M3/c2 ),
    .ZN(\V3/A1/A1/A1/c3 ));
 AND2_X1 \V3/A1/A1/A1/M4/M1/_0_  (.A1(\V3/v2 [3]),
    .A2(\V3/v3 [3]),
    .ZN(\V3/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A1/A1/A1/M4/M1/_1_  (.A(\V3/v2 [3]),
    .B(\V3/v3 [3]),
    .Z(\V3/A1/A1/A1/M4/s1 ));
 AND2_X1 \V3/A1/A1/A1/M4/M2/_0_  (.A1(\V3/A1/A1/A1/M4/s1 ),
    .A2(\V3/A1/A1/A1/c3 ),
    .ZN(\V3/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A1/A1/A1/M4/M2/_1_  (.A(\V3/A1/A1/A1/M4/s1 ),
    .B(\V3/A1/A1/A1/c3 ),
    .Z(\V3/s1 [3]));
 OR2_X1 \V3/A1/A1/A1/M4/_0_  (.A1(\V3/A1/A1/A1/M4/c1 ),
    .A2(\V3/A1/A1/A1/M4/c2 ),
    .ZN(\V3/A1/A1/c1 ));
 AND2_X1 \V3/A1/A1/A2/M1/M1/_0_  (.A1(\V3/v2 [4]),
    .A2(\V3/v3 [4]),
    .ZN(\V3/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M1/M1/_1_  (.A(\V3/v2 [4]),
    .B(\V3/v3 [4]),
    .Z(\V3/A1/A1/A2/M1/s1 ));
 AND2_X1 \V3/A1/A1/A2/M1/M2/_0_  (.A1(\V3/A1/A1/A2/M1/s1 ),
    .A2(\V3/A1/A1/c1 ),
    .ZN(\V3/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M1/M2/_1_  (.A(\V3/A1/A1/A2/M1/s1 ),
    .B(\V3/A1/A1/c1 ),
    .Z(\V3/s1 [4]));
 OR2_X1 \V3/A1/A1/A2/M1/_0_  (.A1(\V3/A1/A1/A2/M1/c1 ),
    .A2(\V3/A1/A1/A2/M1/c2 ),
    .ZN(\V3/A1/A1/A2/c1 ));
 AND2_X1 \V3/A1/A1/A2/M2/M1/_0_  (.A1(\V3/v2 [5]),
    .A2(\V3/v3 [5]),
    .ZN(\V3/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M2/M1/_1_  (.A(\V3/v2 [5]),
    .B(\V3/v3 [5]),
    .Z(\V3/A1/A1/A2/M2/s1 ));
 AND2_X1 \V3/A1/A1/A2/M2/M2/_0_  (.A1(\V3/A1/A1/A2/M2/s1 ),
    .A2(\V3/A1/A1/A2/c1 ),
    .ZN(\V3/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M2/M2/_1_  (.A(\V3/A1/A1/A2/M2/s1 ),
    .B(\V3/A1/A1/A2/c1 ),
    .Z(\V3/s1 [5]));
 OR2_X1 \V3/A1/A1/A2/M2/_0_  (.A1(\V3/A1/A1/A2/M2/c1 ),
    .A2(\V3/A1/A1/A2/M2/c2 ),
    .ZN(\V3/A1/A1/A2/c2 ));
 AND2_X1 \V3/A1/A1/A2/M3/M1/_0_  (.A1(\V3/v2 [6]),
    .A2(\V3/v3 [6]),
    .ZN(\V3/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M3/M1/_1_  (.A(\V3/v2 [6]),
    .B(\V3/v3 [6]),
    .Z(\V3/A1/A1/A2/M3/s1 ));
 AND2_X1 \V3/A1/A1/A2/M3/M2/_0_  (.A1(\V3/A1/A1/A2/M3/s1 ),
    .A2(\V3/A1/A1/A2/c2 ),
    .ZN(\V3/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M3/M2/_1_  (.A(\V3/A1/A1/A2/M3/s1 ),
    .B(\V3/A1/A1/A2/c2 ),
    .Z(\V3/s1 [6]));
 OR2_X1 \V3/A1/A1/A2/M3/_0_  (.A1(\V3/A1/A1/A2/M3/c1 ),
    .A2(\V3/A1/A1/A2/M3/c2 ),
    .ZN(\V3/A1/A1/A2/c3 ));
 AND2_X1 \V3/A1/A1/A2/M4/M1/_0_  (.A1(\V3/v2 [7]),
    .A2(\V3/v3 [7]),
    .ZN(\V3/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A1/A1/A2/M4/M1/_1_  (.A(\V3/v2 [7]),
    .B(\V3/v3 [7]),
    .Z(\V3/A1/A1/A2/M4/s1 ));
 AND2_X1 \V3/A1/A1/A2/M4/M2/_0_  (.A1(\V3/A1/A1/A2/M4/s1 ),
    .A2(\V3/A1/A1/A2/c3 ),
    .ZN(\V3/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A1/A1/A2/M4/M2/_1_  (.A(\V3/A1/A1/A2/M4/s1 ),
    .B(\V3/A1/A1/A2/c3 ),
    .Z(\V3/s1 [7]));
 OR2_X1 \V3/A1/A1/A2/M4/_0_  (.A1(\V3/A1/A1/A2/M4/c1 ),
    .A2(\V3/A1/A1/A2/M4/c2 ),
    .ZN(\V3/A1/c1 ));
 AND2_X1 \V3/A1/A2/A1/M1/M1/_0_  (.A1(\V3/v2 [8]),
    .A2(\V3/v3 [8]),
    .ZN(\V3/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M1/M1/_1_  (.A(\V3/v2 [8]),
    .B(\V3/v3 [8]),
    .Z(\V3/A1/A2/A1/M1/s1 ));
 AND2_X1 \V3/A1/A2/A1/M1/M2/_0_  (.A1(\V3/A1/A2/A1/M1/s1 ),
    .A2(\V3/A1/c1 ),
    .ZN(\V3/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M1/M2/_1_  (.A(\V3/A1/A2/A1/M1/s1 ),
    .B(\V3/A1/c1 ),
    .Z(\V3/s1 [8]));
 OR2_X1 \V3/A1/A2/A1/M1/_0_  (.A1(\V3/A1/A2/A1/M1/c1 ),
    .A2(\V3/A1/A2/A1/M1/c2 ),
    .ZN(\V3/A1/A2/A1/c1 ));
 AND2_X1 \V3/A1/A2/A1/M2/M1/_0_  (.A1(\V3/v2 [9]),
    .A2(\V3/v3 [9]),
    .ZN(\V3/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M2/M1/_1_  (.A(\V3/v2 [9]),
    .B(\V3/v3 [9]),
    .Z(\V3/A1/A2/A1/M2/s1 ));
 AND2_X1 \V3/A1/A2/A1/M2/M2/_0_  (.A1(\V3/A1/A2/A1/M2/s1 ),
    .A2(\V3/A1/A2/A1/c1 ),
    .ZN(\V3/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M2/M2/_1_  (.A(\V3/A1/A2/A1/M2/s1 ),
    .B(\V3/A1/A2/A1/c1 ),
    .Z(\V3/s1 [9]));
 OR2_X1 \V3/A1/A2/A1/M2/_0_  (.A1(\V3/A1/A2/A1/M2/c1 ),
    .A2(\V3/A1/A2/A1/M2/c2 ),
    .ZN(\V3/A1/A2/A1/c2 ));
 AND2_X1 \V3/A1/A2/A1/M3/M1/_0_  (.A1(\V3/v2 [10]),
    .A2(\V3/v3 [10]),
    .ZN(\V3/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M3/M1/_1_  (.A(\V3/v2 [10]),
    .B(\V3/v3 [10]),
    .Z(\V3/A1/A2/A1/M3/s1 ));
 AND2_X1 \V3/A1/A2/A1/M3/M2/_0_  (.A1(\V3/A1/A2/A1/M3/s1 ),
    .A2(\V3/A1/A2/A1/c2 ),
    .ZN(\V3/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M3/M2/_1_  (.A(\V3/A1/A2/A1/M3/s1 ),
    .B(\V3/A1/A2/A1/c2 ),
    .Z(\V3/s1 [10]));
 OR2_X1 \V3/A1/A2/A1/M3/_0_  (.A1(\V3/A1/A2/A1/M3/c1 ),
    .A2(\V3/A1/A2/A1/M3/c2 ),
    .ZN(\V3/A1/A2/A1/c3 ));
 AND2_X1 \V3/A1/A2/A1/M4/M1/_0_  (.A1(\V3/v2 [11]),
    .A2(\V3/v3 [11]),
    .ZN(\V3/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A1/A2/A1/M4/M1/_1_  (.A(\V3/v2 [11]),
    .B(\V3/v3 [11]),
    .Z(\V3/A1/A2/A1/M4/s1 ));
 AND2_X1 \V3/A1/A2/A1/M4/M2/_0_  (.A1(\V3/A1/A2/A1/M4/s1 ),
    .A2(\V3/A1/A2/A1/c3 ),
    .ZN(\V3/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A1/A2/A1/M4/M2/_1_  (.A(\V3/A1/A2/A1/M4/s1 ),
    .B(\V3/A1/A2/A1/c3 ),
    .Z(\V3/s1 [11]));
 OR2_X1 \V3/A1/A2/A1/M4/_0_  (.A1(\V3/A1/A2/A1/M4/c1 ),
    .A2(\V3/A1/A2/A1/M4/c2 ),
    .ZN(\V3/A1/A2/c1 ));
 AND2_X1 \V3/A1/A2/A2/M1/M1/_0_  (.A1(\V3/v2 [12]),
    .A2(\V3/v3 [12]),
    .ZN(\V3/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M1/M1/_1_  (.A(\V3/v2 [12]),
    .B(\V3/v3 [12]),
    .Z(\V3/A1/A2/A2/M1/s1 ));
 AND2_X1 \V3/A1/A2/A2/M1/M2/_0_  (.A1(\V3/A1/A2/A2/M1/s1 ),
    .A2(\V3/A1/A2/c1 ),
    .ZN(\V3/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M1/M2/_1_  (.A(\V3/A1/A2/A2/M1/s1 ),
    .B(\V3/A1/A2/c1 ),
    .Z(\V3/s1 [12]));
 OR2_X1 \V3/A1/A2/A2/M1/_0_  (.A1(\V3/A1/A2/A2/M1/c1 ),
    .A2(\V3/A1/A2/A2/M1/c2 ),
    .ZN(\V3/A1/A2/A2/c1 ));
 AND2_X1 \V3/A1/A2/A2/M2/M1/_0_  (.A1(\V3/v2 [13]),
    .A2(\V3/v3 [13]),
    .ZN(\V3/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M2/M1/_1_  (.A(\V3/v2 [13]),
    .B(\V3/v3 [13]),
    .Z(\V3/A1/A2/A2/M2/s1 ));
 AND2_X1 \V3/A1/A2/A2/M2/M2/_0_  (.A1(\V3/A1/A2/A2/M2/s1 ),
    .A2(\V3/A1/A2/A2/c1 ),
    .ZN(\V3/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M2/M2/_1_  (.A(\V3/A1/A2/A2/M2/s1 ),
    .B(\V3/A1/A2/A2/c1 ),
    .Z(\V3/s1 [13]));
 OR2_X1 \V3/A1/A2/A2/M2/_0_  (.A1(\V3/A1/A2/A2/M2/c1 ),
    .A2(\V3/A1/A2/A2/M2/c2 ),
    .ZN(\V3/A1/A2/A2/c2 ));
 AND2_X1 \V3/A1/A2/A2/M3/M1/_0_  (.A1(\V3/v2 [14]),
    .A2(\V3/v3 [14]),
    .ZN(\V3/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M3/M1/_1_  (.A(\V3/v2 [14]),
    .B(\V3/v3 [14]),
    .Z(\V3/A1/A2/A2/M3/s1 ));
 AND2_X1 \V3/A1/A2/A2/M3/M2/_0_  (.A1(\V3/A1/A2/A2/M3/s1 ),
    .A2(\V3/A1/A2/A2/c2 ),
    .ZN(\V3/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M3/M2/_1_  (.A(\V3/A1/A2/A2/M3/s1 ),
    .B(\V3/A1/A2/A2/c2 ),
    .Z(\V3/s1 [14]));
 OR2_X1 \V3/A1/A2/A2/M3/_0_  (.A1(\V3/A1/A2/A2/M3/c1 ),
    .A2(\V3/A1/A2/A2/M3/c2 ),
    .ZN(\V3/A1/A2/A2/c3 ));
 AND2_X1 \V3/A1/A2/A2/M4/M1/_0_  (.A1(\V3/v2 [15]),
    .A2(\V3/v3 [15]),
    .ZN(\V3/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A1/A2/A2/M4/M1/_1_  (.A(\V3/v2 [15]),
    .B(\V3/v3 [15]),
    .Z(\V3/A1/A2/A2/M4/s1 ));
 AND2_X1 \V3/A1/A2/A2/M4/M2/_0_  (.A1(\V3/A1/A2/A2/M4/s1 ),
    .A2(\V3/A1/A2/A2/c3 ),
    .ZN(\V3/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A1/A2/A2/M4/M2/_1_  (.A(\V3/A1/A2/A2/M4/s1 ),
    .B(\V3/A1/A2/A2/c3 ),
    .Z(\V3/s1 [15]));
 OR2_X1 \V3/A1/A2/A2/M4/_0_  (.A1(\V3/A1/A2/A2/M4/c1 ),
    .A2(\V3/A1/A2/A2/M4/c2 ),
    .ZN(\V3/c1 ));
 AND2_X1 \V3/A2/A1/A1/M1/M1/_0_  (.A1(\V3/s1 [0]),
    .A2(\V3/v1 [8]),
    .ZN(\V3/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M1/M1/_1_  (.A(\V3/s1 [0]),
    .B(\V3/v1 [8]),
    .Z(\V3/A2/A1/A1/M1/s1 ));
 AND2_X1 \V3/A2/A1/A1/M1/M2/_0_  (.A1(\V3/A2/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M1/M2/_1_  (.A(\V3/A2/A1/A1/M1/s1 ),
    .B(net6),
    .Z(v3[8]));
 OR2_X1 \V3/A2/A1/A1/M1/_0_  (.A1(\V3/A2/A1/A1/M1/c1 ),
    .A2(\V3/A2/A1/A1/M1/c2 ),
    .ZN(\V3/A2/A1/A1/c1 ));
 AND2_X1 \V3/A2/A1/A1/M2/M1/_0_  (.A1(\V3/s1 [1]),
    .A2(\V3/v1 [9]),
    .ZN(\V3/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M2/M1/_1_  (.A(\V3/s1 [1]),
    .B(\V3/v1 [9]),
    .Z(\V3/A2/A1/A1/M2/s1 ));
 AND2_X1 \V3/A2/A1/A1/M2/M2/_0_  (.A1(\V3/A2/A1/A1/M2/s1 ),
    .A2(\V3/A2/A1/A1/c1 ),
    .ZN(\V3/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M2/M2/_1_  (.A(\V3/A2/A1/A1/M2/s1 ),
    .B(\V3/A2/A1/A1/c1 ),
    .Z(v3[9]));
 OR2_X1 \V3/A2/A1/A1/M2/_0_  (.A1(\V3/A2/A1/A1/M2/c1 ),
    .A2(\V3/A2/A1/A1/M2/c2 ),
    .ZN(\V3/A2/A1/A1/c2 ));
 AND2_X1 \V3/A2/A1/A1/M3/M1/_0_  (.A1(\V3/s1 [2]),
    .A2(\V3/v1 [10]),
    .ZN(\V3/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M3/M1/_1_  (.A(\V3/s1 [2]),
    .B(\V3/v1 [10]),
    .Z(\V3/A2/A1/A1/M3/s1 ));
 AND2_X1 \V3/A2/A1/A1/M3/M2/_0_  (.A1(\V3/A2/A1/A1/M3/s1 ),
    .A2(\V3/A2/A1/A1/c2 ),
    .ZN(\V3/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M3/M2/_1_  (.A(\V3/A2/A1/A1/M3/s1 ),
    .B(\V3/A2/A1/A1/c2 ),
    .Z(v3[10]));
 OR2_X1 \V3/A2/A1/A1/M3/_0_  (.A1(\V3/A2/A1/A1/M3/c1 ),
    .A2(\V3/A2/A1/A1/M3/c2 ),
    .ZN(\V3/A2/A1/A1/c3 ));
 AND2_X1 \V3/A2/A1/A1/M4/M1/_0_  (.A1(\V3/s1 [3]),
    .A2(\V3/v1 [11]),
    .ZN(\V3/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A2/A1/A1/M4/M1/_1_  (.A(\V3/s1 [3]),
    .B(\V3/v1 [11]),
    .Z(\V3/A2/A1/A1/M4/s1 ));
 AND2_X1 \V3/A2/A1/A1/M4/M2/_0_  (.A1(\V3/A2/A1/A1/M4/s1 ),
    .A2(\V3/A2/A1/A1/c3 ),
    .ZN(\V3/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A2/A1/A1/M4/M2/_1_  (.A(\V3/A2/A1/A1/M4/s1 ),
    .B(\V3/A2/A1/A1/c3 ),
    .Z(v3[11]));
 OR2_X1 \V3/A2/A1/A1/M4/_0_  (.A1(\V3/A2/A1/A1/M4/c1 ),
    .A2(\V3/A2/A1/A1/M4/c2 ),
    .ZN(\V3/A2/A1/c1 ));
 AND2_X1 \V3/A2/A1/A2/M1/M1/_0_  (.A1(\V3/s1 [4]),
    .A2(\V3/v1 [12]),
    .ZN(\V3/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M1/M1/_1_  (.A(\V3/s1 [4]),
    .B(\V3/v1 [12]),
    .Z(\V3/A2/A1/A2/M1/s1 ));
 AND2_X1 \V3/A2/A1/A2/M1/M2/_0_  (.A1(\V3/A2/A1/A2/M1/s1 ),
    .A2(\V3/A2/A1/c1 ),
    .ZN(\V3/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M1/M2/_1_  (.A(\V3/A2/A1/A2/M1/s1 ),
    .B(\V3/A2/A1/c1 ),
    .Z(v3[12]));
 OR2_X1 \V3/A2/A1/A2/M1/_0_  (.A1(\V3/A2/A1/A2/M1/c1 ),
    .A2(\V3/A2/A1/A2/M1/c2 ),
    .ZN(\V3/A2/A1/A2/c1 ));
 AND2_X1 \V3/A2/A1/A2/M2/M1/_0_  (.A1(\V3/s1 [5]),
    .A2(\V3/v1 [13]),
    .ZN(\V3/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M2/M1/_1_  (.A(\V3/s1 [5]),
    .B(\V3/v1 [13]),
    .Z(\V3/A2/A1/A2/M2/s1 ));
 AND2_X1 \V3/A2/A1/A2/M2/M2/_0_  (.A1(\V3/A2/A1/A2/M2/s1 ),
    .A2(\V3/A2/A1/A2/c1 ),
    .ZN(\V3/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M2/M2/_1_  (.A(\V3/A2/A1/A2/M2/s1 ),
    .B(\V3/A2/A1/A2/c1 ),
    .Z(v3[13]));
 OR2_X1 \V3/A2/A1/A2/M2/_0_  (.A1(\V3/A2/A1/A2/M2/c1 ),
    .A2(\V3/A2/A1/A2/M2/c2 ),
    .ZN(\V3/A2/A1/A2/c2 ));
 AND2_X1 \V3/A2/A1/A2/M3/M1/_0_  (.A1(\V3/s1 [6]),
    .A2(\V3/v1 [14]),
    .ZN(\V3/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M3/M1/_1_  (.A(\V3/s1 [6]),
    .B(\V3/v1 [14]),
    .Z(\V3/A2/A1/A2/M3/s1 ));
 AND2_X1 \V3/A2/A1/A2/M3/M2/_0_  (.A1(\V3/A2/A1/A2/M3/s1 ),
    .A2(\V3/A2/A1/A2/c2 ),
    .ZN(\V3/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M3/M2/_1_  (.A(\V3/A2/A1/A2/M3/s1 ),
    .B(\V3/A2/A1/A2/c2 ),
    .Z(v3[14]));
 OR2_X1 \V3/A2/A1/A2/M3/_0_  (.A1(\V3/A2/A1/A2/M3/c1 ),
    .A2(\V3/A2/A1/A2/M3/c2 ),
    .ZN(\V3/A2/A1/A2/c3 ));
 AND2_X1 \V3/A2/A1/A2/M4/M1/_0_  (.A1(\V3/s1 [7]),
    .A2(\V3/v1 [15]),
    .ZN(\V3/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A2/A1/A2/M4/M1/_1_  (.A(\V3/s1 [7]),
    .B(\V3/v1 [15]),
    .Z(\V3/A2/A1/A2/M4/s1 ));
 AND2_X1 \V3/A2/A1/A2/M4/M2/_0_  (.A1(\V3/A2/A1/A2/M4/s1 ),
    .A2(\V3/A2/A1/A2/c3 ),
    .ZN(\V3/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A2/A1/A2/M4/M2/_1_  (.A(\V3/A2/A1/A2/M4/s1 ),
    .B(\V3/A2/A1/A2/c3 ),
    .Z(v3[15]));
 OR2_X2 \V3/A2/A1/A2/M4/_0_  (.A1(\V3/A2/A1/A2/M4/c1 ),
    .A2(\V3/A2/A1/A2/M4/c2 ),
    .ZN(\V3/A2/c1 ));
 AND2_X1 \V3/A2/A2/A1/M1/M1/_0_  (.A1(\V3/s1 [8]),
    .A2(net6),
    .ZN(\V3/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M1/M1/_1_  (.A(\V3/s1 [8]),
    .B(net6),
    .Z(\V3/A2/A2/A1/M1/s1 ));
 AND2_X1 \V3/A2/A2/A1/M1/M2/_0_  (.A1(\V3/A2/A2/A1/M1/s1 ),
    .A2(\V3/A2/c1 ),
    .ZN(\V3/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M1/M2/_1_  (.A(\V3/A2/A2/A1/M1/s1 ),
    .B(\V3/A2/c1 ),
    .Z(\V3/s2 [8]));
 OR2_X1 \V3/A2/A2/A1/M1/_0_  (.A1(\V3/A2/A2/A1/M1/c1 ),
    .A2(\V3/A2/A2/A1/M1/c2 ),
    .ZN(\V3/A2/A2/A1/c1 ));
 AND2_X1 \V3/A2/A2/A1/M2/M1/_0_  (.A1(\V3/s1 [9]),
    .A2(net6),
    .ZN(\V3/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M2/M1/_1_  (.A(\V3/s1 [9]),
    .B(net6),
    .Z(\V3/A2/A2/A1/M2/s1 ));
 AND2_X1 \V3/A2/A2/A1/M2/M2/_0_  (.A1(\V3/A2/A2/A1/M2/s1 ),
    .A2(\V3/A2/A2/A1/c1 ),
    .ZN(\V3/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M2/M2/_1_  (.A(\V3/A2/A2/A1/M2/s1 ),
    .B(\V3/A2/A2/A1/c1 ),
    .Z(\V3/s2 [9]));
 OR2_X1 \V3/A2/A2/A1/M2/_0_  (.A1(\V3/A2/A2/A1/M2/c1 ),
    .A2(\V3/A2/A2/A1/M2/c2 ),
    .ZN(\V3/A2/A2/A1/c2 ));
 AND2_X1 \V3/A2/A2/A1/M3/M1/_0_  (.A1(\V3/s1 [10]),
    .A2(net6),
    .ZN(\V3/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M3/M1/_1_  (.A(\V3/s1 [10]),
    .B(net6),
    .Z(\V3/A2/A2/A1/M3/s1 ));
 AND2_X1 \V3/A2/A2/A1/M3/M2/_0_  (.A1(\V3/A2/A2/A1/M3/s1 ),
    .A2(\V3/A2/A2/A1/c2 ),
    .ZN(\V3/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M3/M2/_1_  (.A(\V3/A2/A2/A1/M3/s1 ),
    .B(\V3/A2/A2/A1/c2 ),
    .Z(\V3/s2 [10]));
 OR2_X1 \V3/A2/A2/A1/M3/_0_  (.A1(\V3/A2/A2/A1/M3/c1 ),
    .A2(\V3/A2/A2/A1/M3/c2 ),
    .ZN(\V3/A2/A2/A1/c3 ));
 AND2_X1 \V3/A2/A2/A1/M4/M1/_0_  (.A1(\V3/s1 [11]),
    .A2(net6),
    .ZN(\V3/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A2/A2/A1/M4/M1/_1_  (.A(\V3/s1 [11]),
    .B(net6),
    .Z(\V3/A2/A2/A1/M4/s1 ));
 AND2_X1 \V3/A2/A2/A1/M4/M2/_0_  (.A1(\V3/A2/A2/A1/M4/s1 ),
    .A2(\V3/A2/A2/A1/c3 ),
    .ZN(\V3/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A2/A2/A1/M4/M2/_1_  (.A(\V3/A2/A2/A1/M4/s1 ),
    .B(\V3/A2/A2/A1/c3 ),
    .Z(\V3/s2 [11]));
 OR2_X1 \V3/A2/A2/A1/M4/_0_  (.A1(\V3/A2/A2/A1/M4/c1 ),
    .A2(\V3/A2/A2/A1/M4/c2 ),
    .ZN(\V3/A2/A2/c1 ));
 AND2_X1 \V3/A2/A2/A2/M1/M1/_0_  (.A1(\V3/s1 [12]),
    .A2(net5),
    .ZN(\V3/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M1/M1/_1_  (.A(\V3/s1 [12]),
    .B(net5),
    .Z(\V3/A2/A2/A2/M1/s1 ));
 AND2_X1 \V3/A2/A2/A2/M1/M2/_0_  (.A1(\V3/A2/A2/A2/M1/s1 ),
    .A2(\V3/A2/A2/c1 ),
    .ZN(\V3/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M1/M2/_1_  (.A(\V3/A2/A2/A2/M1/s1 ),
    .B(\V3/A2/A2/c1 ),
    .Z(\V3/s2 [12]));
 OR2_X1 \V3/A2/A2/A2/M1/_0_  (.A1(\V3/A2/A2/A2/M1/c1 ),
    .A2(\V3/A2/A2/A2/M1/c2 ),
    .ZN(\V3/A2/A2/A2/c1 ));
 AND2_X1 \V3/A2/A2/A2/M2/M1/_0_  (.A1(\V3/s1 [13]),
    .A2(net8),
    .ZN(\V3/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M2/M1/_1_  (.A(\V3/s1 [13]),
    .B(net8),
    .Z(\V3/A2/A2/A2/M2/s1 ));
 AND2_X1 \V3/A2/A2/A2/M2/M2/_0_  (.A1(\V3/A2/A2/A2/M2/s1 ),
    .A2(\V3/A2/A2/A2/c1 ),
    .ZN(\V3/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M2/M2/_1_  (.A(\V3/A2/A2/A2/M2/s1 ),
    .B(\V3/A2/A2/A2/c1 ),
    .Z(\V3/s2 [13]));
 OR2_X1 \V3/A2/A2/A2/M2/_0_  (.A1(\V3/A2/A2/A2/M2/c1 ),
    .A2(\V3/A2/A2/A2/M2/c2 ),
    .ZN(\V3/A2/A2/A2/c2 ));
 AND2_X1 \V3/A2/A2/A2/M3/M1/_0_  (.A1(\V3/s1 [14]),
    .A2(net8),
    .ZN(\V3/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M3/M1/_1_  (.A(\V3/s1 [14]),
    .B(net8),
    .Z(\V3/A2/A2/A2/M3/s1 ));
 AND2_X1 \V3/A2/A2/A2/M3/M2/_0_  (.A1(\V3/A2/A2/A2/M3/s1 ),
    .A2(\V3/A2/A2/A2/c2 ),
    .ZN(\V3/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M3/M2/_1_  (.A(\V3/A2/A2/A2/M3/s1 ),
    .B(\V3/A2/A2/A2/c2 ),
    .Z(\V3/s2 [14]));
 OR2_X1 \V3/A2/A2/A2/M3/_0_  (.A1(\V3/A2/A2/A2/M3/c1 ),
    .A2(\V3/A2/A2/A2/M3/c2 ),
    .ZN(\V3/A2/A2/A2/c3 ));
 AND2_X1 \V3/A2/A2/A2/M4/M1/_0_  (.A1(\V3/s1 [15]),
    .A2(net8),
    .ZN(\V3/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A2/A2/A2/M4/M1/_1_  (.A(\V3/s1 [15]),
    .B(net8),
    .Z(\V3/A2/A2/A2/M4/s1 ));
 AND2_X1 \V3/A2/A2/A2/M4/M2/_0_  (.A1(\V3/A2/A2/A2/M4/s1 ),
    .A2(\V3/A2/A2/A2/c3 ),
    .ZN(\V3/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A2/A2/A2/M4/M2/_1_  (.A(\V3/A2/A2/A2/M4/s1 ),
    .B(\V3/A2/A2/A2/c3 ),
    .Z(\V3/s2 [15]));
 OR2_X1 \V3/A2/A2/A2/M4/_0_  (.A1(\V3/A2/A2/A2/M4/c1 ),
    .A2(\V3/A2/A2/A2/M4/c2 ),
    .ZN(\V3/c2 ));
 AND2_X1 \V3/A3/A1/A1/M1/M1/_0_  (.A1(\V3/v4 [0]),
    .A2(\V3/s2 [8]),
    .ZN(\V3/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M1/M1/_1_  (.A(\V3/v4 [0]),
    .B(\V3/s2 [8]),
    .Z(\V3/A3/A1/A1/M1/s1 ));
 AND2_X1 \V3/A3/A1/A1/M1/M2/_0_  (.A1(\V3/A3/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M1/M2/_1_  (.A(\V3/A3/A1/A1/M1/s1 ),
    .B(net6),
    .Z(v3[16]));
 OR2_X1 \V3/A3/A1/A1/M1/_0_  (.A1(\V3/A3/A1/A1/M1/c1 ),
    .A2(\V3/A3/A1/A1/M1/c2 ),
    .ZN(\V3/A3/A1/A1/c1 ));
 AND2_X1 \V3/A3/A1/A1/M2/M1/_0_  (.A1(\V3/v4 [1]),
    .A2(\V3/s2 [9]),
    .ZN(\V3/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M2/M1/_1_  (.A(\V3/v4 [1]),
    .B(\V3/s2 [9]),
    .Z(\V3/A3/A1/A1/M2/s1 ));
 AND2_X1 \V3/A3/A1/A1/M2/M2/_0_  (.A1(\V3/A3/A1/A1/M2/s1 ),
    .A2(\V3/A3/A1/A1/c1 ),
    .ZN(\V3/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M2/M2/_1_  (.A(\V3/A3/A1/A1/M2/s1 ),
    .B(\V3/A3/A1/A1/c1 ),
    .Z(v3[17]));
 OR2_X1 \V3/A3/A1/A1/M2/_0_  (.A1(\V3/A3/A1/A1/M2/c1 ),
    .A2(\V3/A3/A1/A1/M2/c2 ),
    .ZN(\V3/A3/A1/A1/c2 ));
 AND2_X1 \V3/A3/A1/A1/M3/M1/_0_  (.A1(\V3/v4 [2]),
    .A2(\V3/s2 [10]),
    .ZN(\V3/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M3/M1/_1_  (.A(\V3/v4 [2]),
    .B(\V3/s2 [10]),
    .Z(\V3/A3/A1/A1/M3/s1 ));
 AND2_X1 \V3/A3/A1/A1/M3/M2/_0_  (.A1(\V3/A3/A1/A1/M3/s1 ),
    .A2(\V3/A3/A1/A1/c2 ),
    .ZN(\V3/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M3/M2/_1_  (.A(\V3/A3/A1/A1/M3/s1 ),
    .B(\V3/A3/A1/A1/c2 ),
    .Z(v3[18]));
 OR2_X1 \V3/A3/A1/A1/M3/_0_  (.A1(\V3/A3/A1/A1/M3/c1 ),
    .A2(\V3/A3/A1/A1/M3/c2 ),
    .ZN(\V3/A3/A1/A1/c3 ));
 AND2_X1 \V3/A3/A1/A1/M4/M1/_0_  (.A1(\V3/v4 [3]),
    .A2(\V3/s2 [11]),
    .ZN(\V3/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V3/A3/A1/A1/M4/M1/_1_  (.A(\V3/v4 [3]),
    .B(\V3/s2 [11]),
    .Z(\V3/A3/A1/A1/M4/s1 ));
 AND2_X1 \V3/A3/A1/A1/M4/M2/_0_  (.A1(\V3/A3/A1/A1/M4/s1 ),
    .A2(\V3/A3/A1/A1/c3 ),
    .ZN(\V3/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V3/A3/A1/A1/M4/M2/_1_  (.A(\V3/A3/A1/A1/M4/s1 ),
    .B(\V3/A3/A1/A1/c3 ),
    .Z(v3[19]));
 OR2_X1 \V3/A3/A1/A1/M4/_0_  (.A1(\V3/A3/A1/A1/M4/c1 ),
    .A2(\V3/A3/A1/A1/M4/c2 ),
    .ZN(\V3/A3/A1/c1 ));
 AND2_X1 \V3/A3/A1/A2/M1/M1/_0_  (.A1(\V3/v4 [4]),
    .A2(\V3/s2 [12]),
    .ZN(\V3/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M1/M1/_1_  (.A(\V3/v4 [4]),
    .B(\V3/s2 [12]),
    .Z(\V3/A3/A1/A2/M1/s1 ));
 AND2_X1 \V3/A3/A1/A2/M1/M2/_0_  (.A1(\V3/A3/A1/A2/M1/s1 ),
    .A2(\V3/A3/A1/c1 ),
    .ZN(\V3/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M1/M2/_1_  (.A(\V3/A3/A1/A2/M1/s1 ),
    .B(\V3/A3/A1/c1 ),
    .Z(v3[20]));
 OR2_X1 \V3/A3/A1/A2/M1/_0_  (.A1(\V3/A3/A1/A2/M1/c1 ),
    .A2(\V3/A3/A1/A2/M1/c2 ),
    .ZN(\V3/A3/A1/A2/c1 ));
 AND2_X1 \V3/A3/A1/A2/M2/M1/_0_  (.A1(\V3/v4 [5]),
    .A2(\V3/s2 [13]),
    .ZN(\V3/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M2/M1/_1_  (.A(\V3/v4 [5]),
    .B(\V3/s2 [13]),
    .Z(\V3/A3/A1/A2/M2/s1 ));
 AND2_X1 \V3/A3/A1/A2/M2/M2/_0_  (.A1(\V3/A3/A1/A2/M2/s1 ),
    .A2(\V3/A3/A1/A2/c1 ),
    .ZN(\V3/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M2/M2/_1_  (.A(\V3/A3/A1/A2/M2/s1 ),
    .B(\V3/A3/A1/A2/c1 ),
    .Z(v3[21]));
 OR2_X1 \V3/A3/A1/A2/M2/_0_  (.A1(\V3/A3/A1/A2/M2/c1 ),
    .A2(\V3/A3/A1/A2/M2/c2 ),
    .ZN(\V3/A3/A1/A2/c2 ));
 AND2_X1 \V3/A3/A1/A2/M3/M1/_0_  (.A1(\V3/v4 [6]),
    .A2(\V3/s2 [14]),
    .ZN(\V3/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M3/M1/_1_  (.A(\V3/v4 [6]),
    .B(\V3/s2 [14]),
    .Z(\V3/A3/A1/A2/M3/s1 ));
 AND2_X1 \V3/A3/A1/A2/M3/M2/_0_  (.A1(\V3/A3/A1/A2/M3/s1 ),
    .A2(\V3/A3/A1/A2/c2 ),
    .ZN(\V3/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M3/M2/_1_  (.A(\V3/A3/A1/A2/M3/s1 ),
    .B(\V3/A3/A1/A2/c2 ),
    .Z(v3[22]));
 OR2_X1 \V3/A3/A1/A2/M3/_0_  (.A1(\V3/A3/A1/A2/M3/c1 ),
    .A2(\V3/A3/A1/A2/M3/c2 ),
    .ZN(\V3/A3/A1/A2/c3 ));
 AND2_X1 \V3/A3/A1/A2/M4/M1/_0_  (.A1(\V3/v4 [7]),
    .A2(\V3/s2 [15]),
    .ZN(\V3/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V3/A3/A1/A2/M4/M1/_1_  (.A(\V3/v4 [7]),
    .B(\V3/s2 [15]),
    .Z(\V3/A3/A1/A2/M4/s1 ));
 AND2_X1 \V3/A3/A1/A2/M4/M2/_0_  (.A1(\V3/A3/A1/A2/M4/s1 ),
    .A2(\V3/A3/A1/A2/c3 ),
    .ZN(\V3/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V3/A3/A1/A2/M4/M2/_1_  (.A(\V3/A3/A1/A2/M4/s1 ),
    .B(\V3/A3/A1/A2/c3 ),
    .Z(v3[23]));
 OR2_X1 \V3/A3/A1/A2/M4/_0_  (.A1(\V3/A3/A1/A2/M4/c1 ),
    .A2(\V3/A3/A1/A2/M4/c2 ),
    .ZN(\V3/A3/c1 ));
 AND2_X1 \V3/A3/A2/A1/M1/M1/_0_  (.A1(\V3/v4 [8]),
    .A2(\V3/c3 ),
    .ZN(\V3/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M1/M1/_1_  (.A(\V3/v4 [8]),
    .B(\V3/c3 ),
    .Z(\V3/A3/A2/A1/M1/s1 ));
 AND2_X1 \V3/A3/A2/A1/M1/M2/_0_  (.A1(\V3/A3/A2/A1/M1/s1 ),
    .A2(\V3/A3/c1 ),
    .ZN(\V3/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M1/M2/_1_  (.A(\V3/A3/A2/A1/M1/s1 ),
    .B(\V3/A3/c1 ),
    .Z(v3[24]));
 OR2_X1 \V3/A3/A2/A1/M1/_0_  (.A1(\V3/A3/A2/A1/M1/c1 ),
    .A2(\V3/A3/A2/A1/M1/c2 ),
    .ZN(\V3/A3/A2/A1/c1 ));
 AND2_X1 \V3/A3/A2/A1/M2/M1/_0_  (.A1(\V3/v4 [9]),
    .A2(net6),
    .ZN(\V3/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M2/M1/_1_  (.A(\V3/v4 [9]),
    .B(net6),
    .Z(\V3/A3/A2/A1/M2/s1 ));
 AND2_X1 \V3/A3/A2/A1/M2/M2/_0_  (.A1(\V3/A3/A2/A1/M2/s1 ),
    .A2(\V3/A3/A2/A1/c1 ),
    .ZN(\V3/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M2/M2/_1_  (.A(\V3/A3/A2/A1/M2/s1 ),
    .B(\V3/A3/A2/A1/c1 ),
    .Z(v3[25]));
 OR2_X1 \V3/A3/A2/A1/M2/_0_  (.A1(\V3/A3/A2/A1/M2/c1 ),
    .A2(\V3/A3/A2/A1/M2/c2 ),
    .ZN(\V3/A3/A2/A1/c2 ));
 AND2_X1 \V3/A3/A2/A1/M3/M1/_0_  (.A1(\V3/v4 [10]),
    .A2(net6),
    .ZN(\V3/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M3/M1/_1_  (.A(\V3/v4 [10]),
    .B(net6),
    .Z(\V3/A3/A2/A1/M3/s1 ));
 AND2_X1 \V3/A3/A2/A1/M3/M2/_0_  (.A1(\V3/A3/A2/A1/M3/s1 ),
    .A2(\V3/A3/A2/A1/c2 ),
    .ZN(\V3/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M3/M2/_1_  (.A(\V3/A3/A2/A1/M3/s1 ),
    .B(\V3/A3/A2/A1/c2 ),
    .Z(v3[26]));
 OR2_X1 \V3/A3/A2/A1/M3/_0_  (.A1(\V3/A3/A2/A1/M3/c1 ),
    .A2(\V3/A3/A2/A1/M3/c2 ),
    .ZN(\V3/A3/A2/A1/c3 ));
 AND2_X1 \V3/A3/A2/A1/M4/M1/_0_  (.A1(\V3/v4 [11]),
    .A2(net6),
    .ZN(\V3/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V3/A3/A2/A1/M4/M1/_1_  (.A(\V3/v4 [11]),
    .B(net6),
    .Z(\V3/A3/A2/A1/M4/s1 ));
 AND2_X1 \V3/A3/A2/A1/M4/M2/_0_  (.A1(\V3/A3/A2/A1/M4/s1 ),
    .A2(\V3/A3/A2/A1/c3 ),
    .ZN(\V3/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V3/A3/A2/A1/M4/M2/_1_  (.A(\V3/A3/A2/A1/M4/s1 ),
    .B(\V3/A3/A2/A1/c3 ),
    .Z(v3[27]));
 OR2_X1 \V3/A3/A2/A1/M4/_0_  (.A1(\V3/A3/A2/A1/M4/c1 ),
    .A2(\V3/A3/A2/A1/M4/c2 ),
    .ZN(\V3/A3/A2/c1 ));
 AND2_X1 \V3/A3/A2/A2/M1/M1/_0_  (.A1(\V3/v4 [12]),
    .A2(net7),
    .ZN(\V3/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M1/M1/_1_  (.A(\V3/v4 [12]),
    .B(net7),
    .Z(\V3/A3/A2/A2/M1/s1 ));
 AND2_X1 \V3/A3/A2/A2/M1/M2/_0_  (.A1(\V3/A3/A2/A2/M1/s1 ),
    .A2(\V3/A3/A2/c1 ),
    .ZN(\V3/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M1/M2/_1_  (.A(\V3/A3/A2/A2/M1/s1 ),
    .B(\V3/A3/A2/c1 ),
    .Z(v3[28]));
 OR2_X1 \V3/A3/A2/A2/M1/_0_  (.A1(\V3/A3/A2/A2/M1/c1 ),
    .A2(\V3/A3/A2/A2/M1/c2 ),
    .ZN(\V3/A3/A2/A2/c1 ));
 AND2_X1 \V3/A3/A2/A2/M2/M1/_0_  (.A1(\V3/v4 [13]),
    .A2(net7),
    .ZN(\V3/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M2/M1/_1_  (.A(\V3/v4 [13]),
    .B(net7),
    .Z(\V3/A3/A2/A2/M2/s1 ));
 AND2_X1 \V3/A3/A2/A2/M2/M2/_0_  (.A1(\V3/A3/A2/A2/M2/s1 ),
    .A2(\V3/A3/A2/A2/c1 ),
    .ZN(\V3/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M2/M2/_1_  (.A(\V3/A3/A2/A2/M2/s1 ),
    .B(\V3/A3/A2/A2/c1 ),
    .Z(v3[29]));
 OR2_X1 \V3/A3/A2/A2/M2/_0_  (.A1(\V3/A3/A2/A2/M2/c1 ),
    .A2(\V3/A3/A2/A2/M2/c2 ),
    .ZN(\V3/A3/A2/A2/c2 ));
 AND2_X1 \V3/A3/A2/A2/M3/M1/_0_  (.A1(\V3/v4 [14]),
    .A2(net7),
    .ZN(\V3/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M3/M1/_1_  (.A(\V3/v4 [14]),
    .B(net7),
    .Z(\V3/A3/A2/A2/M3/s1 ));
 AND2_X1 \V3/A3/A2/A2/M3/M2/_0_  (.A1(\V3/A3/A2/A2/M3/s1 ),
    .A2(\V3/A3/A2/A2/c2 ),
    .ZN(\V3/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M3/M2/_1_  (.A(\V3/A3/A2/A2/M3/s1 ),
    .B(\V3/A3/A2/A2/c2 ),
    .Z(v3[30]));
 OR2_X1 \V3/A3/A2/A2/M3/_0_  (.A1(\V3/A3/A2/A2/M3/c1 ),
    .A2(\V3/A3/A2/A2/M3/c2 ),
    .ZN(\V3/A3/A2/A2/c3 ));
 AND2_X1 \V3/A3/A2/A2/M4/M1/_0_  (.A1(\V3/v4 [15]),
    .A2(net7),
    .ZN(\V3/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V3/A3/A2/A2/M4/M1/_1_  (.A(\V3/v4 [15]),
    .B(net7),
    .Z(\V3/A3/A2/A2/M4/s1 ));
 AND2_X1 \V3/A3/A2/A2/M4/M2/_0_  (.A1(\V3/A3/A2/A2/M4/s1 ),
    .A2(\V3/A3/A2/A2/c3 ),
    .ZN(\V3/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V3/A3/A2/A2/M4/M2/_1_  (.A(\V3/A3/A2/A2/M4/s1 ),
    .B(\V3/A3/A2/A2/c3 ),
    .Z(v3[31]));
 OR2_X1 \V3/A3/A2/A2/M4/_0_  (.A1(\V3/A3/A2/A2/M4/c1 ),
    .A2(\V3/A3/A2/A2/M4/c2 ),
    .ZN(\V3/overflow ));
 AND2_X1 \V3/V1/A1/A1/M1/M1/_0_  (.A1(\V3/V1/v2 [0]),
    .A2(\V3/V1/v3 [0]),
    .ZN(\V3/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M1/M1/_1_  (.A(\V3/V1/v2 [0]),
    .B(\V3/V1/v3 [0]),
    .Z(\V3/V1/A1/A1/M1/s1 ));
 AND2_X1 \V3/V1/A1/A1/M1/M2/_0_  (.A1(\V3/V1/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M1/M2/_1_  (.A(\V3/V1/A1/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/V1/s1 [0]));
 OR2_X1 \V3/V1/A1/A1/M1/_0_  (.A1(\V3/V1/A1/A1/M1/c1 ),
    .A2(\V3/V1/A1/A1/M1/c2 ),
    .ZN(\V3/V1/A1/A1/c1 ));
 AND2_X1 \V3/V1/A1/A1/M2/M1/_0_  (.A1(\V3/V1/v2 [1]),
    .A2(\V3/V1/v3 [1]),
    .ZN(\V3/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M2/M1/_1_  (.A(\V3/V1/v2 [1]),
    .B(\V3/V1/v3 [1]),
    .Z(\V3/V1/A1/A1/M2/s1 ));
 AND2_X1 \V3/V1/A1/A1/M2/M2/_0_  (.A1(\V3/V1/A1/A1/M2/s1 ),
    .A2(\V3/V1/A1/A1/c1 ),
    .ZN(\V3/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M2/M2/_1_  (.A(\V3/V1/A1/A1/M2/s1 ),
    .B(\V3/V1/A1/A1/c1 ),
    .Z(\V3/V1/s1 [1]));
 OR2_X1 \V3/V1/A1/A1/M2/_0_  (.A1(\V3/V1/A1/A1/M2/c1 ),
    .A2(\V3/V1/A1/A1/M2/c2 ),
    .ZN(\V3/V1/A1/A1/c2 ));
 AND2_X1 \V3/V1/A1/A1/M3/M1/_0_  (.A1(\V3/V1/v2 [2]),
    .A2(\V3/V1/v3 [2]),
    .ZN(\V3/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M3/M1/_1_  (.A(\V3/V1/v2 [2]),
    .B(\V3/V1/v3 [2]),
    .Z(\V3/V1/A1/A1/M3/s1 ));
 AND2_X1 \V3/V1/A1/A1/M3/M2/_0_  (.A1(\V3/V1/A1/A1/M3/s1 ),
    .A2(\V3/V1/A1/A1/c2 ),
    .ZN(\V3/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M3/M2/_1_  (.A(\V3/V1/A1/A1/M3/s1 ),
    .B(\V3/V1/A1/A1/c2 ),
    .Z(\V3/V1/s1 [2]));
 OR2_X1 \V3/V1/A1/A1/M3/_0_  (.A1(\V3/V1/A1/A1/M3/c1 ),
    .A2(\V3/V1/A1/A1/M3/c2 ),
    .ZN(\V3/V1/A1/A1/c3 ));
 AND2_X1 \V3/V1/A1/A1/M4/M1/_0_  (.A1(\V3/V1/v2 [3]),
    .A2(\V3/V1/v3 [3]),
    .ZN(\V3/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A1/A1/M4/M1/_1_  (.A(\V3/V1/v2 [3]),
    .B(\V3/V1/v3 [3]),
    .Z(\V3/V1/A1/A1/M4/s1 ));
 AND2_X1 \V3/V1/A1/A1/M4/M2/_0_  (.A1(\V3/V1/A1/A1/M4/s1 ),
    .A2(\V3/V1/A1/A1/c3 ),
    .ZN(\V3/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A1/A1/M4/M2/_1_  (.A(\V3/V1/A1/A1/M4/s1 ),
    .B(\V3/V1/A1/A1/c3 ),
    .Z(\V3/V1/s1 [3]));
 OR2_X1 \V3/V1/A1/A1/M4/_0_  (.A1(\V3/V1/A1/A1/M4/c1 ),
    .A2(\V3/V1/A1/A1/M4/c2 ),
    .ZN(\V3/V1/A1/c1 ));
 AND2_X1 \V3/V1/A1/A2/M1/M1/_0_  (.A1(\V3/V1/v2 [4]),
    .A2(\V3/V1/v3 [4]),
    .ZN(\V3/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M1/M1/_1_  (.A(\V3/V1/v2 [4]),
    .B(\V3/V1/v3 [4]),
    .Z(\V3/V1/A1/A2/M1/s1 ));
 AND2_X1 \V3/V1/A1/A2/M1/M2/_0_  (.A1(\V3/V1/A1/A2/M1/s1 ),
    .A2(\V3/V1/A1/c1 ),
    .ZN(\V3/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M1/M2/_1_  (.A(\V3/V1/A1/A2/M1/s1 ),
    .B(\V3/V1/A1/c1 ),
    .Z(\V3/V1/s1 [4]));
 OR2_X1 \V3/V1/A1/A2/M1/_0_  (.A1(\V3/V1/A1/A2/M1/c1 ),
    .A2(\V3/V1/A1/A2/M1/c2 ),
    .ZN(\V3/V1/A1/A2/c1 ));
 AND2_X1 \V3/V1/A1/A2/M2/M1/_0_  (.A1(\V3/V1/v2 [5]),
    .A2(\V3/V1/v3 [5]),
    .ZN(\V3/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M2/M1/_1_  (.A(\V3/V1/v2 [5]),
    .B(\V3/V1/v3 [5]),
    .Z(\V3/V1/A1/A2/M2/s1 ));
 AND2_X1 \V3/V1/A1/A2/M2/M2/_0_  (.A1(\V3/V1/A1/A2/M2/s1 ),
    .A2(\V3/V1/A1/A2/c1 ),
    .ZN(\V3/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M2/M2/_1_  (.A(\V3/V1/A1/A2/M2/s1 ),
    .B(\V3/V1/A1/A2/c1 ),
    .Z(\V3/V1/s1 [5]));
 OR2_X1 \V3/V1/A1/A2/M2/_0_  (.A1(\V3/V1/A1/A2/M2/c1 ),
    .A2(\V3/V1/A1/A2/M2/c2 ),
    .ZN(\V3/V1/A1/A2/c2 ));
 AND2_X1 \V3/V1/A1/A2/M3/M1/_0_  (.A1(\V3/V1/v2 [6]),
    .A2(\V3/V1/v3 [6]),
    .ZN(\V3/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M3/M1/_1_  (.A(\V3/V1/v2 [6]),
    .B(\V3/V1/v3 [6]),
    .Z(\V3/V1/A1/A2/M3/s1 ));
 AND2_X1 \V3/V1/A1/A2/M3/M2/_0_  (.A1(\V3/V1/A1/A2/M3/s1 ),
    .A2(\V3/V1/A1/A2/c2 ),
    .ZN(\V3/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M3/M2/_1_  (.A(\V3/V1/A1/A2/M3/s1 ),
    .B(\V3/V1/A1/A2/c2 ),
    .Z(\V3/V1/s1 [6]));
 OR2_X1 \V3/V1/A1/A2/M3/_0_  (.A1(\V3/V1/A1/A2/M3/c1 ),
    .A2(\V3/V1/A1/A2/M3/c2 ),
    .ZN(\V3/V1/A1/A2/c3 ));
 AND2_X1 \V3/V1/A1/A2/M4/M1/_0_  (.A1(\V3/V1/v2 [7]),
    .A2(\V3/V1/v3 [7]),
    .ZN(\V3/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A1/A2/M4/M1/_1_  (.A(\V3/V1/v2 [7]),
    .B(\V3/V1/v3 [7]),
    .Z(\V3/V1/A1/A2/M4/s1 ));
 AND2_X1 \V3/V1/A1/A2/M4/M2/_0_  (.A1(\V3/V1/A1/A2/M4/s1 ),
    .A2(\V3/V1/A1/A2/c3 ),
    .ZN(\V3/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A1/A2/M4/M2/_1_  (.A(\V3/V1/A1/A2/M4/s1 ),
    .B(\V3/V1/A1/A2/c3 ),
    .Z(\V3/V1/s1 [7]));
 OR2_X1 \V3/V1/A1/A2/M4/_0_  (.A1(\V3/V1/A1/A2/M4/c1 ),
    .A2(\V3/V1/A1/A2/M4/c2 ),
    .ZN(\V3/V1/c1 ));
 AND2_X1 \V3/V1/A2/A1/M1/M1/_0_  (.A1(\V3/V1/s1 [0]),
    .A2(\V3/V1/v1 [4]),
    .ZN(\V3/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M1/M1/_1_  (.A(\V3/V1/s1 [0]),
    .B(\V3/V1/v1 [4]),
    .Z(\V3/V1/A2/A1/M1/s1 ));
 AND2_X1 \V3/V1/A2/A1/M1/M2/_0_  (.A1(\V3/V1/A2/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M1/M2/_1_  (.A(\V3/V1/A2/A1/M1/s1 ),
    .B(net4),
    .Z(v3[4]));
 OR2_X1 \V3/V1/A2/A1/M1/_0_  (.A1(\V3/V1/A2/A1/M1/c1 ),
    .A2(\V3/V1/A2/A1/M1/c2 ),
    .ZN(\V3/V1/A2/A1/c1 ));
 AND2_X1 \V3/V1/A2/A1/M2/M1/_0_  (.A1(\V3/V1/s1 [1]),
    .A2(\V3/V1/v1 [5]),
    .ZN(\V3/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M2/M1/_1_  (.A(\V3/V1/s1 [1]),
    .B(\V3/V1/v1 [5]),
    .Z(\V3/V1/A2/A1/M2/s1 ));
 AND2_X1 \V3/V1/A2/A1/M2/M2/_0_  (.A1(\V3/V1/A2/A1/M2/s1 ),
    .A2(\V3/V1/A2/A1/c1 ),
    .ZN(\V3/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M2/M2/_1_  (.A(\V3/V1/A2/A1/M2/s1 ),
    .B(\V3/V1/A2/A1/c1 ),
    .Z(v3[5]));
 OR2_X1 \V3/V1/A2/A1/M2/_0_  (.A1(\V3/V1/A2/A1/M2/c1 ),
    .A2(\V3/V1/A2/A1/M2/c2 ),
    .ZN(\V3/V1/A2/A1/c2 ));
 AND2_X1 \V3/V1/A2/A1/M3/M1/_0_  (.A1(\V3/V1/s1 [2]),
    .A2(\V3/V1/v1 [6]),
    .ZN(\V3/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M3/M1/_1_  (.A(\V3/V1/s1 [2]),
    .B(\V3/V1/v1 [6]),
    .Z(\V3/V1/A2/A1/M3/s1 ));
 AND2_X1 \V3/V1/A2/A1/M3/M2/_0_  (.A1(\V3/V1/A2/A1/M3/s1 ),
    .A2(\V3/V1/A2/A1/c2 ),
    .ZN(\V3/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M3/M2/_1_  (.A(\V3/V1/A2/A1/M3/s1 ),
    .B(\V3/V1/A2/A1/c2 ),
    .Z(v3[6]));
 OR2_X1 \V3/V1/A2/A1/M3/_0_  (.A1(\V3/V1/A2/A1/M3/c1 ),
    .A2(\V3/V1/A2/A1/M3/c2 ),
    .ZN(\V3/V1/A2/A1/c3 ));
 AND2_X1 \V3/V1/A2/A1/M4/M1/_0_  (.A1(\V3/V1/s1 [3]),
    .A2(\V3/V1/v1 [7]),
    .ZN(\V3/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A2/A1/M4/M1/_1_  (.A(\V3/V1/s1 [3]),
    .B(\V3/V1/v1 [7]),
    .Z(\V3/V1/A2/A1/M4/s1 ));
 AND2_X1 \V3/V1/A2/A1/M4/M2/_0_  (.A1(\V3/V1/A2/A1/M4/s1 ),
    .A2(\V3/V1/A2/A1/c3 ),
    .ZN(\V3/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A2/A1/M4/M2/_1_  (.A(\V3/V1/A2/A1/M4/s1 ),
    .B(\V3/V1/A2/A1/c3 ),
    .Z(v3[7]));
 OR2_X1 \V3/V1/A2/A1/M4/_0_  (.A1(\V3/V1/A2/A1/M4/c1 ),
    .A2(\V3/V1/A2/A1/M4/c2 ),
    .ZN(\V3/V1/A2/c1 ));
 AND2_X1 \V3/V1/A2/A2/M1/M1/_0_  (.A1(\V3/V1/s1 [4]),
    .A2(net2),
    .ZN(\V3/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M1/M1/_1_  (.A(\V3/V1/s1 [4]),
    .B(net2),
    .Z(\V3/V1/A2/A2/M1/s1 ));
 AND2_X1 \V3/V1/A2/A2/M1/M2/_0_  (.A1(\V3/V1/A2/A2/M1/s1 ),
    .A2(\V3/V1/A2/c1 ),
    .ZN(\V3/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M1/M2/_1_  (.A(\V3/V1/A2/A2/M1/s1 ),
    .B(\V3/V1/A2/c1 ),
    .Z(\V3/V1/s2 [4]));
 OR2_X1 \V3/V1/A2/A2/M1/_0_  (.A1(\V3/V1/A2/A2/M1/c1 ),
    .A2(\V3/V1/A2/A2/M1/c2 ),
    .ZN(\V3/V1/A2/A2/c1 ));
 AND2_X1 \V3/V1/A2/A2/M2/M1/_0_  (.A1(\V3/V1/s1 [5]),
    .A2(net2),
    .ZN(\V3/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M2/M1/_1_  (.A(\V3/V1/s1 [5]),
    .B(net2),
    .Z(\V3/V1/A2/A2/M2/s1 ));
 AND2_X1 \V3/V1/A2/A2/M2/M2/_0_  (.A1(\V3/V1/A2/A2/M2/s1 ),
    .A2(\V3/V1/A2/A2/c1 ),
    .ZN(\V3/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M2/M2/_1_  (.A(\V3/V1/A2/A2/M2/s1 ),
    .B(\V3/V1/A2/A2/c1 ),
    .Z(\V3/V1/s2 [5]));
 OR2_X1 \V3/V1/A2/A2/M2/_0_  (.A1(\V3/V1/A2/A2/M2/c1 ),
    .A2(\V3/V1/A2/A2/M2/c2 ),
    .ZN(\V3/V1/A2/A2/c2 ));
 AND2_X1 \V3/V1/A2/A2/M3/M1/_0_  (.A1(\V3/V1/s1 [6]),
    .A2(net2),
    .ZN(\V3/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M3/M1/_1_  (.A(\V3/V1/s1 [6]),
    .B(net2),
    .Z(\V3/V1/A2/A2/M3/s1 ));
 AND2_X1 \V3/V1/A2/A2/M3/M2/_0_  (.A1(\V3/V1/A2/A2/M3/s1 ),
    .A2(\V3/V1/A2/A2/c2 ),
    .ZN(\V3/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M3/M2/_1_  (.A(\V3/V1/A2/A2/M3/s1 ),
    .B(\V3/V1/A2/A2/c2 ),
    .Z(\V3/V1/s2 [6]));
 OR2_X1 \V3/V1/A2/A2/M3/_0_  (.A1(\V3/V1/A2/A2/M3/c1 ),
    .A2(\V3/V1/A2/A2/M3/c2 ),
    .ZN(\V3/V1/A2/A2/c3 ));
 AND2_X1 \V3/V1/A2/A2/M4/M1/_0_  (.A1(\V3/V1/s1 [7]),
    .A2(net2),
    .ZN(\V3/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A2/A2/M4/M1/_1_  (.A(\V3/V1/s1 [7]),
    .B(net2),
    .Z(\V3/V1/A2/A2/M4/s1 ));
 AND2_X1 \V3/V1/A2/A2/M4/M2/_0_  (.A1(\V3/V1/A2/A2/M4/s1 ),
    .A2(\V3/V1/A2/A2/c3 ),
    .ZN(\V3/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A2/A2/M4/M2/_1_  (.A(\V3/V1/A2/A2/M4/s1 ),
    .B(\V3/V1/A2/A2/c3 ),
    .Z(\V3/V1/s2 [7]));
 OR2_X1 \V3/V1/A2/A2/M4/_0_  (.A1(\V3/V1/A2/A2/M4/c1 ),
    .A2(\V3/V1/A2/A2/M4/c2 ),
    .ZN(\V3/V1/c2 ));
 AND2_X1 \V3/V1/A3/A1/M1/M1/_0_  (.A1(\V3/V1/v4 [0]),
    .A2(\V3/V1/s2 [4]),
    .ZN(\V3/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M1/M1/_1_  (.A(\V3/V1/v4 [0]),
    .B(\V3/V1/s2 [4]),
    .Z(\V3/V1/A3/A1/M1/s1 ));
 AND2_X1 \V3/V1/A3/A1/M1/M2/_0_  (.A1(\V3/V1/A3/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M1/M2/_1_  (.A(\V3/V1/A3/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/v1 [8]));
 OR2_X1 \V3/V1/A3/A1/M1/_0_  (.A1(\V3/V1/A3/A1/M1/c1 ),
    .A2(\V3/V1/A3/A1/M1/c2 ),
    .ZN(\V3/V1/A3/A1/c1 ));
 AND2_X1 \V3/V1/A3/A1/M2/M1/_0_  (.A1(\V3/V1/v4 [1]),
    .A2(\V3/V1/s2 [5]),
    .ZN(\V3/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M2/M1/_1_  (.A(\V3/V1/v4 [1]),
    .B(\V3/V1/s2 [5]),
    .Z(\V3/V1/A3/A1/M2/s1 ));
 AND2_X1 \V3/V1/A3/A1/M2/M2/_0_  (.A1(\V3/V1/A3/A1/M2/s1 ),
    .A2(\V3/V1/A3/A1/c1 ),
    .ZN(\V3/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M2/M2/_1_  (.A(\V3/V1/A3/A1/M2/s1 ),
    .B(\V3/V1/A3/A1/c1 ),
    .Z(\V3/v1 [9]));
 OR2_X1 \V3/V1/A3/A1/M2/_0_  (.A1(\V3/V1/A3/A1/M2/c1 ),
    .A2(\V3/V1/A3/A1/M2/c2 ),
    .ZN(\V3/V1/A3/A1/c2 ));
 AND2_X1 \V3/V1/A3/A1/M3/M1/_0_  (.A1(\V3/V1/v4 [2]),
    .A2(\V3/V1/s2 [6]),
    .ZN(\V3/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M3/M1/_1_  (.A(\V3/V1/v4 [2]),
    .B(\V3/V1/s2 [6]),
    .Z(\V3/V1/A3/A1/M3/s1 ));
 AND2_X1 \V3/V1/A3/A1/M3/M2/_0_  (.A1(\V3/V1/A3/A1/M3/s1 ),
    .A2(\V3/V1/A3/A1/c2 ),
    .ZN(\V3/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M3/M2/_1_  (.A(\V3/V1/A3/A1/M3/s1 ),
    .B(\V3/V1/A3/A1/c2 ),
    .Z(\V3/v1 [10]));
 OR2_X1 \V3/V1/A3/A1/M3/_0_  (.A1(\V3/V1/A3/A1/M3/c1 ),
    .A2(\V3/V1/A3/A1/M3/c2 ),
    .ZN(\V3/V1/A3/A1/c3 ));
 AND2_X1 \V3/V1/A3/A1/M4/M1/_0_  (.A1(\V3/V1/v4 [3]),
    .A2(\V3/V1/s2 [7]),
    .ZN(\V3/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V1/A3/A1/M4/M1/_1_  (.A(\V3/V1/v4 [3]),
    .B(\V3/V1/s2 [7]),
    .Z(\V3/V1/A3/A1/M4/s1 ));
 AND2_X1 \V3/V1/A3/A1/M4/M2/_0_  (.A1(\V3/V1/A3/A1/M4/s1 ),
    .A2(\V3/V1/A3/A1/c3 ),
    .ZN(\V3/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V1/A3/A1/M4/M2/_1_  (.A(\V3/V1/A3/A1/M4/s1 ),
    .B(\V3/V1/A3/A1/c3 ),
    .Z(\V3/v1 [11]));
 OR2_X1 \V3/V1/A3/A1/M4/_0_  (.A1(\V3/V1/A3/A1/M4/c1 ),
    .A2(\V3/V1/A3/A1/M4/c2 ),
    .ZN(\V3/V1/A3/c1 ));
 AND2_X1 \V3/V1/A3/A2/M1/M1/_0_  (.A1(\V3/V1/v4 [4]),
    .A2(\V3/V1/c3 ),
    .ZN(\V3/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M1/M1/_1_  (.A(\V3/V1/v4 [4]),
    .B(\V3/V1/c3 ),
    .Z(\V3/V1/A3/A2/M1/s1 ));
 AND2_X1 \V3/V1/A3/A2/M1/M2/_0_  (.A1(\V3/V1/A3/A2/M1/s1 ),
    .A2(\V3/V1/A3/c1 ),
    .ZN(\V3/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M1/M2/_1_  (.A(\V3/V1/A3/A2/M1/s1 ),
    .B(\V3/V1/A3/c1 ),
    .Z(\V3/v1 [12]));
 OR2_X1 \V3/V1/A3/A2/M1/_0_  (.A1(\V3/V1/A3/A2/M1/c1 ),
    .A2(\V3/V1/A3/A2/M1/c2 ),
    .ZN(\V3/V1/A3/A2/c1 ));
 AND2_X1 \V3/V1/A3/A2/M2/M1/_0_  (.A1(\V3/V1/v4 [5]),
    .A2(net2),
    .ZN(\V3/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M2/M1/_1_  (.A(\V3/V1/v4 [5]),
    .B(net2),
    .Z(\V3/V1/A3/A2/M2/s1 ));
 AND2_X1 \V3/V1/A3/A2/M2/M2/_0_  (.A1(\V3/V1/A3/A2/M2/s1 ),
    .A2(\V3/V1/A3/A2/c1 ),
    .ZN(\V3/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M2/M2/_1_  (.A(\V3/V1/A3/A2/M2/s1 ),
    .B(\V3/V1/A3/A2/c1 ),
    .Z(\V3/v1 [13]));
 OR2_X1 \V3/V1/A3/A2/M2/_0_  (.A1(\V3/V1/A3/A2/M2/c1 ),
    .A2(\V3/V1/A3/A2/M2/c2 ),
    .ZN(\V3/V1/A3/A2/c2 ));
 AND2_X1 \V3/V1/A3/A2/M3/M1/_0_  (.A1(\V3/V1/v4 [6]),
    .A2(net2),
    .ZN(\V3/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M3/M1/_1_  (.A(\V3/V1/v4 [6]),
    .B(net2),
    .Z(\V3/V1/A3/A2/M3/s1 ));
 AND2_X1 \V3/V1/A3/A2/M3/M2/_0_  (.A1(\V3/V1/A3/A2/M3/s1 ),
    .A2(\V3/V1/A3/A2/c2 ),
    .ZN(\V3/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M3/M2/_1_  (.A(\V3/V1/A3/A2/M3/s1 ),
    .B(\V3/V1/A3/A2/c2 ),
    .Z(\V3/v1 [14]));
 OR2_X1 \V3/V1/A3/A2/M3/_0_  (.A1(\V3/V1/A3/A2/M3/c1 ),
    .A2(\V3/V1/A3/A2/M3/c2 ),
    .ZN(\V3/V1/A3/A2/c3 ));
 AND2_X1 \V3/V1/A3/A2/M4/M1/_0_  (.A1(\V3/V1/v4 [7]),
    .A2(net2),
    .ZN(\V3/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V1/A3/A2/M4/M1/_1_  (.A(\V3/V1/v4 [7]),
    .B(net2),
    .Z(\V3/V1/A3/A2/M4/s1 ));
 AND2_X1 \V3/V1/A3/A2/M4/M2/_0_  (.A1(\V3/V1/A3/A2/M4/s1 ),
    .A2(\V3/V1/A3/A2/c3 ),
    .ZN(\V3/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V1/A3/A2/M4/M2/_1_  (.A(\V3/V1/A3/A2/M4/s1 ),
    .B(\V3/V1/A3/A2/c3 ),
    .Z(\V3/v1 [15]));
 OR2_X1 \V3/V1/A3/A2/M4/_0_  (.A1(\V3/V1/A3/A2/M4/c1 ),
    .A2(\V3/V1/A3/A2/M4/c2 ),
    .ZN(\V3/V1/overflow ));
 AND2_X1 \V3/V1/V1/A1/M1/M1/_0_  (.A1(\V3/V1/V1/v2 [0]),
    .A2(\V3/V1/V1/v3 [0]),
    .ZN(\V3/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M1/M1/_1_  (.A(\V3/V1/V1/v2 [0]),
    .B(\V3/V1/V1/v3 [0]),
    .Z(\V3/V1/V1/A1/M1/s1 ));
 AND2_X1 \V3/V1/V1/A1/M1/M2/_0_  (.A1(\V3/V1/V1/A1/M1/s1 ),
    .A2(net4),
    .ZN(\V3/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M1/M2/_1_  (.A(\V3/V1/V1/A1/M1/s1 ),
    .B(net4),
    .Z(\V3/V1/V1/s1 [0]));
 OR2_X1 \V3/V1/V1/A1/M1/_0_  (.A1(\V3/V1/V1/A1/M1/c1 ),
    .A2(\V3/V1/V1/A1/M1/c2 ),
    .ZN(\V3/V1/V1/A1/c1 ));
 AND2_X1 \V3/V1/V1/A1/M2/M1/_0_  (.A1(\V3/V1/V1/v2 [1]),
    .A2(\V3/V1/V1/v3 [1]),
    .ZN(\V3/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M2/M1/_1_  (.A(\V3/V1/V1/v2 [1]),
    .B(\V3/V1/V1/v3 [1]),
    .Z(\V3/V1/V1/A1/M2/s1 ));
 AND2_X1 \V3/V1/V1/A1/M2/M2/_0_  (.A1(\V3/V1/V1/A1/M2/s1 ),
    .A2(\V3/V1/V1/A1/c1 ),
    .ZN(\V3/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M2/M2/_1_  (.A(\V3/V1/V1/A1/M2/s1 ),
    .B(\V3/V1/V1/A1/c1 ),
    .Z(\V3/V1/V1/s1 [1]));
 OR2_X1 \V3/V1/V1/A1/M2/_0_  (.A1(\V3/V1/V1/A1/M2/c1 ),
    .A2(\V3/V1/V1/A1/M2/c2 ),
    .ZN(\V3/V1/V1/A1/c2 ));
 AND2_X1 \V3/V1/V1/A1/M3/M1/_0_  (.A1(\V3/V1/V1/v2 [2]),
    .A2(\V3/V1/V1/v3 [2]),
    .ZN(\V3/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M3/M1/_1_  (.A(\V3/V1/V1/v2 [2]),
    .B(\V3/V1/V1/v3 [2]),
    .Z(\V3/V1/V1/A1/M3/s1 ));
 AND2_X1 \V3/V1/V1/A1/M3/M2/_0_  (.A1(\V3/V1/V1/A1/M3/s1 ),
    .A2(\V3/V1/V1/A1/c2 ),
    .ZN(\V3/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M3/M2/_1_  (.A(\V3/V1/V1/A1/M3/s1 ),
    .B(\V3/V1/V1/A1/c2 ),
    .Z(\V3/V1/V1/s1 [2]));
 OR2_X1 \V3/V1/V1/A1/M3/_0_  (.A1(\V3/V1/V1/A1/M3/c1 ),
    .A2(\V3/V1/V1/A1/M3/c2 ),
    .ZN(\V3/V1/V1/A1/c3 ));
 AND2_X1 \V3/V1/V1/A1/M4/M1/_0_  (.A1(\V3/V1/V1/v2 [3]),
    .A2(\V3/V1/V1/v3 [3]),
    .ZN(\V3/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A1/M4/M1/_1_  (.A(\V3/V1/V1/v2 [3]),
    .B(\V3/V1/V1/v3 [3]),
    .Z(\V3/V1/V1/A1/M4/s1 ));
 AND2_X1 \V3/V1/V1/A1/M4/M2/_0_  (.A1(\V3/V1/V1/A1/M4/s1 ),
    .A2(\V3/V1/V1/A1/c3 ),
    .ZN(\V3/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A1/M4/M2/_1_  (.A(\V3/V1/V1/A1/M4/s1 ),
    .B(\V3/V1/V1/A1/c3 ),
    .Z(\V3/V1/V1/s1 [3]));
 OR2_X1 \V3/V1/V1/A1/M4/_0_  (.A1(\V3/V1/V1/A1/M4/c1 ),
    .A2(\V3/V1/V1/A1/M4/c2 ),
    .ZN(\V3/V1/V1/c1 ));
 AND2_X1 \V3/V1/V1/A2/M1/M1/_0_  (.A1(\V3/V1/V1/s1 [0]),
    .A2(\V3/V1/V1/v1 [2]),
    .ZN(\V3/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M1/M1/_1_  (.A(\V3/V1/V1/s1 [0]),
    .B(\V3/V1/V1/v1 [2]),
    .Z(\V3/V1/V1/A2/M1/s1 ));
 AND2_X1 \V3/V1/V1/A2/M1/M2/_0_  (.A1(\V3/V1/V1/A2/M1/s1 ),
    .A2(net4),
    .ZN(\V3/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M1/M2/_1_  (.A(\V3/V1/V1/A2/M1/s1 ),
    .B(net4),
    .Z(v3[2]));
 OR2_X1 \V3/V1/V1/A2/M1/_0_  (.A1(\V3/V1/V1/A2/M1/c1 ),
    .A2(\V3/V1/V1/A2/M1/c2 ),
    .ZN(\V3/V1/V1/A2/c1 ));
 AND2_X1 \V3/V1/V1/A2/M2/M1/_0_  (.A1(\V3/V1/V1/s1 [1]),
    .A2(\V3/V1/V1/v1 [3]),
    .ZN(\V3/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M2/M1/_1_  (.A(\V3/V1/V1/s1 [1]),
    .B(\V3/V1/V1/v1 [3]),
    .Z(\V3/V1/V1/A2/M2/s1 ));
 AND2_X1 \V3/V1/V1/A2/M2/M2/_0_  (.A1(\V3/V1/V1/A2/M2/s1 ),
    .A2(\V3/V1/V1/A2/c1 ),
    .ZN(\V3/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M2/M2/_1_  (.A(\V3/V1/V1/A2/M2/s1 ),
    .B(\V3/V1/V1/A2/c1 ),
    .Z(v3[3]));
 OR2_X1 \V3/V1/V1/A2/M2/_0_  (.A1(\V3/V1/V1/A2/M2/c1 ),
    .A2(\V3/V1/V1/A2/M2/c2 ),
    .ZN(\V3/V1/V1/A2/c2 ));
 AND2_X1 \V3/V1/V1/A2/M3/M1/_0_  (.A1(\V3/V1/V1/s1 [2]),
    .A2(net6),
    .ZN(\V3/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M3/M1/_1_  (.A(\V3/V1/V1/s1 [2]),
    .B(net6),
    .Z(\V3/V1/V1/A2/M3/s1 ));
 AND2_X1 \V3/V1/V1/A2/M3/M2/_0_  (.A1(\V3/V1/V1/A2/M3/s1 ),
    .A2(\V3/V1/V1/A2/c2 ),
    .ZN(\V3/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M3/M2/_1_  (.A(\V3/V1/V1/A2/M3/s1 ),
    .B(\V3/V1/V1/A2/c2 ),
    .Z(\V3/V1/V1/s2 [2]));
 OR2_X1 \V3/V1/V1/A2/M3/_0_  (.A1(\V3/V1/V1/A2/M3/c1 ),
    .A2(\V3/V1/V1/A2/M3/c2 ),
    .ZN(\V3/V1/V1/A2/c3 ));
 AND2_X1 \V3/V1/V1/A2/M4/M1/_0_  (.A1(\V3/V1/V1/s1 [3]),
    .A2(net6),
    .ZN(\V3/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A2/M4/M1/_1_  (.A(\V3/V1/V1/s1 [3]),
    .B(net6),
    .Z(\V3/V1/V1/A2/M4/s1 ));
 AND2_X1 \V3/V1/V1/A2/M4/M2/_0_  (.A1(\V3/V1/V1/A2/M4/s1 ),
    .A2(\V3/V1/V1/A2/c3 ),
    .ZN(\V3/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A2/M4/M2/_1_  (.A(\V3/V1/V1/A2/M4/s1 ),
    .B(\V3/V1/V1/A2/c3 ),
    .Z(\V3/V1/V1/s2 [3]));
 OR2_X1 \V3/V1/V1/A2/M4/_0_  (.A1(\V3/V1/V1/A2/M4/c1 ),
    .A2(\V3/V1/V1/A2/M4/c2 ),
    .ZN(\V3/V1/V1/c2 ));
 AND2_X1 \V3/V1/V1/A3/M1/M1/_0_  (.A1(\V3/V1/V1/v4 [0]),
    .A2(\V3/V1/V1/s2 [2]),
    .ZN(\V3/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M1/M1/_1_  (.A(\V3/V1/V1/v4 [0]),
    .B(\V3/V1/V1/s2 [2]),
    .Z(\V3/V1/V1/A3/M1/s1 ));
 AND2_X1 \V3/V1/V1/A3/M1/M2/_0_  (.A1(\V3/V1/V1/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M1/M2/_1_  (.A(\V3/V1/V1/A3/M1/s1 ),
    .B(net6),
    .Z(\V3/V1/v1 [4]));
 OR2_X1 \V3/V1/V1/A3/M1/_0_  (.A1(\V3/V1/V1/A3/M1/c1 ),
    .A2(\V3/V1/V1/A3/M1/c2 ),
    .ZN(\V3/V1/V1/A3/c1 ));
 AND2_X1 \V3/V1/V1/A3/M2/M1/_0_  (.A1(\V3/V1/V1/v4 [1]),
    .A2(\V3/V1/V1/s2 [3]),
    .ZN(\V3/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M2/M1/_1_  (.A(\V3/V1/V1/v4 [1]),
    .B(\V3/V1/V1/s2 [3]),
    .Z(\V3/V1/V1/A3/M2/s1 ));
 AND2_X1 \V3/V1/V1/A3/M2/M2/_0_  (.A1(\V3/V1/V1/A3/M2/s1 ),
    .A2(\V3/V1/V1/A3/c1 ),
    .ZN(\V3/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M2/M2/_1_  (.A(\V3/V1/V1/A3/M2/s1 ),
    .B(\V3/V1/V1/A3/c1 ),
    .Z(\V3/V1/v1 [5]));
 OR2_X1 \V3/V1/V1/A3/M2/_0_  (.A1(\V3/V1/V1/A3/M2/c1 ),
    .A2(\V3/V1/V1/A3/M2/c2 ),
    .ZN(\V3/V1/V1/A3/c2 ));
 AND2_X1 \V3/V1/V1/A3/M3/M1/_0_  (.A1(\V3/V1/V1/v4 [2]),
    .A2(\V3/V1/V1/c3 ),
    .ZN(\V3/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M3/M1/_1_  (.A(\V3/V1/V1/v4 [2]),
    .B(\V3/V1/V1/c3 ),
    .Z(\V3/V1/V1/A3/M3/s1 ));
 AND2_X1 \V3/V1/V1/A3/M3/M2/_0_  (.A1(\V3/V1/V1/A3/M3/s1 ),
    .A2(\V3/V1/V1/A3/c2 ),
    .ZN(\V3/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M3/M2/_1_  (.A(\V3/V1/V1/A3/M3/s1 ),
    .B(\V3/V1/V1/A3/c2 ),
    .Z(\V3/V1/v1 [6]));
 OR2_X1 \V3/V1/V1/A3/M3/_0_  (.A1(\V3/V1/V1/A3/M3/c1 ),
    .A2(\V3/V1/V1/A3/M3/c2 ),
    .ZN(\V3/V1/V1/A3/c3 ));
 AND2_X1 \V3/V1/V1/A3/M4/M1/_0_  (.A1(\V3/V1/V1/v4 [3]),
    .A2(net6),
    .ZN(\V3/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V1/A3/M4/M1/_1_  (.A(\V3/V1/V1/v4 [3]),
    .B(net6),
    .Z(\V3/V1/V1/A3/M4/s1 ));
 AND2_X1 \V3/V1/V1/A3/M4/M2/_0_  (.A1(\V3/V1/V1/A3/M4/s1 ),
    .A2(\V3/V1/V1/A3/c3 ),
    .ZN(\V3/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V1/A3/M4/M2/_1_  (.A(\V3/V1/V1/A3/M4/s1 ),
    .B(\V3/V1/V1/A3/c3 ),
    .Z(\V3/V1/v1 [7]));
 OR2_X1 \V3/V1/V1/A3/M4/_0_  (.A1(\V3/V1/V1/A3/M4/c1 ),
    .A2(\V3/V1/V1/A3/M4/c2 ),
    .ZN(\V3/V1/V1/overflow ));
 AND2_X1 \V3/V1/V1/V1/HA1/_0_  (.A1(\V3/V1/V1/V1/w2 ),
    .A2(\V3/V1/V1/V1/w1 ),
    .ZN(\V3/V1/V1/V1/w4 ));
 XOR2_X2 \V3/V1/V1/V1/HA1/_1_  (.A(\V3/V1/V1/V1/w2 ),
    .B(\V3/V1/V1/V1/w1 ),
    .Z(v3[1]));
 AND2_X1 \V3/V1/V1/V1/HA2/_0_  (.A1(\V3/V1/V1/V1/w4 ),
    .A2(\V3/V1/V1/V1/w3 ),
    .ZN(\V3/V1/V1/v1 [3]));
 XOR2_X2 \V3/V1/V1/V1/HA2/_1_  (.A(\V3/V1/V1/V1/w4 ),
    .B(\V3/V1/V1/V1/w3 ),
    .Z(\V3/V1/V1/v1 [2]));
 AND2_X1 \V3/V1/V1/V1/_0_  (.A1(net48),
    .A2(B[16]),
    .ZN(v3[0]));
 AND2_X1 \V3/V1/V1/V1/_1_  (.A1(net48),
    .A2(net21),
    .ZN(\V3/V1/V1/V1/w1 ));
 AND2_X1 \V3/V1/V1/V1/_2_  (.A1(net22),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V1/w2 ));
 AND2_X1 \V3/V1/V1/V1/_3_  (.A1(net21),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V1/w3 ));
 AND2_X1 \V3/V1/V1/V2/HA1/_0_  (.A1(\V3/V1/V1/V2/w2 ),
    .A2(\V3/V1/V1/V2/w1 ),
    .ZN(\V3/V1/V1/V2/w4 ));
 XOR2_X2 \V3/V1/V1/V2/HA1/_1_  (.A(\V3/V1/V1/V2/w2 ),
    .B(\V3/V1/V1/V2/w1 ),
    .Z(\V3/V1/V1/v2 [1]));
 AND2_X1 \V3/V1/V1/V2/HA2/_0_  (.A1(\V3/V1/V1/V2/w4 ),
    .A2(\V3/V1/V1/V2/w3 ),
    .ZN(\V3/V1/V1/v2 [3]));
 XOR2_X2 \V3/V1/V1/V2/HA2/_1_  (.A(\V3/V1/V1/V2/w4 ),
    .B(\V3/V1/V1/V2/w3 ),
    .Z(\V3/V1/V1/v2 [2]));
 AND2_X1 \V3/V1/V1/V2/_0_  (.A1(A[2]),
    .A2(net22),
    .ZN(\V3/V1/V1/v2 [0]));
 AND2_X1 \V3/V1/V1/V2/_1_  (.A1(A[2]),
    .A2(net21),
    .ZN(\V3/V1/V1/V2/w1 ));
 AND2_X1 \V3/V1/V1/V2/_2_  (.A1(net22),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V2/w2 ));
 AND2_X1 \V3/V1/V1/V2/_3_  (.A1(net21),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V2/w3 ));
 AND2_X1 \V3/V1/V1/V3/HA1/_0_  (.A1(\V3/V1/V1/V3/w2 ),
    .A2(\V3/V1/V1/V3/w1 ),
    .ZN(\V3/V1/V1/V3/w4 ));
 XOR2_X2 \V3/V1/V1/V3/HA1/_1_  (.A(\V3/V1/V1/V3/w2 ),
    .B(\V3/V1/V1/V3/w1 ),
    .Z(\V3/V1/V1/v3 [1]));
 AND2_X1 \V3/V1/V1/V3/HA2/_0_  (.A1(\V3/V1/V1/V3/w4 ),
    .A2(\V3/V1/V1/V3/w3 ),
    .ZN(\V3/V1/V1/v3 [3]));
 XOR2_X2 \V3/V1/V1/V3/HA2/_1_  (.A(\V3/V1/V1/V3/w4 ),
    .B(\V3/V1/V1/V3/w3 ),
    .Z(\V3/V1/V1/v3 [2]));
 AND2_X1 \V3/V1/V1/V3/_0_  (.A1(net48),
    .A2(net20),
    .ZN(\V3/V1/V1/v3 [0]));
 AND2_X1 \V3/V1/V1/V3/_1_  (.A1(net48),
    .A2(net19),
    .ZN(\V3/V1/V1/V3/w1 ));
 AND2_X1 \V3/V1/V1/V3/_2_  (.A1(net20),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V3/w2 ));
 AND2_X1 \V3/V1/V1/V3/_3_  (.A1(net19),
    .A2(A[1]),
    .ZN(\V3/V1/V1/V3/w3 ));
 AND2_X1 \V3/V1/V1/V4/HA1/_0_  (.A1(\V3/V1/V1/V4/w2 ),
    .A2(\V3/V1/V1/V4/w1 ),
    .ZN(\V3/V1/V1/V4/w4 ));
 XOR2_X2 \V3/V1/V1/V4/HA1/_1_  (.A(\V3/V1/V1/V4/w2 ),
    .B(\V3/V1/V1/V4/w1 ),
    .Z(\V3/V1/V1/v4 [1]));
 AND2_X1 \V3/V1/V1/V4/HA2/_0_  (.A1(\V3/V1/V1/V4/w4 ),
    .A2(\V3/V1/V1/V4/w3 ),
    .ZN(\V3/V1/V1/v4 [3]));
 XOR2_X2 \V3/V1/V1/V4/HA2/_1_  (.A(\V3/V1/V1/V4/w4 ),
    .B(\V3/V1/V1/V4/w3 ),
    .Z(\V3/V1/V1/v4 [2]));
 AND2_X1 \V3/V1/V1/V4/_0_  (.A1(A[2]),
    .A2(net20),
    .ZN(\V3/V1/V1/v4 [0]));
 AND2_X1 \V3/V1/V1/V4/_1_  (.A1(A[2]),
    .A2(net19),
    .ZN(\V3/V1/V1/V4/w1 ));
 AND2_X1 \V3/V1/V1/V4/_2_  (.A1(net20),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V4/w2 ));
 AND2_X1 \V3/V1/V1/V4/_3_  (.A1(net19),
    .A2(A[3]),
    .ZN(\V3/V1/V1/V4/w3 ));
 OR2_X1 \V3/V1/V1/_0_  (.A1(\V3/V1/V1/c1 ),
    .A2(\V3/V1/V1/c2 ),
    .ZN(\V3/V1/V1/c3 ));
 AND2_X1 \V3/V1/V2/A1/M1/M1/_0_  (.A1(\V3/V1/V2/v2 [0]),
    .A2(\V3/V1/V2/v3 [0]),
    .ZN(\V3/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M1/M1/_1_  (.A(\V3/V1/V2/v2 [0]),
    .B(\V3/V1/V2/v3 [0]),
    .Z(\V3/V1/V2/A1/M1/s1 ));
 AND2_X1 \V3/V1/V2/A1/M1/M2/_0_  (.A1(\V3/V1/V2/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M1/M2/_1_  (.A(\V3/V1/V2/A1/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/V2/s1 [0]));
 OR2_X1 \V3/V1/V2/A1/M1/_0_  (.A1(\V3/V1/V2/A1/M1/c1 ),
    .A2(\V3/V1/V2/A1/M1/c2 ),
    .ZN(\V3/V1/V2/A1/c1 ));
 AND2_X1 \V3/V1/V2/A1/M2/M1/_0_  (.A1(\V3/V1/V2/v2 [1]),
    .A2(\V3/V1/V2/v3 [1]),
    .ZN(\V3/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M2/M1/_1_  (.A(\V3/V1/V2/v2 [1]),
    .B(\V3/V1/V2/v3 [1]),
    .Z(\V3/V1/V2/A1/M2/s1 ));
 AND2_X1 \V3/V1/V2/A1/M2/M2/_0_  (.A1(\V3/V1/V2/A1/M2/s1 ),
    .A2(\V3/V1/V2/A1/c1 ),
    .ZN(\V3/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M2/M2/_1_  (.A(\V3/V1/V2/A1/M2/s1 ),
    .B(\V3/V1/V2/A1/c1 ),
    .Z(\V3/V1/V2/s1 [1]));
 OR2_X1 \V3/V1/V2/A1/M2/_0_  (.A1(\V3/V1/V2/A1/M2/c1 ),
    .A2(\V3/V1/V2/A1/M2/c2 ),
    .ZN(\V3/V1/V2/A1/c2 ));
 AND2_X1 \V3/V1/V2/A1/M3/M1/_0_  (.A1(\V3/V1/V2/v2 [2]),
    .A2(\V3/V1/V2/v3 [2]),
    .ZN(\V3/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M3/M1/_1_  (.A(\V3/V1/V2/v2 [2]),
    .B(\V3/V1/V2/v3 [2]),
    .Z(\V3/V1/V2/A1/M3/s1 ));
 AND2_X1 \V3/V1/V2/A1/M3/M2/_0_  (.A1(\V3/V1/V2/A1/M3/s1 ),
    .A2(\V3/V1/V2/A1/c2 ),
    .ZN(\V3/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M3/M2/_1_  (.A(\V3/V1/V2/A1/M3/s1 ),
    .B(\V3/V1/V2/A1/c2 ),
    .Z(\V3/V1/V2/s1 [2]));
 OR2_X1 \V3/V1/V2/A1/M3/_0_  (.A1(\V3/V1/V2/A1/M3/c1 ),
    .A2(\V3/V1/V2/A1/M3/c2 ),
    .ZN(\V3/V1/V2/A1/c3 ));
 AND2_X1 \V3/V1/V2/A1/M4/M1/_0_  (.A1(\V3/V1/V2/v2 [3]),
    .A2(\V3/V1/V2/v3 [3]),
    .ZN(\V3/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A1/M4/M1/_1_  (.A(\V3/V1/V2/v2 [3]),
    .B(\V3/V1/V2/v3 [3]),
    .Z(\V3/V1/V2/A1/M4/s1 ));
 AND2_X1 \V3/V1/V2/A1/M4/M2/_0_  (.A1(\V3/V1/V2/A1/M4/s1 ),
    .A2(\V3/V1/V2/A1/c3 ),
    .ZN(\V3/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A1/M4/M2/_1_  (.A(\V3/V1/V2/A1/M4/s1 ),
    .B(\V3/V1/V2/A1/c3 ),
    .Z(\V3/V1/V2/s1 [3]));
 OR2_X1 \V3/V1/V2/A1/M4/_0_  (.A1(\V3/V1/V2/A1/M4/c1 ),
    .A2(\V3/V1/V2/A1/M4/c2 ),
    .ZN(\V3/V1/V2/c1 ));
 AND2_X1 \V3/V1/V2/A2/M1/M1/_0_  (.A1(\V3/V1/V2/s1 [0]),
    .A2(\V3/V1/V2/v1 [2]),
    .ZN(\V3/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M1/M1/_1_  (.A(\V3/V1/V2/s1 [0]),
    .B(\V3/V1/V2/v1 [2]),
    .Z(\V3/V1/V2/A2/M1/s1 ));
 AND2_X1 \V3/V1/V2/A2/M1/M2/_0_  (.A1(\V3/V1/V2/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M1/M2/_1_  (.A(\V3/V1/V2/A2/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v2 [2]));
 OR2_X1 \V3/V1/V2/A2/M1/_0_  (.A1(\V3/V1/V2/A2/M1/c1 ),
    .A2(\V3/V1/V2/A2/M1/c2 ),
    .ZN(\V3/V1/V2/A2/c1 ));
 AND2_X1 \V3/V1/V2/A2/M2/M1/_0_  (.A1(\V3/V1/V2/s1 [1]),
    .A2(\V3/V1/V2/v1 [3]),
    .ZN(\V3/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M2/M1/_1_  (.A(\V3/V1/V2/s1 [1]),
    .B(\V3/V1/V2/v1 [3]),
    .Z(\V3/V1/V2/A2/M2/s1 ));
 AND2_X1 \V3/V1/V2/A2/M2/M2/_0_  (.A1(\V3/V1/V2/A2/M2/s1 ),
    .A2(\V3/V1/V2/A2/c1 ),
    .ZN(\V3/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M2/M2/_1_  (.A(\V3/V1/V2/A2/M2/s1 ),
    .B(\V3/V1/V2/A2/c1 ),
    .Z(\V3/V1/v2 [3]));
 OR2_X1 \V3/V1/V2/A2/M2/_0_  (.A1(\V3/V1/V2/A2/M2/c1 ),
    .A2(\V3/V1/V2/A2/M2/c2 ),
    .ZN(\V3/V1/V2/A2/c2 ));
 AND2_X1 \V3/V1/V2/A2/M3/M1/_0_  (.A1(\V3/V1/V2/s1 [2]),
    .A2(net2),
    .ZN(\V3/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M3/M1/_1_  (.A(\V3/V1/V2/s1 [2]),
    .B(net2),
    .Z(\V3/V1/V2/A2/M3/s1 ));
 AND2_X1 \V3/V1/V2/A2/M3/M2/_0_  (.A1(\V3/V1/V2/A2/M3/s1 ),
    .A2(\V3/V1/V2/A2/c2 ),
    .ZN(\V3/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M3/M2/_1_  (.A(\V3/V1/V2/A2/M3/s1 ),
    .B(\V3/V1/V2/A2/c2 ),
    .Z(\V3/V1/V2/s2 [2]));
 OR2_X1 \V3/V1/V2/A2/M3/_0_  (.A1(\V3/V1/V2/A2/M3/c1 ),
    .A2(\V3/V1/V2/A2/M3/c2 ),
    .ZN(\V3/V1/V2/A2/c3 ));
 AND2_X1 \V3/V1/V2/A2/M4/M1/_0_  (.A1(\V3/V1/V2/s1 [3]),
    .A2(net2),
    .ZN(\V3/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A2/M4/M1/_1_  (.A(\V3/V1/V2/s1 [3]),
    .B(net2),
    .Z(\V3/V1/V2/A2/M4/s1 ));
 AND2_X1 \V3/V1/V2/A2/M4/M2/_0_  (.A1(\V3/V1/V2/A2/M4/s1 ),
    .A2(\V3/V1/V2/A2/c3 ),
    .ZN(\V3/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A2/M4/M2/_1_  (.A(\V3/V1/V2/A2/M4/s1 ),
    .B(\V3/V1/V2/A2/c3 ),
    .Z(\V3/V1/V2/s2 [3]));
 OR2_X1 \V3/V1/V2/A2/M4/_0_  (.A1(\V3/V1/V2/A2/M4/c1 ),
    .A2(\V3/V1/V2/A2/M4/c2 ),
    .ZN(\V3/V1/V2/c2 ));
 AND2_X1 \V3/V1/V2/A3/M1/M1/_0_  (.A1(\V3/V1/V2/v4 [0]),
    .A2(\V3/V1/V2/s2 [2]),
    .ZN(\V3/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M1/M1/_1_  (.A(\V3/V1/V2/v4 [0]),
    .B(\V3/V1/V2/s2 [2]),
    .Z(\V3/V1/V2/A3/M1/s1 ));
 AND2_X1 \V3/V1/V2/A3/M1/M2/_0_  (.A1(\V3/V1/V2/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M1/M2/_1_  (.A(\V3/V1/V2/A3/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v2 [4]));
 OR2_X1 \V3/V1/V2/A3/M1/_0_  (.A1(\V3/V1/V2/A3/M1/c1 ),
    .A2(\V3/V1/V2/A3/M1/c2 ),
    .ZN(\V3/V1/V2/A3/c1 ));
 AND2_X1 \V3/V1/V2/A3/M2/M1/_0_  (.A1(\V3/V1/V2/v4 [1]),
    .A2(\V3/V1/V2/s2 [3]),
    .ZN(\V3/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M2/M1/_1_  (.A(\V3/V1/V2/v4 [1]),
    .B(\V3/V1/V2/s2 [3]),
    .Z(\V3/V1/V2/A3/M2/s1 ));
 AND2_X1 \V3/V1/V2/A3/M2/M2/_0_  (.A1(\V3/V1/V2/A3/M2/s1 ),
    .A2(\V3/V1/V2/A3/c1 ),
    .ZN(\V3/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M2/M2/_1_  (.A(\V3/V1/V2/A3/M2/s1 ),
    .B(\V3/V1/V2/A3/c1 ),
    .Z(\V3/V1/v2 [5]));
 OR2_X1 \V3/V1/V2/A3/M2/_0_  (.A1(\V3/V1/V2/A3/M2/c1 ),
    .A2(\V3/V1/V2/A3/M2/c2 ),
    .ZN(\V3/V1/V2/A3/c2 ));
 AND2_X1 \V3/V1/V2/A3/M3/M1/_0_  (.A1(\V3/V1/V2/v4 [2]),
    .A2(\V3/V1/V2/c3 ),
    .ZN(\V3/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M3/M1/_1_  (.A(\V3/V1/V2/v4 [2]),
    .B(\V3/V1/V2/c3 ),
    .Z(\V3/V1/V2/A3/M3/s1 ));
 AND2_X1 \V3/V1/V2/A3/M3/M2/_0_  (.A1(\V3/V1/V2/A3/M3/s1 ),
    .A2(\V3/V1/V2/A3/c2 ),
    .ZN(\V3/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M3/M2/_1_  (.A(\V3/V1/V2/A3/M3/s1 ),
    .B(\V3/V1/V2/A3/c2 ),
    .Z(\V3/V1/v2 [6]));
 OR2_X1 \V3/V1/V2/A3/M3/_0_  (.A1(\V3/V1/V2/A3/M3/c1 ),
    .A2(\V3/V1/V2/A3/M3/c2 ),
    .ZN(\V3/V1/V2/A3/c3 ));
 AND2_X1 \V3/V1/V2/A3/M4/M1/_0_  (.A1(\V3/V1/V2/v4 [3]),
    .A2(net2),
    .ZN(\V3/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V2/A3/M4/M1/_1_  (.A(\V3/V1/V2/v4 [3]),
    .B(net2),
    .Z(\V3/V1/V2/A3/M4/s1 ));
 AND2_X1 \V3/V1/V2/A3/M4/M2/_0_  (.A1(\V3/V1/V2/A3/M4/s1 ),
    .A2(\V3/V1/V2/A3/c3 ),
    .ZN(\V3/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V2/A3/M4/M2/_1_  (.A(\V3/V1/V2/A3/M4/s1 ),
    .B(\V3/V1/V2/A3/c3 ),
    .Z(\V3/V1/v2 [7]));
 OR2_X1 \V3/V1/V2/A3/M4/_0_  (.A1(\V3/V1/V2/A3/M4/c1 ),
    .A2(\V3/V1/V2/A3/M4/c2 ),
    .ZN(\V3/V1/V2/overflow ));
 AND2_X1 \V3/V1/V2/V1/HA1/_0_  (.A1(\V3/V1/V2/V1/w2 ),
    .A2(\V3/V1/V2/V1/w1 ),
    .ZN(\V3/V1/V2/V1/w4 ));
 XOR2_X2 \V3/V1/V2/V1/HA1/_1_  (.A(\V3/V1/V2/V1/w2 ),
    .B(\V3/V1/V2/V1/w1 ),
    .Z(\V3/V1/v2 [1]));
 AND2_X1 \V3/V1/V2/V1/HA2/_0_  (.A1(\V3/V1/V2/V1/w4 ),
    .A2(\V3/V1/V2/V1/w3 ),
    .ZN(\V3/V1/V2/v1 [3]));
 XOR2_X2 \V3/V1/V2/V1/HA2/_1_  (.A(\V3/V1/V2/V1/w4 ),
    .B(\V3/V1/V2/V1/w3 ),
    .Z(\V3/V1/V2/v1 [2]));
 AND2_X1 \V3/V1/V2/V1/_0_  (.A1(A[4]),
    .A2(net22),
    .ZN(\V3/V1/v2 [0]));
 AND2_X1 \V3/V1/V2/V1/_1_  (.A1(A[4]),
    .A2(net21),
    .ZN(\V3/V1/V2/V1/w1 ));
 AND2_X1 \V3/V1/V2/V1/_2_  (.A1(net22),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V1/w2 ));
 AND2_X1 \V3/V1/V2/V1/_3_  (.A1(net21),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V1/w3 ));
 AND2_X1 \V3/V1/V2/V2/HA1/_0_  (.A1(\V3/V1/V2/V2/w2 ),
    .A2(\V3/V1/V2/V2/w1 ),
    .ZN(\V3/V1/V2/V2/w4 ));
 XOR2_X2 \V3/V1/V2/V2/HA1/_1_  (.A(\V3/V1/V2/V2/w2 ),
    .B(\V3/V1/V2/V2/w1 ),
    .Z(\V3/V1/V2/v2 [1]));
 AND2_X1 \V3/V1/V2/V2/HA2/_0_  (.A1(\V3/V1/V2/V2/w4 ),
    .A2(\V3/V1/V2/V2/w3 ),
    .ZN(\V3/V1/V2/v2 [3]));
 XOR2_X2 \V3/V1/V2/V2/HA2/_1_  (.A(\V3/V1/V2/V2/w4 ),
    .B(\V3/V1/V2/V2/w3 ),
    .Z(\V3/V1/V2/v2 [2]));
 AND2_X1 \V3/V1/V2/V2/_0_  (.A1(A[6]),
    .A2(net22),
    .ZN(\V3/V1/V2/v2 [0]));
 AND2_X1 \V3/V1/V2/V2/_1_  (.A1(A[6]),
    .A2(net21),
    .ZN(\V3/V1/V2/V2/w1 ));
 AND2_X1 \V3/V1/V2/V2/_2_  (.A1(net22),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V2/w2 ));
 AND2_X1 \V3/V1/V2/V2/_3_  (.A1(net21),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V2/w3 ));
 AND2_X1 \V3/V1/V2/V3/HA1/_0_  (.A1(\V3/V1/V2/V3/w2 ),
    .A2(\V3/V1/V2/V3/w1 ),
    .ZN(\V3/V1/V2/V3/w4 ));
 XOR2_X2 \V3/V1/V2/V3/HA1/_1_  (.A(\V3/V1/V2/V3/w2 ),
    .B(\V3/V1/V2/V3/w1 ),
    .Z(\V3/V1/V2/v3 [1]));
 AND2_X1 \V3/V1/V2/V3/HA2/_0_  (.A1(\V3/V1/V2/V3/w4 ),
    .A2(\V3/V1/V2/V3/w3 ),
    .ZN(\V3/V1/V2/v3 [3]));
 XOR2_X2 \V3/V1/V2/V3/HA2/_1_  (.A(\V3/V1/V2/V3/w4 ),
    .B(\V3/V1/V2/V3/w3 ),
    .Z(\V3/V1/V2/v3 [2]));
 AND2_X1 \V3/V1/V2/V3/_0_  (.A1(A[4]),
    .A2(net20),
    .ZN(\V3/V1/V2/v3 [0]));
 AND2_X1 \V3/V1/V2/V3/_1_  (.A1(A[4]),
    .A2(net19),
    .ZN(\V3/V1/V2/V3/w1 ));
 AND2_X1 \V3/V1/V2/V3/_2_  (.A1(net20),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V3/w2 ));
 AND2_X1 \V3/V1/V2/V3/_3_  (.A1(net19),
    .A2(A[5]),
    .ZN(\V3/V1/V2/V3/w3 ));
 AND2_X1 \V3/V1/V2/V4/HA1/_0_  (.A1(\V3/V1/V2/V4/w2 ),
    .A2(\V3/V1/V2/V4/w1 ),
    .ZN(\V3/V1/V2/V4/w4 ));
 XOR2_X2 \V3/V1/V2/V4/HA1/_1_  (.A(\V3/V1/V2/V4/w2 ),
    .B(\V3/V1/V2/V4/w1 ),
    .Z(\V3/V1/V2/v4 [1]));
 AND2_X1 \V3/V1/V2/V4/HA2/_0_  (.A1(\V3/V1/V2/V4/w4 ),
    .A2(\V3/V1/V2/V4/w3 ),
    .ZN(\V3/V1/V2/v4 [3]));
 XOR2_X2 \V3/V1/V2/V4/HA2/_1_  (.A(\V3/V1/V2/V4/w4 ),
    .B(\V3/V1/V2/V4/w3 ),
    .Z(\V3/V1/V2/v4 [2]));
 AND2_X1 \V3/V1/V2/V4/_0_  (.A1(A[6]),
    .A2(net20),
    .ZN(\V3/V1/V2/v4 [0]));
 AND2_X1 \V3/V1/V2/V4/_1_  (.A1(A[6]),
    .A2(net19),
    .ZN(\V3/V1/V2/V4/w1 ));
 AND2_X1 \V3/V1/V2/V4/_2_  (.A1(net20),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V4/w2 ));
 AND2_X1 \V3/V1/V2/V4/_3_  (.A1(net19),
    .A2(A[7]),
    .ZN(\V3/V1/V2/V4/w3 ));
 OR2_X1 \V3/V1/V2/_0_  (.A1(\V3/V1/V2/c1 ),
    .A2(\V3/V1/V2/c2 ),
    .ZN(\V3/V1/V2/c3 ));
 AND2_X1 \V3/V1/V3/A1/M1/M1/_0_  (.A1(\V3/V1/V3/v2 [0]),
    .A2(\V3/V1/V3/v3 [0]),
    .ZN(\V3/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M1/M1/_1_  (.A(\V3/V1/V3/v2 [0]),
    .B(\V3/V1/V3/v3 [0]),
    .Z(\V3/V1/V3/A1/M1/s1 ));
 AND2_X1 \V3/V1/V3/A1/M1/M2/_0_  (.A1(\V3/V1/V3/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M1/M2/_1_  (.A(\V3/V1/V3/A1/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/V3/s1 [0]));
 OR2_X1 \V3/V1/V3/A1/M1/_0_  (.A1(\V3/V1/V3/A1/M1/c1 ),
    .A2(\V3/V1/V3/A1/M1/c2 ),
    .ZN(\V3/V1/V3/A1/c1 ));
 AND2_X1 \V3/V1/V3/A1/M2/M1/_0_  (.A1(\V3/V1/V3/v2 [1]),
    .A2(\V3/V1/V3/v3 [1]),
    .ZN(\V3/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M2/M1/_1_  (.A(\V3/V1/V3/v2 [1]),
    .B(\V3/V1/V3/v3 [1]),
    .Z(\V3/V1/V3/A1/M2/s1 ));
 AND2_X1 \V3/V1/V3/A1/M2/M2/_0_  (.A1(\V3/V1/V3/A1/M2/s1 ),
    .A2(\V3/V1/V3/A1/c1 ),
    .ZN(\V3/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M2/M2/_1_  (.A(\V3/V1/V3/A1/M2/s1 ),
    .B(\V3/V1/V3/A1/c1 ),
    .Z(\V3/V1/V3/s1 [1]));
 OR2_X1 \V3/V1/V3/A1/M2/_0_  (.A1(\V3/V1/V3/A1/M2/c1 ),
    .A2(\V3/V1/V3/A1/M2/c2 ),
    .ZN(\V3/V1/V3/A1/c2 ));
 AND2_X1 \V3/V1/V3/A1/M3/M1/_0_  (.A1(\V3/V1/V3/v2 [2]),
    .A2(\V3/V1/V3/v3 [2]),
    .ZN(\V3/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M3/M1/_1_  (.A(\V3/V1/V3/v2 [2]),
    .B(\V3/V1/V3/v3 [2]),
    .Z(\V3/V1/V3/A1/M3/s1 ));
 AND2_X1 \V3/V1/V3/A1/M3/M2/_0_  (.A1(\V3/V1/V3/A1/M3/s1 ),
    .A2(\V3/V1/V3/A1/c2 ),
    .ZN(\V3/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M3/M2/_1_  (.A(\V3/V1/V3/A1/M3/s1 ),
    .B(\V3/V1/V3/A1/c2 ),
    .Z(\V3/V1/V3/s1 [2]));
 OR2_X1 \V3/V1/V3/A1/M3/_0_  (.A1(\V3/V1/V3/A1/M3/c1 ),
    .A2(\V3/V1/V3/A1/M3/c2 ),
    .ZN(\V3/V1/V3/A1/c3 ));
 AND2_X1 \V3/V1/V3/A1/M4/M1/_0_  (.A1(\V3/V1/V3/v2 [3]),
    .A2(\V3/V1/V3/v3 [3]),
    .ZN(\V3/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A1/M4/M1/_1_  (.A(\V3/V1/V3/v2 [3]),
    .B(\V3/V1/V3/v3 [3]),
    .Z(\V3/V1/V3/A1/M4/s1 ));
 AND2_X1 \V3/V1/V3/A1/M4/M2/_0_  (.A1(\V3/V1/V3/A1/M4/s1 ),
    .A2(\V3/V1/V3/A1/c3 ),
    .ZN(\V3/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A1/M4/M2/_1_  (.A(\V3/V1/V3/A1/M4/s1 ),
    .B(\V3/V1/V3/A1/c3 ),
    .Z(\V3/V1/V3/s1 [3]));
 OR2_X1 \V3/V1/V3/A1/M4/_0_  (.A1(\V3/V1/V3/A1/M4/c1 ),
    .A2(\V3/V1/V3/A1/M4/c2 ),
    .ZN(\V3/V1/V3/c1 ));
 AND2_X1 \V3/V1/V3/A2/M1/M1/_0_  (.A1(\V3/V1/V3/s1 [0]),
    .A2(\V3/V1/V3/v1 [2]),
    .ZN(\V3/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M1/M1/_1_  (.A(\V3/V1/V3/s1 [0]),
    .B(\V3/V1/V3/v1 [2]),
    .Z(\V3/V1/V3/A2/M1/s1 ));
 AND2_X1 \V3/V1/V3/A2/M1/M2/_0_  (.A1(\V3/V1/V3/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M1/M2/_1_  (.A(\V3/V1/V3/A2/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v3 [2]));
 OR2_X1 \V3/V1/V3/A2/M1/_0_  (.A1(\V3/V1/V3/A2/M1/c1 ),
    .A2(\V3/V1/V3/A2/M1/c2 ),
    .ZN(\V3/V1/V3/A2/c1 ));
 AND2_X1 \V3/V1/V3/A2/M2/M1/_0_  (.A1(\V3/V1/V3/s1 [1]),
    .A2(\V3/V1/V3/v1 [3]),
    .ZN(\V3/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M2/M1/_1_  (.A(\V3/V1/V3/s1 [1]),
    .B(\V3/V1/V3/v1 [3]),
    .Z(\V3/V1/V3/A2/M2/s1 ));
 AND2_X1 \V3/V1/V3/A2/M2/M2/_0_  (.A1(\V3/V1/V3/A2/M2/s1 ),
    .A2(\V3/V1/V3/A2/c1 ),
    .ZN(\V3/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M2/M2/_1_  (.A(\V3/V1/V3/A2/M2/s1 ),
    .B(\V3/V1/V3/A2/c1 ),
    .Z(\V3/V1/v3 [3]));
 OR2_X1 \V3/V1/V3/A2/M2/_0_  (.A1(\V3/V1/V3/A2/M2/c1 ),
    .A2(\V3/V1/V3/A2/M2/c2 ),
    .ZN(\V3/V1/V3/A2/c2 ));
 AND2_X1 \V3/V1/V3/A2/M3/M1/_0_  (.A1(\V3/V1/V3/s1 [2]),
    .A2(net2),
    .ZN(\V3/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M3/M1/_1_  (.A(\V3/V1/V3/s1 [2]),
    .B(net2),
    .Z(\V3/V1/V3/A2/M3/s1 ));
 AND2_X1 \V3/V1/V3/A2/M3/M2/_0_  (.A1(\V3/V1/V3/A2/M3/s1 ),
    .A2(\V3/V1/V3/A2/c2 ),
    .ZN(\V3/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M3/M2/_1_  (.A(\V3/V1/V3/A2/M3/s1 ),
    .B(\V3/V1/V3/A2/c2 ),
    .Z(\V3/V1/V3/s2 [2]));
 OR2_X1 \V3/V1/V3/A2/M3/_0_  (.A1(\V3/V1/V3/A2/M3/c1 ),
    .A2(\V3/V1/V3/A2/M3/c2 ),
    .ZN(\V3/V1/V3/A2/c3 ));
 AND2_X1 \V3/V1/V3/A2/M4/M1/_0_  (.A1(\V3/V1/V3/s1 [3]),
    .A2(net2),
    .ZN(\V3/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A2/M4/M1/_1_  (.A(\V3/V1/V3/s1 [3]),
    .B(net2),
    .Z(\V3/V1/V3/A2/M4/s1 ));
 AND2_X1 \V3/V1/V3/A2/M4/M2/_0_  (.A1(\V3/V1/V3/A2/M4/s1 ),
    .A2(\V3/V1/V3/A2/c3 ),
    .ZN(\V3/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A2/M4/M2/_1_  (.A(\V3/V1/V3/A2/M4/s1 ),
    .B(\V3/V1/V3/A2/c3 ),
    .Z(\V3/V1/V3/s2 [3]));
 OR2_X1 \V3/V1/V3/A2/M4/_0_  (.A1(\V3/V1/V3/A2/M4/c1 ),
    .A2(\V3/V1/V3/A2/M4/c2 ),
    .ZN(\V3/V1/V3/c2 ));
 AND2_X1 \V3/V1/V3/A3/M1/M1/_0_  (.A1(\V3/V1/V3/v4 [0]),
    .A2(\V3/V1/V3/s2 [2]),
    .ZN(\V3/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M1/M1/_1_  (.A(\V3/V1/V3/v4 [0]),
    .B(\V3/V1/V3/s2 [2]),
    .Z(\V3/V1/V3/A3/M1/s1 ));
 AND2_X1 \V3/V1/V3/A3/M1/M2/_0_  (.A1(\V3/V1/V3/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M1/M2/_1_  (.A(\V3/V1/V3/A3/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v3 [4]));
 OR2_X1 \V3/V1/V3/A3/M1/_0_  (.A1(\V3/V1/V3/A3/M1/c1 ),
    .A2(\V3/V1/V3/A3/M1/c2 ),
    .ZN(\V3/V1/V3/A3/c1 ));
 AND2_X1 \V3/V1/V3/A3/M2/M1/_0_  (.A1(\V3/V1/V3/v4 [1]),
    .A2(\V3/V1/V3/s2 [3]),
    .ZN(\V3/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M2/M1/_1_  (.A(\V3/V1/V3/v4 [1]),
    .B(\V3/V1/V3/s2 [3]),
    .Z(\V3/V1/V3/A3/M2/s1 ));
 AND2_X1 \V3/V1/V3/A3/M2/M2/_0_  (.A1(\V3/V1/V3/A3/M2/s1 ),
    .A2(\V3/V1/V3/A3/c1 ),
    .ZN(\V3/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M2/M2/_1_  (.A(\V3/V1/V3/A3/M2/s1 ),
    .B(\V3/V1/V3/A3/c1 ),
    .Z(\V3/V1/v3 [5]));
 OR2_X1 \V3/V1/V3/A3/M2/_0_  (.A1(\V3/V1/V3/A3/M2/c1 ),
    .A2(\V3/V1/V3/A3/M2/c2 ),
    .ZN(\V3/V1/V3/A3/c2 ));
 AND2_X1 \V3/V1/V3/A3/M3/M1/_0_  (.A1(\V3/V1/V3/v4 [2]),
    .A2(\V3/V1/V3/c3 ),
    .ZN(\V3/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M3/M1/_1_  (.A(\V3/V1/V3/v4 [2]),
    .B(\V3/V1/V3/c3 ),
    .Z(\V3/V1/V3/A3/M3/s1 ));
 AND2_X1 \V3/V1/V3/A3/M3/M2/_0_  (.A1(\V3/V1/V3/A3/M3/s1 ),
    .A2(\V3/V1/V3/A3/c2 ),
    .ZN(\V3/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M3/M2/_1_  (.A(\V3/V1/V3/A3/M3/s1 ),
    .B(\V3/V1/V3/A3/c2 ),
    .Z(\V3/V1/v3 [6]));
 OR2_X1 \V3/V1/V3/A3/M3/_0_  (.A1(\V3/V1/V3/A3/M3/c1 ),
    .A2(\V3/V1/V3/A3/M3/c2 ),
    .ZN(\V3/V1/V3/A3/c3 ));
 AND2_X1 \V3/V1/V3/A3/M4/M1/_0_  (.A1(\V3/V1/V3/v4 [3]),
    .A2(net2),
    .ZN(\V3/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V3/A3/M4/M1/_1_  (.A(\V3/V1/V3/v4 [3]),
    .B(net2),
    .Z(\V3/V1/V3/A3/M4/s1 ));
 AND2_X1 \V3/V1/V3/A3/M4/M2/_0_  (.A1(\V3/V1/V3/A3/M4/s1 ),
    .A2(\V3/V1/V3/A3/c3 ),
    .ZN(\V3/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V3/A3/M4/M2/_1_  (.A(\V3/V1/V3/A3/M4/s1 ),
    .B(\V3/V1/V3/A3/c3 ),
    .Z(\V3/V1/v3 [7]));
 OR2_X1 \V3/V1/V3/A3/M4/_0_  (.A1(\V3/V1/V3/A3/M4/c1 ),
    .A2(\V3/V1/V3/A3/M4/c2 ),
    .ZN(\V3/V1/V3/overflow ));
 AND2_X1 \V3/V1/V3/V1/HA1/_0_  (.A1(\V3/V1/V3/V1/w2 ),
    .A2(\V3/V1/V3/V1/w1 ),
    .ZN(\V3/V1/V3/V1/w4 ));
 XOR2_X2 \V3/V1/V3/V1/HA1/_1_  (.A(\V3/V1/V3/V1/w2 ),
    .B(\V3/V1/V3/V1/w1 ),
    .Z(\V3/V1/v3 [1]));
 AND2_X1 \V3/V1/V3/V1/HA2/_0_  (.A1(\V3/V1/V3/V1/w4 ),
    .A2(\V3/V1/V3/V1/w3 ),
    .ZN(\V3/V1/V3/v1 [3]));
 XOR2_X2 \V3/V1/V3/V1/HA2/_1_  (.A(\V3/V1/V3/V1/w4 ),
    .B(\V3/V1/V3/V1/w3 ),
    .Z(\V3/V1/V3/v1 [2]));
 AND2_X1 \V3/V1/V3/V1/_0_  (.A1(net48),
    .A2(net18),
    .ZN(\V3/V1/v3 [0]));
 AND2_X1 \V3/V1/V3/V1/_1_  (.A1(net48),
    .A2(net17),
    .ZN(\V3/V1/V3/V1/w1 ));
 AND2_X1 \V3/V1/V3/V1/_2_  (.A1(net18),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V1/w2 ));
 AND2_X1 \V3/V1/V3/V1/_3_  (.A1(net17),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V1/w3 ));
 AND2_X1 \V3/V1/V3/V2/HA1/_0_  (.A1(\V3/V1/V3/V2/w2 ),
    .A2(\V3/V1/V3/V2/w1 ),
    .ZN(\V3/V1/V3/V2/w4 ));
 XOR2_X2 \V3/V1/V3/V2/HA1/_1_  (.A(\V3/V1/V3/V2/w2 ),
    .B(\V3/V1/V3/V2/w1 ),
    .Z(\V3/V1/V3/v2 [1]));
 AND2_X1 \V3/V1/V3/V2/HA2/_0_  (.A1(\V3/V1/V3/V2/w4 ),
    .A2(\V3/V1/V3/V2/w3 ),
    .ZN(\V3/V1/V3/v2 [3]));
 XOR2_X2 \V3/V1/V3/V2/HA2/_1_  (.A(\V3/V1/V3/V2/w4 ),
    .B(\V3/V1/V3/V2/w3 ),
    .Z(\V3/V1/V3/v2 [2]));
 AND2_X1 \V3/V1/V3/V2/_0_  (.A1(A[2]),
    .A2(net18),
    .ZN(\V3/V1/V3/v2 [0]));
 AND2_X1 \V3/V1/V3/V2/_1_  (.A1(A[2]),
    .A2(net17),
    .ZN(\V3/V1/V3/V2/w1 ));
 AND2_X1 \V3/V1/V3/V2/_2_  (.A1(net18),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V2/w2 ));
 AND2_X1 \V3/V1/V3/V2/_3_  (.A1(net17),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V2/w3 ));
 AND2_X1 \V3/V1/V3/V3/HA1/_0_  (.A1(\V3/V1/V3/V3/w2 ),
    .A2(\V3/V1/V3/V3/w1 ),
    .ZN(\V3/V1/V3/V3/w4 ));
 XOR2_X2 \V3/V1/V3/V3/HA1/_1_  (.A(\V3/V1/V3/V3/w2 ),
    .B(\V3/V1/V3/V3/w1 ),
    .Z(\V3/V1/V3/v3 [1]));
 AND2_X1 \V3/V1/V3/V3/HA2/_0_  (.A1(\V3/V1/V3/V3/w4 ),
    .A2(\V3/V1/V3/V3/w3 ),
    .ZN(\V3/V1/V3/v3 [3]));
 XOR2_X2 \V3/V1/V3/V3/HA2/_1_  (.A(\V3/V1/V3/V3/w4 ),
    .B(\V3/V1/V3/V3/w3 ),
    .Z(\V3/V1/V3/v3 [2]));
 AND2_X1 \V3/V1/V3/V3/_0_  (.A1(net48),
    .A2(B[22]),
    .ZN(\V3/V1/V3/v3 [0]));
 AND2_X1 \V3/V1/V3/V3/_1_  (.A1(net48),
    .A2(B[23]),
    .ZN(\V3/V1/V3/V3/w1 ));
 AND2_X1 \V3/V1/V3/V3/_2_  (.A1(B[22]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V3/w2 ));
 AND2_X1 \V3/V1/V3/V3/_3_  (.A1(B[23]),
    .A2(A[1]),
    .ZN(\V3/V1/V3/V3/w3 ));
 AND2_X1 \V3/V1/V3/V4/HA1/_0_  (.A1(\V3/V1/V3/V4/w2 ),
    .A2(\V3/V1/V3/V4/w1 ),
    .ZN(\V3/V1/V3/V4/w4 ));
 XOR2_X2 \V3/V1/V3/V4/HA1/_1_  (.A(\V3/V1/V3/V4/w2 ),
    .B(\V3/V1/V3/V4/w1 ),
    .Z(\V3/V1/V3/v4 [1]));
 AND2_X1 \V3/V1/V3/V4/HA2/_0_  (.A1(\V3/V1/V3/V4/w4 ),
    .A2(\V3/V1/V3/V4/w3 ),
    .ZN(\V3/V1/V3/v4 [3]));
 XOR2_X2 \V3/V1/V3/V4/HA2/_1_  (.A(\V3/V1/V3/V4/w4 ),
    .B(\V3/V1/V3/V4/w3 ),
    .Z(\V3/V1/V3/v4 [2]));
 AND2_X1 \V3/V1/V3/V4/_0_  (.A1(A[2]),
    .A2(B[22]),
    .ZN(\V3/V1/V3/v4 [0]));
 AND2_X1 \V3/V1/V3/V4/_1_  (.A1(A[2]),
    .A2(B[23]),
    .ZN(\V3/V1/V3/V4/w1 ));
 AND2_X1 \V3/V1/V3/V4/_2_  (.A1(B[22]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V4/w2 ));
 AND2_X1 \V3/V1/V3/V4/_3_  (.A1(B[23]),
    .A2(A[3]),
    .ZN(\V3/V1/V3/V4/w3 ));
 OR2_X1 \V3/V1/V3/_0_  (.A1(\V3/V1/V3/c1 ),
    .A2(\V3/V1/V3/c2 ),
    .ZN(\V3/V1/V3/c3 ));
 AND2_X1 \V3/V1/V4/A1/M1/M1/_0_  (.A1(\V3/V1/V4/v2 [0]),
    .A2(\V3/V1/V4/v3 [0]),
    .ZN(\V3/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M1/M1/_1_  (.A(\V3/V1/V4/v2 [0]),
    .B(\V3/V1/V4/v3 [0]),
    .Z(\V3/V1/V4/A1/M1/s1 ));
 AND2_X1 \V3/V1/V4/A1/M1/M2/_0_  (.A1(\V3/V1/V4/A1/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M1/M2/_1_  (.A(\V3/V1/V4/A1/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/V4/s1 [0]));
 OR2_X1 \V3/V1/V4/A1/M1/_0_  (.A1(\V3/V1/V4/A1/M1/c1 ),
    .A2(\V3/V1/V4/A1/M1/c2 ),
    .ZN(\V3/V1/V4/A1/c1 ));
 AND2_X1 \V3/V1/V4/A1/M2/M1/_0_  (.A1(\V3/V1/V4/v2 [1]),
    .A2(\V3/V1/V4/v3 [1]),
    .ZN(\V3/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M2/M1/_1_  (.A(\V3/V1/V4/v2 [1]),
    .B(\V3/V1/V4/v3 [1]),
    .Z(\V3/V1/V4/A1/M2/s1 ));
 AND2_X1 \V3/V1/V4/A1/M2/M2/_0_  (.A1(\V3/V1/V4/A1/M2/s1 ),
    .A2(\V3/V1/V4/A1/c1 ),
    .ZN(\V3/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M2/M2/_1_  (.A(\V3/V1/V4/A1/M2/s1 ),
    .B(\V3/V1/V4/A1/c1 ),
    .Z(\V3/V1/V4/s1 [1]));
 OR2_X1 \V3/V1/V4/A1/M2/_0_  (.A1(\V3/V1/V4/A1/M2/c1 ),
    .A2(\V3/V1/V4/A1/M2/c2 ),
    .ZN(\V3/V1/V4/A1/c2 ));
 AND2_X1 \V3/V1/V4/A1/M3/M1/_0_  (.A1(\V3/V1/V4/v2 [2]),
    .A2(\V3/V1/V4/v3 [2]),
    .ZN(\V3/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M3/M1/_1_  (.A(\V3/V1/V4/v2 [2]),
    .B(\V3/V1/V4/v3 [2]),
    .Z(\V3/V1/V4/A1/M3/s1 ));
 AND2_X1 \V3/V1/V4/A1/M3/M2/_0_  (.A1(\V3/V1/V4/A1/M3/s1 ),
    .A2(\V3/V1/V4/A1/c2 ),
    .ZN(\V3/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M3/M2/_1_  (.A(\V3/V1/V4/A1/M3/s1 ),
    .B(\V3/V1/V4/A1/c2 ),
    .Z(\V3/V1/V4/s1 [2]));
 OR2_X1 \V3/V1/V4/A1/M3/_0_  (.A1(\V3/V1/V4/A1/M3/c1 ),
    .A2(\V3/V1/V4/A1/M3/c2 ),
    .ZN(\V3/V1/V4/A1/c3 ));
 AND2_X1 \V3/V1/V4/A1/M4/M1/_0_  (.A1(\V3/V1/V4/v2 [3]),
    .A2(\V3/V1/V4/v3 [3]),
    .ZN(\V3/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A1/M4/M1/_1_  (.A(\V3/V1/V4/v2 [3]),
    .B(\V3/V1/V4/v3 [3]),
    .Z(\V3/V1/V4/A1/M4/s1 ));
 AND2_X1 \V3/V1/V4/A1/M4/M2/_0_  (.A1(\V3/V1/V4/A1/M4/s1 ),
    .A2(\V3/V1/V4/A1/c3 ),
    .ZN(\V3/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A1/M4/M2/_1_  (.A(\V3/V1/V4/A1/M4/s1 ),
    .B(\V3/V1/V4/A1/c3 ),
    .Z(\V3/V1/V4/s1 [3]));
 OR2_X1 \V3/V1/V4/A1/M4/_0_  (.A1(\V3/V1/V4/A1/M4/c1 ),
    .A2(\V3/V1/V4/A1/M4/c2 ),
    .ZN(\V3/V1/V4/c1 ));
 AND2_X1 \V3/V1/V4/A2/M1/M1/_0_  (.A1(\V3/V1/V4/s1 [0]),
    .A2(\V3/V1/V4/v1 [2]),
    .ZN(\V3/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M1/M1/_1_  (.A(\V3/V1/V4/s1 [0]),
    .B(\V3/V1/V4/v1 [2]),
    .Z(\V3/V1/V4/A2/M1/s1 ));
 AND2_X1 \V3/V1/V4/A2/M1/M2/_0_  (.A1(\V3/V1/V4/A2/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M1/M2/_1_  (.A(\V3/V1/V4/A2/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v4 [2]));
 OR2_X1 \V3/V1/V4/A2/M1/_0_  (.A1(\V3/V1/V4/A2/M1/c1 ),
    .A2(\V3/V1/V4/A2/M1/c2 ),
    .ZN(\V3/V1/V4/A2/c1 ));
 AND2_X1 \V3/V1/V4/A2/M2/M1/_0_  (.A1(\V3/V1/V4/s1 [1]),
    .A2(\V3/V1/V4/v1 [3]),
    .ZN(\V3/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M2/M1/_1_  (.A(\V3/V1/V4/s1 [1]),
    .B(\V3/V1/V4/v1 [3]),
    .Z(\V3/V1/V4/A2/M2/s1 ));
 AND2_X1 \V3/V1/V4/A2/M2/M2/_0_  (.A1(\V3/V1/V4/A2/M2/s1 ),
    .A2(\V3/V1/V4/A2/c1 ),
    .ZN(\V3/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M2/M2/_1_  (.A(\V3/V1/V4/A2/M2/s1 ),
    .B(\V3/V1/V4/A2/c1 ),
    .Z(\V3/V1/v4 [3]));
 OR2_X1 \V3/V1/V4/A2/M2/_0_  (.A1(\V3/V1/V4/A2/M2/c1 ),
    .A2(\V3/V1/V4/A2/M2/c2 ),
    .ZN(\V3/V1/V4/A2/c2 ));
 AND2_X1 \V3/V1/V4/A2/M3/M1/_0_  (.A1(\V3/V1/V4/s1 [2]),
    .A2(net2),
    .ZN(\V3/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M3/M1/_1_  (.A(\V3/V1/V4/s1 [2]),
    .B(net2),
    .Z(\V3/V1/V4/A2/M3/s1 ));
 AND2_X1 \V3/V1/V4/A2/M3/M2/_0_  (.A1(\V3/V1/V4/A2/M3/s1 ),
    .A2(\V3/V1/V4/A2/c2 ),
    .ZN(\V3/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M3/M2/_1_  (.A(\V3/V1/V4/A2/M3/s1 ),
    .B(\V3/V1/V4/A2/c2 ),
    .Z(\V3/V1/V4/s2 [2]));
 OR2_X1 \V3/V1/V4/A2/M3/_0_  (.A1(\V3/V1/V4/A2/M3/c1 ),
    .A2(\V3/V1/V4/A2/M3/c2 ),
    .ZN(\V3/V1/V4/A2/c3 ));
 AND2_X1 \V3/V1/V4/A2/M4/M1/_0_  (.A1(\V3/V1/V4/s1 [3]),
    .A2(net2),
    .ZN(\V3/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A2/M4/M1/_1_  (.A(\V3/V1/V4/s1 [3]),
    .B(net2),
    .Z(\V3/V1/V4/A2/M4/s1 ));
 AND2_X1 \V3/V1/V4/A2/M4/M2/_0_  (.A1(\V3/V1/V4/A2/M4/s1 ),
    .A2(\V3/V1/V4/A2/c3 ),
    .ZN(\V3/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A2/M4/M2/_1_  (.A(\V3/V1/V4/A2/M4/s1 ),
    .B(\V3/V1/V4/A2/c3 ),
    .Z(\V3/V1/V4/s2 [3]));
 OR2_X1 \V3/V1/V4/A2/M4/_0_  (.A1(\V3/V1/V4/A2/M4/c1 ),
    .A2(\V3/V1/V4/A2/M4/c2 ),
    .ZN(\V3/V1/V4/c2 ));
 AND2_X1 \V3/V1/V4/A3/M1/M1/_0_  (.A1(\V3/V1/V4/v4 [0]),
    .A2(\V3/V1/V4/s2 [2]),
    .ZN(\V3/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M1/M1/_1_  (.A(\V3/V1/V4/v4 [0]),
    .B(\V3/V1/V4/s2 [2]),
    .Z(\V3/V1/V4/A3/M1/s1 ));
 AND2_X1 \V3/V1/V4/A3/M1/M2/_0_  (.A1(\V3/V1/V4/A3/M1/s1 ),
    .A2(net2),
    .ZN(\V3/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M1/M2/_1_  (.A(\V3/V1/V4/A3/M1/s1 ),
    .B(net2),
    .Z(\V3/V1/v4 [4]));
 OR2_X1 \V3/V1/V4/A3/M1/_0_  (.A1(\V3/V1/V4/A3/M1/c1 ),
    .A2(\V3/V1/V4/A3/M1/c2 ),
    .ZN(\V3/V1/V4/A3/c1 ));
 AND2_X1 \V3/V1/V4/A3/M2/M1/_0_  (.A1(\V3/V1/V4/v4 [1]),
    .A2(\V3/V1/V4/s2 [3]),
    .ZN(\V3/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M2/M1/_1_  (.A(\V3/V1/V4/v4 [1]),
    .B(\V3/V1/V4/s2 [3]),
    .Z(\V3/V1/V4/A3/M2/s1 ));
 AND2_X1 \V3/V1/V4/A3/M2/M2/_0_  (.A1(\V3/V1/V4/A3/M2/s1 ),
    .A2(\V3/V1/V4/A3/c1 ),
    .ZN(\V3/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M2/M2/_1_  (.A(\V3/V1/V4/A3/M2/s1 ),
    .B(\V3/V1/V4/A3/c1 ),
    .Z(\V3/V1/v4 [5]));
 OR2_X1 \V3/V1/V4/A3/M2/_0_  (.A1(\V3/V1/V4/A3/M2/c1 ),
    .A2(\V3/V1/V4/A3/M2/c2 ),
    .ZN(\V3/V1/V4/A3/c2 ));
 AND2_X1 \V3/V1/V4/A3/M3/M1/_0_  (.A1(\V3/V1/V4/v4 [2]),
    .A2(\V3/V1/V4/c3 ),
    .ZN(\V3/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M3/M1/_1_  (.A(\V3/V1/V4/v4 [2]),
    .B(\V3/V1/V4/c3 ),
    .Z(\V3/V1/V4/A3/M3/s1 ));
 AND2_X1 \V3/V1/V4/A3/M3/M2/_0_  (.A1(\V3/V1/V4/A3/M3/s1 ),
    .A2(\V3/V1/V4/A3/c2 ),
    .ZN(\V3/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M3/M2/_1_  (.A(\V3/V1/V4/A3/M3/s1 ),
    .B(\V3/V1/V4/A3/c2 ),
    .Z(\V3/V1/v4 [6]));
 OR2_X1 \V3/V1/V4/A3/M3/_0_  (.A1(\V3/V1/V4/A3/M3/c1 ),
    .A2(\V3/V1/V4/A3/M3/c2 ),
    .ZN(\V3/V1/V4/A3/c3 ));
 AND2_X1 \V3/V1/V4/A3/M4/M1/_0_  (.A1(\V3/V1/V4/v4 [3]),
    .A2(net2),
    .ZN(\V3/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V1/V4/A3/M4/M1/_1_  (.A(\V3/V1/V4/v4 [3]),
    .B(net2),
    .Z(\V3/V1/V4/A3/M4/s1 ));
 AND2_X1 \V3/V1/V4/A3/M4/M2/_0_  (.A1(\V3/V1/V4/A3/M4/s1 ),
    .A2(\V3/V1/V4/A3/c3 ),
    .ZN(\V3/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V1/V4/A3/M4/M2/_1_  (.A(\V3/V1/V4/A3/M4/s1 ),
    .B(\V3/V1/V4/A3/c3 ),
    .Z(\V3/V1/v4 [7]));
 OR2_X1 \V3/V1/V4/A3/M4/_0_  (.A1(\V3/V1/V4/A3/M4/c1 ),
    .A2(\V3/V1/V4/A3/M4/c2 ),
    .ZN(\V3/V1/V4/overflow ));
 AND2_X1 \V3/V1/V4/V1/HA1/_0_  (.A1(\V3/V1/V4/V1/w2 ),
    .A2(\V3/V1/V4/V1/w1 ),
    .ZN(\V3/V1/V4/V1/w4 ));
 XOR2_X2 \V3/V1/V4/V1/HA1/_1_  (.A(\V3/V1/V4/V1/w2 ),
    .B(\V3/V1/V4/V1/w1 ),
    .Z(\V3/V1/v4 [1]));
 AND2_X1 \V3/V1/V4/V1/HA2/_0_  (.A1(\V3/V1/V4/V1/w4 ),
    .A2(\V3/V1/V4/V1/w3 ),
    .ZN(\V3/V1/V4/v1 [3]));
 XOR2_X2 \V3/V1/V4/V1/HA2/_1_  (.A(\V3/V1/V4/V1/w4 ),
    .B(\V3/V1/V4/V1/w3 ),
    .Z(\V3/V1/V4/v1 [2]));
 AND2_X1 \V3/V1/V4/V1/_0_  (.A1(A[4]),
    .A2(net18),
    .ZN(\V3/V1/v4 [0]));
 AND2_X1 \V3/V1/V4/V1/_1_  (.A1(A[4]),
    .A2(net17),
    .ZN(\V3/V1/V4/V1/w1 ));
 AND2_X1 \V3/V1/V4/V1/_2_  (.A1(net18),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V1/w2 ));
 AND2_X1 \V3/V1/V4/V1/_3_  (.A1(net17),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V1/w3 ));
 AND2_X1 \V3/V1/V4/V2/HA1/_0_  (.A1(\V3/V1/V4/V2/w2 ),
    .A2(\V3/V1/V4/V2/w1 ),
    .ZN(\V3/V1/V4/V2/w4 ));
 XOR2_X2 \V3/V1/V4/V2/HA1/_1_  (.A(\V3/V1/V4/V2/w2 ),
    .B(\V3/V1/V4/V2/w1 ),
    .Z(\V3/V1/V4/v2 [1]));
 AND2_X1 \V3/V1/V4/V2/HA2/_0_  (.A1(\V3/V1/V4/V2/w4 ),
    .A2(\V3/V1/V4/V2/w3 ),
    .ZN(\V3/V1/V4/v2 [3]));
 XOR2_X2 \V3/V1/V4/V2/HA2/_1_  (.A(\V3/V1/V4/V2/w4 ),
    .B(\V3/V1/V4/V2/w3 ),
    .Z(\V3/V1/V4/v2 [2]));
 AND2_X1 \V3/V1/V4/V2/_0_  (.A1(A[6]),
    .A2(net18),
    .ZN(\V3/V1/V4/v2 [0]));
 AND2_X1 \V3/V1/V4/V2/_1_  (.A1(A[6]),
    .A2(net17),
    .ZN(\V3/V1/V4/V2/w1 ));
 AND2_X1 \V3/V1/V4/V2/_2_  (.A1(net18),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V2/w2 ));
 AND2_X1 \V3/V1/V4/V2/_3_  (.A1(net17),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V2/w3 ));
 AND2_X1 \V3/V1/V4/V3/HA1/_0_  (.A1(\V3/V1/V4/V3/w2 ),
    .A2(\V3/V1/V4/V3/w1 ),
    .ZN(\V3/V1/V4/V3/w4 ));
 XOR2_X2 \V3/V1/V4/V3/HA1/_1_  (.A(\V3/V1/V4/V3/w2 ),
    .B(\V3/V1/V4/V3/w1 ),
    .Z(\V3/V1/V4/v3 [1]));
 AND2_X1 \V3/V1/V4/V3/HA2/_0_  (.A1(\V3/V1/V4/V3/w4 ),
    .A2(\V3/V1/V4/V3/w3 ),
    .ZN(\V3/V1/V4/v3 [3]));
 XOR2_X2 \V3/V1/V4/V3/HA2/_1_  (.A(\V3/V1/V4/V3/w4 ),
    .B(\V3/V1/V4/V3/w3 ),
    .Z(\V3/V1/V4/v3 [2]));
 AND2_X1 \V3/V1/V4/V3/_0_  (.A1(A[4]),
    .A2(B[22]),
    .ZN(\V3/V1/V4/v3 [0]));
 AND2_X1 \V3/V1/V4/V3/_1_  (.A1(A[4]),
    .A2(B[23]),
    .ZN(\V3/V1/V4/V3/w1 ));
 AND2_X1 \V3/V1/V4/V3/_2_  (.A1(B[22]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V3/w2 ));
 AND2_X1 \V3/V1/V4/V3/_3_  (.A1(B[23]),
    .A2(A[5]),
    .ZN(\V3/V1/V4/V3/w3 ));
 AND2_X1 \V3/V1/V4/V4/HA1/_0_  (.A1(\V3/V1/V4/V4/w2 ),
    .A2(\V3/V1/V4/V4/w1 ),
    .ZN(\V3/V1/V4/V4/w4 ));
 XOR2_X2 \V3/V1/V4/V4/HA1/_1_  (.A(\V3/V1/V4/V4/w2 ),
    .B(\V3/V1/V4/V4/w1 ),
    .Z(\V3/V1/V4/v4 [1]));
 AND2_X1 \V3/V1/V4/V4/HA2/_0_  (.A1(\V3/V1/V4/V4/w4 ),
    .A2(\V3/V1/V4/V4/w3 ),
    .ZN(\V3/V1/V4/v4 [3]));
 XOR2_X2 \V3/V1/V4/V4/HA2/_1_  (.A(\V3/V1/V4/V4/w4 ),
    .B(\V3/V1/V4/V4/w3 ),
    .Z(\V3/V1/V4/v4 [2]));
 AND2_X1 \V3/V1/V4/V4/_0_  (.A1(A[6]),
    .A2(B[22]),
    .ZN(\V3/V1/V4/v4 [0]));
 AND2_X1 \V3/V1/V4/V4/_1_  (.A1(A[6]),
    .A2(B[23]),
    .ZN(\V3/V1/V4/V4/w1 ));
 AND2_X1 \V3/V1/V4/V4/_2_  (.A1(B[22]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V4/w2 ));
 AND2_X1 \V3/V1/V4/V4/_3_  (.A1(B[23]),
    .A2(A[7]),
    .ZN(\V3/V1/V4/V4/w3 ));
 OR2_X1 \V3/V1/V4/_0_  (.A1(\V3/V1/V4/c1 ),
    .A2(\V3/V1/V4/c2 ),
    .ZN(\V3/V1/V4/c3 ));
 OR2_X1 \V3/V1/_0_  (.A1(\V3/V1/c1 ),
    .A2(\V3/V1/c2 ),
    .ZN(\V3/V1/c3 ));
 AND2_X1 \V3/V2/A1/A1/M1/M1/_0_  (.A1(\V3/V2/v2 [0]),
    .A2(\V3/V2/v3 [0]),
    .ZN(\V3/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M1/M1/_1_  (.A(\V3/V2/v2 [0]),
    .B(\V3/V2/v3 [0]),
    .Z(\V3/V2/A1/A1/M1/s1 ));
 AND2_X1 \V3/V2/A1/A1/M1/M2/_0_  (.A1(\V3/V2/A1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M1/M2/_1_  (.A(\V3/V2/A1/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/V2/s1 [0]));
 OR2_X1 \V3/V2/A1/A1/M1/_0_  (.A1(\V3/V2/A1/A1/M1/c1 ),
    .A2(\V3/V2/A1/A1/M1/c2 ),
    .ZN(\V3/V2/A1/A1/c1 ));
 AND2_X1 \V3/V2/A1/A1/M2/M1/_0_  (.A1(\V3/V2/v2 [1]),
    .A2(\V3/V2/v3 [1]),
    .ZN(\V3/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M2/M1/_1_  (.A(\V3/V2/v2 [1]),
    .B(\V3/V2/v3 [1]),
    .Z(\V3/V2/A1/A1/M2/s1 ));
 AND2_X1 \V3/V2/A1/A1/M2/M2/_0_  (.A1(\V3/V2/A1/A1/M2/s1 ),
    .A2(\V3/V2/A1/A1/c1 ),
    .ZN(\V3/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M2/M2/_1_  (.A(\V3/V2/A1/A1/M2/s1 ),
    .B(\V3/V2/A1/A1/c1 ),
    .Z(\V3/V2/s1 [1]));
 OR2_X1 \V3/V2/A1/A1/M2/_0_  (.A1(\V3/V2/A1/A1/M2/c1 ),
    .A2(\V3/V2/A1/A1/M2/c2 ),
    .ZN(\V3/V2/A1/A1/c2 ));
 AND2_X1 \V3/V2/A1/A1/M3/M1/_0_  (.A1(\V3/V2/v2 [2]),
    .A2(\V3/V2/v3 [2]),
    .ZN(\V3/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M3/M1/_1_  (.A(\V3/V2/v2 [2]),
    .B(\V3/V2/v3 [2]),
    .Z(\V3/V2/A1/A1/M3/s1 ));
 AND2_X1 \V3/V2/A1/A1/M3/M2/_0_  (.A1(\V3/V2/A1/A1/M3/s1 ),
    .A2(\V3/V2/A1/A1/c2 ),
    .ZN(\V3/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M3/M2/_1_  (.A(\V3/V2/A1/A1/M3/s1 ),
    .B(\V3/V2/A1/A1/c2 ),
    .Z(\V3/V2/s1 [2]));
 OR2_X1 \V3/V2/A1/A1/M3/_0_  (.A1(\V3/V2/A1/A1/M3/c1 ),
    .A2(\V3/V2/A1/A1/M3/c2 ),
    .ZN(\V3/V2/A1/A1/c3 ));
 AND2_X1 \V3/V2/A1/A1/M4/M1/_0_  (.A1(\V3/V2/v2 [3]),
    .A2(\V3/V2/v3 [3]),
    .ZN(\V3/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A1/A1/M4/M1/_1_  (.A(\V3/V2/v2 [3]),
    .B(\V3/V2/v3 [3]),
    .Z(\V3/V2/A1/A1/M4/s1 ));
 AND2_X1 \V3/V2/A1/A1/M4/M2/_0_  (.A1(\V3/V2/A1/A1/M4/s1 ),
    .A2(\V3/V2/A1/A1/c3 ),
    .ZN(\V3/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A1/A1/M4/M2/_1_  (.A(\V3/V2/A1/A1/M4/s1 ),
    .B(\V3/V2/A1/A1/c3 ),
    .Z(\V3/V2/s1 [3]));
 OR2_X1 \V3/V2/A1/A1/M4/_0_  (.A1(\V3/V2/A1/A1/M4/c1 ),
    .A2(\V3/V2/A1/A1/M4/c2 ),
    .ZN(\V3/V2/A1/c1 ));
 AND2_X1 \V3/V2/A1/A2/M1/M1/_0_  (.A1(\V3/V2/v2 [4]),
    .A2(\V3/V2/v3 [4]),
    .ZN(\V3/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M1/M1/_1_  (.A(\V3/V2/v2 [4]),
    .B(\V3/V2/v3 [4]),
    .Z(\V3/V2/A1/A2/M1/s1 ));
 AND2_X1 \V3/V2/A1/A2/M1/M2/_0_  (.A1(\V3/V2/A1/A2/M1/s1 ),
    .A2(\V3/V2/A1/c1 ),
    .ZN(\V3/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M1/M2/_1_  (.A(\V3/V2/A1/A2/M1/s1 ),
    .B(\V3/V2/A1/c1 ),
    .Z(\V3/V2/s1 [4]));
 OR2_X1 \V3/V2/A1/A2/M1/_0_  (.A1(\V3/V2/A1/A2/M1/c1 ),
    .A2(\V3/V2/A1/A2/M1/c2 ),
    .ZN(\V3/V2/A1/A2/c1 ));
 AND2_X1 \V3/V2/A1/A2/M2/M1/_0_  (.A1(\V3/V2/v2 [5]),
    .A2(\V3/V2/v3 [5]),
    .ZN(\V3/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M2/M1/_1_  (.A(\V3/V2/v2 [5]),
    .B(\V3/V2/v3 [5]),
    .Z(\V3/V2/A1/A2/M2/s1 ));
 AND2_X1 \V3/V2/A1/A2/M2/M2/_0_  (.A1(\V3/V2/A1/A2/M2/s1 ),
    .A2(\V3/V2/A1/A2/c1 ),
    .ZN(\V3/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M2/M2/_1_  (.A(\V3/V2/A1/A2/M2/s1 ),
    .B(\V3/V2/A1/A2/c1 ),
    .Z(\V3/V2/s1 [5]));
 OR2_X1 \V3/V2/A1/A2/M2/_0_  (.A1(\V3/V2/A1/A2/M2/c1 ),
    .A2(\V3/V2/A1/A2/M2/c2 ),
    .ZN(\V3/V2/A1/A2/c2 ));
 AND2_X1 \V3/V2/A1/A2/M3/M1/_0_  (.A1(\V3/V2/v2 [6]),
    .A2(\V3/V2/v3 [6]),
    .ZN(\V3/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M3/M1/_1_  (.A(\V3/V2/v2 [6]),
    .B(\V3/V2/v3 [6]),
    .Z(\V3/V2/A1/A2/M3/s1 ));
 AND2_X1 \V3/V2/A1/A2/M3/M2/_0_  (.A1(\V3/V2/A1/A2/M3/s1 ),
    .A2(\V3/V2/A1/A2/c2 ),
    .ZN(\V3/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M3/M2/_1_  (.A(\V3/V2/A1/A2/M3/s1 ),
    .B(\V3/V2/A1/A2/c2 ),
    .Z(\V3/V2/s1 [6]));
 OR2_X1 \V3/V2/A1/A2/M3/_0_  (.A1(\V3/V2/A1/A2/M3/c1 ),
    .A2(\V3/V2/A1/A2/M3/c2 ),
    .ZN(\V3/V2/A1/A2/c3 ));
 AND2_X1 \V3/V2/A1/A2/M4/M1/_0_  (.A1(\V3/V2/v2 [7]),
    .A2(\V3/V2/v3 [7]),
    .ZN(\V3/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A1/A2/M4/M1/_1_  (.A(\V3/V2/v2 [7]),
    .B(\V3/V2/v3 [7]),
    .Z(\V3/V2/A1/A2/M4/s1 ));
 AND2_X1 \V3/V2/A1/A2/M4/M2/_0_  (.A1(\V3/V2/A1/A2/M4/s1 ),
    .A2(\V3/V2/A1/A2/c3 ),
    .ZN(\V3/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A1/A2/M4/M2/_1_  (.A(\V3/V2/A1/A2/M4/s1 ),
    .B(\V3/V2/A1/A2/c3 ),
    .Z(\V3/V2/s1 [7]));
 OR2_X1 \V3/V2/A1/A2/M4/_0_  (.A1(\V3/V2/A1/A2/M4/c1 ),
    .A2(\V3/V2/A1/A2/M4/c2 ),
    .ZN(\V3/V2/c1 ));
 AND2_X1 \V3/V2/A2/A1/M1/M1/_0_  (.A1(\V3/V2/s1 [0]),
    .A2(\V3/V2/v1 [4]),
    .ZN(\V3/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M1/M1/_1_  (.A(\V3/V2/s1 [0]),
    .B(\V3/V2/v1 [4]),
    .Z(\V3/V2/A2/A1/M1/s1 ));
 AND2_X1 \V3/V2/A2/A1/M1/M2/_0_  (.A1(\V3/V2/A2/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M1/M2/_1_  (.A(\V3/V2/A2/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/v2 [4]));
 OR2_X1 \V3/V2/A2/A1/M1/_0_  (.A1(\V3/V2/A2/A1/M1/c1 ),
    .A2(\V3/V2/A2/A1/M1/c2 ),
    .ZN(\V3/V2/A2/A1/c1 ));
 AND2_X1 \V3/V2/A2/A1/M2/M1/_0_  (.A1(\V3/V2/s1 [1]),
    .A2(\V3/V2/v1 [5]),
    .ZN(\V3/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M2/M1/_1_  (.A(\V3/V2/s1 [1]),
    .B(\V3/V2/v1 [5]),
    .Z(\V3/V2/A2/A1/M2/s1 ));
 AND2_X1 \V3/V2/A2/A1/M2/M2/_0_  (.A1(\V3/V2/A2/A1/M2/s1 ),
    .A2(\V3/V2/A2/A1/c1 ),
    .ZN(\V3/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M2/M2/_1_  (.A(\V3/V2/A2/A1/M2/s1 ),
    .B(\V3/V2/A2/A1/c1 ),
    .Z(\V3/v2 [5]));
 OR2_X1 \V3/V2/A2/A1/M2/_0_  (.A1(\V3/V2/A2/A1/M2/c1 ),
    .A2(\V3/V2/A2/A1/M2/c2 ),
    .ZN(\V3/V2/A2/A1/c2 ));
 AND2_X1 \V3/V2/A2/A1/M3/M1/_0_  (.A1(\V3/V2/s1 [2]),
    .A2(\V3/V2/v1 [6]),
    .ZN(\V3/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M3/M1/_1_  (.A(\V3/V2/s1 [2]),
    .B(\V3/V2/v1 [6]),
    .Z(\V3/V2/A2/A1/M3/s1 ));
 AND2_X1 \V3/V2/A2/A1/M3/M2/_0_  (.A1(\V3/V2/A2/A1/M3/s1 ),
    .A2(\V3/V2/A2/A1/c2 ),
    .ZN(\V3/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M3/M2/_1_  (.A(\V3/V2/A2/A1/M3/s1 ),
    .B(\V3/V2/A2/A1/c2 ),
    .Z(\V3/v2 [6]));
 OR2_X1 \V3/V2/A2/A1/M3/_0_  (.A1(\V3/V2/A2/A1/M3/c1 ),
    .A2(\V3/V2/A2/A1/M3/c2 ),
    .ZN(\V3/V2/A2/A1/c3 ));
 AND2_X1 \V3/V2/A2/A1/M4/M1/_0_  (.A1(\V3/V2/s1 [3]),
    .A2(\V3/V2/v1 [7]),
    .ZN(\V3/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A2/A1/M4/M1/_1_  (.A(\V3/V2/s1 [3]),
    .B(\V3/V2/v1 [7]),
    .Z(\V3/V2/A2/A1/M4/s1 ));
 AND2_X1 \V3/V2/A2/A1/M4/M2/_0_  (.A1(\V3/V2/A2/A1/M4/s1 ),
    .A2(\V3/V2/A2/A1/c3 ),
    .ZN(\V3/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A2/A1/M4/M2/_1_  (.A(\V3/V2/A2/A1/M4/s1 ),
    .B(\V3/V2/A2/A1/c3 ),
    .Z(\V3/v2 [7]));
 OR2_X1 \V3/V2/A2/A1/M4/_0_  (.A1(\V3/V2/A2/A1/M4/c1 ),
    .A2(\V3/V2/A2/A1/M4/c2 ),
    .ZN(\V3/V2/A2/c1 ));
 AND2_X1 \V3/V2/A2/A2/M1/M1/_0_  (.A1(\V3/V2/s1 [4]),
    .A2(net5),
    .ZN(\V3/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M1/M1/_1_  (.A(\V3/V2/s1 [4]),
    .B(net5),
    .Z(\V3/V2/A2/A2/M1/s1 ));
 AND2_X1 \V3/V2/A2/A2/M1/M2/_0_  (.A1(\V3/V2/A2/A2/M1/s1 ),
    .A2(\V3/V2/A2/c1 ),
    .ZN(\V3/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M1/M2/_1_  (.A(\V3/V2/A2/A2/M1/s1 ),
    .B(\V3/V2/A2/c1 ),
    .Z(\V3/V2/s2 [4]));
 OR2_X1 \V3/V2/A2/A2/M1/_0_  (.A1(\V3/V2/A2/A2/M1/c1 ),
    .A2(\V3/V2/A2/A2/M1/c2 ),
    .ZN(\V3/V2/A2/A2/c1 ));
 AND2_X1 \V3/V2/A2/A2/M2/M1/_0_  (.A1(\V3/V2/s1 [5]),
    .A2(net5),
    .ZN(\V3/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M2/M1/_1_  (.A(\V3/V2/s1 [5]),
    .B(net5),
    .Z(\V3/V2/A2/A2/M2/s1 ));
 AND2_X1 \V3/V2/A2/A2/M2/M2/_0_  (.A1(\V3/V2/A2/A2/M2/s1 ),
    .A2(\V3/V2/A2/A2/c1 ),
    .ZN(\V3/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M2/M2/_1_  (.A(\V3/V2/A2/A2/M2/s1 ),
    .B(\V3/V2/A2/A2/c1 ),
    .Z(\V3/V2/s2 [5]));
 OR2_X1 \V3/V2/A2/A2/M2/_0_  (.A1(\V3/V2/A2/A2/M2/c1 ),
    .A2(\V3/V2/A2/A2/M2/c2 ),
    .ZN(\V3/V2/A2/A2/c2 ));
 AND2_X1 \V3/V2/A2/A2/M3/M1/_0_  (.A1(\V3/V2/s1 [6]),
    .A2(net5),
    .ZN(\V3/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M3/M1/_1_  (.A(\V3/V2/s1 [6]),
    .B(net5),
    .Z(\V3/V2/A2/A2/M3/s1 ));
 AND2_X1 \V3/V2/A2/A2/M3/M2/_0_  (.A1(\V3/V2/A2/A2/M3/s1 ),
    .A2(\V3/V2/A2/A2/c2 ),
    .ZN(\V3/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M3/M2/_1_  (.A(\V3/V2/A2/A2/M3/s1 ),
    .B(\V3/V2/A2/A2/c2 ),
    .Z(\V3/V2/s2 [6]));
 OR2_X1 \V3/V2/A2/A2/M3/_0_  (.A1(\V3/V2/A2/A2/M3/c1 ),
    .A2(\V3/V2/A2/A2/M3/c2 ),
    .ZN(\V3/V2/A2/A2/c3 ));
 AND2_X1 \V3/V2/A2/A2/M4/M1/_0_  (.A1(\V3/V2/s1 [7]),
    .A2(net5),
    .ZN(\V3/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A2/A2/M4/M1/_1_  (.A(\V3/V2/s1 [7]),
    .B(net5),
    .Z(\V3/V2/A2/A2/M4/s1 ));
 AND2_X1 \V3/V2/A2/A2/M4/M2/_0_  (.A1(\V3/V2/A2/A2/M4/s1 ),
    .A2(\V3/V2/A2/A2/c3 ),
    .ZN(\V3/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A2/A2/M4/M2/_1_  (.A(\V3/V2/A2/A2/M4/s1 ),
    .B(\V3/V2/A2/A2/c3 ),
    .Z(\V3/V2/s2 [7]));
 OR2_X1 \V3/V2/A2/A2/M4/_0_  (.A1(\V3/V2/A2/A2/M4/c1 ),
    .A2(\V3/V2/A2/A2/M4/c2 ),
    .ZN(\V3/V2/c2 ));
 AND2_X1 \V3/V2/A3/A1/M1/M1/_0_  (.A1(\V3/V2/v4 [0]),
    .A2(\V3/V2/s2 [4]),
    .ZN(\V3/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M1/M1/_1_  (.A(\V3/V2/v4 [0]),
    .B(\V3/V2/s2 [4]),
    .Z(\V3/V2/A3/A1/M1/s1 ));
 AND2_X1 \V3/V2/A3/A1/M1/M2/_0_  (.A1(\V3/V2/A3/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M1/M2/_1_  (.A(\V3/V2/A3/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/v2 [8]));
 OR2_X1 \V3/V2/A3/A1/M1/_0_  (.A1(\V3/V2/A3/A1/M1/c1 ),
    .A2(\V3/V2/A3/A1/M1/c2 ),
    .ZN(\V3/V2/A3/A1/c1 ));
 AND2_X1 \V3/V2/A3/A1/M2/M1/_0_  (.A1(\V3/V2/v4 [1]),
    .A2(\V3/V2/s2 [5]),
    .ZN(\V3/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M2/M1/_1_  (.A(\V3/V2/v4 [1]),
    .B(\V3/V2/s2 [5]),
    .Z(\V3/V2/A3/A1/M2/s1 ));
 AND2_X1 \V3/V2/A3/A1/M2/M2/_0_  (.A1(\V3/V2/A3/A1/M2/s1 ),
    .A2(\V3/V2/A3/A1/c1 ),
    .ZN(\V3/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M2/M2/_1_  (.A(\V3/V2/A3/A1/M2/s1 ),
    .B(\V3/V2/A3/A1/c1 ),
    .Z(\V3/v2 [9]));
 OR2_X1 \V3/V2/A3/A1/M2/_0_  (.A1(\V3/V2/A3/A1/M2/c1 ),
    .A2(\V3/V2/A3/A1/M2/c2 ),
    .ZN(\V3/V2/A3/A1/c2 ));
 AND2_X1 \V3/V2/A3/A1/M3/M1/_0_  (.A1(\V3/V2/v4 [2]),
    .A2(\V3/V2/s2 [6]),
    .ZN(\V3/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M3/M1/_1_  (.A(\V3/V2/v4 [2]),
    .B(\V3/V2/s2 [6]),
    .Z(\V3/V2/A3/A1/M3/s1 ));
 AND2_X1 \V3/V2/A3/A1/M3/M2/_0_  (.A1(\V3/V2/A3/A1/M3/s1 ),
    .A2(\V3/V2/A3/A1/c2 ),
    .ZN(\V3/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M3/M2/_1_  (.A(\V3/V2/A3/A1/M3/s1 ),
    .B(\V3/V2/A3/A1/c2 ),
    .Z(\V3/v2 [10]));
 OR2_X1 \V3/V2/A3/A1/M3/_0_  (.A1(\V3/V2/A3/A1/M3/c1 ),
    .A2(\V3/V2/A3/A1/M3/c2 ),
    .ZN(\V3/V2/A3/A1/c3 ));
 AND2_X1 \V3/V2/A3/A1/M4/M1/_0_  (.A1(\V3/V2/v4 [3]),
    .A2(\V3/V2/s2 [7]),
    .ZN(\V3/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V2/A3/A1/M4/M1/_1_  (.A(\V3/V2/v4 [3]),
    .B(\V3/V2/s2 [7]),
    .Z(\V3/V2/A3/A1/M4/s1 ));
 AND2_X1 \V3/V2/A3/A1/M4/M2/_0_  (.A1(\V3/V2/A3/A1/M4/s1 ),
    .A2(\V3/V2/A3/A1/c3 ),
    .ZN(\V3/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V2/A3/A1/M4/M2/_1_  (.A(\V3/V2/A3/A1/M4/s1 ),
    .B(\V3/V2/A3/A1/c3 ),
    .Z(\V3/v2 [11]));
 OR2_X1 \V3/V2/A3/A1/M4/_0_  (.A1(\V3/V2/A3/A1/M4/c1 ),
    .A2(\V3/V2/A3/A1/M4/c2 ),
    .ZN(\V3/V2/A3/c1 ));
 AND2_X1 \V3/V2/A3/A2/M1/M1/_0_  (.A1(\V3/V2/v4 [4]),
    .A2(\V3/V2/c3 ),
    .ZN(\V3/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M1/M1/_1_  (.A(\V3/V2/v4 [4]),
    .B(\V3/V2/c3 ),
    .Z(\V3/V2/A3/A2/M1/s1 ));
 AND2_X1 \V3/V2/A3/A2/M1/M2/_0_  (.A1(\V3/V2/A3/A2/M1/s1 ),
    .A2(\V3/V2/A3/c1 ),
    .ZN(\V3/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M1/M2/_1_  (.A(\V3/V2/A3/A2/M1/s1 ),
    .B(\V3/V2/A3/c1 ),
    .Z(\V3/v2 [12]));
 OR2_X1 \V3/V2/A3/A2/M1/_0_  (.A1(\V3/V2/A3/A2/M1/c1 ),
    .A2(\V3/V2/A3/A2/M1/c2 ),
    .ZN(\V3/V2/A3/A2/c1 ));
 AND2_X1 \V3/V2/A3/A2/M2/M1/_0_  (.A1(\V3/V2/v4 [5]),
    .A2(net8),
    .ZN(\V3/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M2/M1/_1_  (.A(\V3/V2/v4 [5]),
    .B(net8),
    .Z(\V3/V2/A3/A2/M2/s1 ));
 AND2_X1 \V3/V2/A3/A2/M2/M2/_0_  (.A1(\V3/V2/A3/A2/M2/s1 ),
    .A2(\V3/V2/A3/A2/c1 ),
    .ZN(\V3/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M2/M2/_1_  (.A(\V3/V2/A3/A2/M2/s1 ),
    .B(\V3/V2/A3/A2/c1 ),
    .Z(\V3/v2 [13]));
 OR2_X1 \V3/V2/A3/A2/M2/_0_  (.A1(\V3/V2/A3/A2/M2/c1 ),
    .A2(\V3/V2/A3/A2/M2/c2 ),
    .ZN(\V3/V2/A3/A2/c2 ));
 AND2_X1 \V3/V2/A3/A2/M3/M1/_0_  (.A1(\V3/V2/v4 [6]),
    .A2(net8),
    .ZN(\V3/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M3/M1/_1_  (.A(\V3/V2/v4 [6]),
    .B(net8),
    .Z(\V3/V2/A3/A2/M3/s1 ));
 AND2_X1 \V3/V2/A3/A2/M3/M2/_0_  (.A1(\V3/V2/A3/A2/M3/s1 ),
    .A2(\V3/V2/A3/A2/c2 ),
    .ZN(\V3/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M3/M2/_1_  (.A(\V3/V2/A3/A2/M3/s1 ),
    .B(\V3/V2/A3/A2/c2 ),
    .Z(\V3/v2 [14]));
 OR2_X1 \V3/V2/A3/A2/M3/_0_  (.A1(\V3/V2/A3/A2/M3/c1 ),
    .A2(\V3/V2/A3/A2/M3/c2 ),
    .ZN(\V3/V2/A3/A2/c3 ));
 AND2_X1 \V3/V2/A3/A2/M4/M1/_0_  (.A1(\V3/V2/v4 [7]),
    .A2(net8),
    .ZN(\V3/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V2/A3/A2/M4/M1/_1_  (.A(\V3/V2/v4 [7]),
    .B(net8),
    .Z(\V3/V2/A3/A2/M4/s1 ));
 AND2_X1 \V3/V2/A3/A2/M4/M2/_0_  (.A1(\V3/V2/A3/A2/M4/s1 ),
    .A2(\V3/V2/A3/A2/c3 ),
    .ZN(\V3/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V2/A3/A2/M4/M2/_1_  (.A(\V3/V2/A3/A2/M4/s1 ),
    .B(\V3/V2/A3/A2/c3 ),
    .Z(\V3/v2 [15]));
 OR2_X1 \V3/V2/A3/A2/M4/_0_  (.A1(\V3/V2/A3/A2/M4/c1 ),
    .A2(\V3/V2/A3/A2/M4/c2 ),
    .ZN(\V3/V2/overflow ));
 AND2_X1 \V3/V2/V1/A1/M1/M1/_0_  (.A1(\V3/V2/V1/v2 [0]),
    .A2(\V3/V2/V1/v3 [0]),
    .ZN(\V3/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M1/M1/_1_  (.A(\V3/V2/V1/v2 [0]),
    .B(\V3/V2/V1/v3 [0]),
    .Z(\V3/V2/V1/A1/M1/s1 ));
 AND2_X1 \V3/V2/V1/A1/M1/M2/_0_  (.A1(\V3/V2/V1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M1/M2/_1_  (.A(\V3/V2/V1/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/V1/s1 [0]));
 OR2_X1 \V3/V2/V1/A1/M1/_0_  (.A1(\V3/V2/V1/A1/M1/c1 ),
    .A2(\V3/V2/V1/A1/M1/c2 ),
    .ZN(\V3/V2/V1/A1/c1 ));
 AND2_X1 \V3/V2/V1/A1/M2/M1/_0_  (.A1(\V3/V2/V1/v2 [1]),
    .A2(\V3/V2/V1/v3 [1]),
    .ZN(\V3/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M2/M1/_1_  (.A(\V3/V2/V1/v2 [1]),
    .B(\V3/V2/V1/v3 [1]),
    .Z(\V3/V2/V1/A1/M2/s1 ));
 AND2_X1 \V3/V2/V1/A1/M2/M2/_0_  (.A1(\V3/V2/V1/A1/M2/s1 ),
    .A2(\V3/V2/V1/A1/c1 ),
    .ZN(\V3/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M2/M2/_1_  (.A(\V3/V2/V1/A1/M2/s1 ),
    .B(\V3/V2/V1/A1/c1 ),
    .Z(\V3/V2/V1/s1 [1]));
 OR2_X1 \V3/V2/V1/A1/M2/_0_  (.A1(\V3/V2/V1/A1/M2/c1 ),
    .A2(\V3/V2/V1/A1/M2/c2 ),
    .ZN(\V3/V2/V1/A1/c2 ));
 AND2_X1 \V3/V2/V1/A1/M3/M1/_0_  (.A1(\V3/V2/V1/v2 [2]),
    .A2(\V3/V2/V1/v3 [2]),
    .ZN(\V3/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M3/M1/_1_  (.A(\V3/V2/V1/v2 [2]),
    .B(\V3/V2/V1/v3 [2]),
    .Z(\V3/V2/V1/A1/M3/s1 ));
 AND2_X1 \V3/V2/V1/A1/M3/M2/_0_  (.A1(\V3/V2/V1/A1/M3/s1 ),
    .A2(\V3/V2/V1/A1/c2 ),
    .ZN(\V3/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M3/M2/_1_  (.A(\V3/V2/V1/A1/M3/s1 ),
    .B(\V3/V2/V1/A1/c2 ),
    .Z(\V3/V2/V1/s1 [2]));
 OR2_X1 \V3/V2/V1/A1/M3/_0_  (.A1(\V3/V2/V1/A1/M3/c1 ),
    .A2(\V3/V2/V1/A1/M3/c2 ),
    .ZN(\V3/V2/V1/A1/c3 ));
 AND2_X1 \V3/V2/V1/A1/M4/M1/_0_  (.A1(\V3/V2/V1/v2 [3]),
    .A2(\V3/V2/V1/v3 [3]),
    .ZN(\V3/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A1/M4/M1/_1_  (.A(\V3/V2/V1/v2 [3]),
    .B(\V3/V2/V1/v3 [3]),
    .Z(\V3/V2/V1/A1/M4/s1 ));
 AND2_X1 \V3/V2/V1/A1/M4/M2/_0_  (.A1(\V3/V2/V1/A1/M4/s1 ),
    .A2(\V3/V2/V1/A1/c3 ),
    .ZN(\V3/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A1/M4/M2/_1_  (.A(\V3/V2/V1/A1/M4/s1 ),
    .B(\V3/V2/V1/A1/c3 ),
    .Z(\V3/V2/V1/s1 [3]));
 OR2_X1 \V3/V2/V1/A1/M4/_0_  (.A1(\V3/V2/V1/A1/M4/c1 ),
    .A2(\V3/V2/V1/A1/M4/c2 ),
    .ZN(\V3/V2/V1/c1 ));
 AND2_X1 \V3/V2/V1/A2/M1/M1/_0_  (.A1(\V3/V2/V1/s1 [0]),
    .A2(\V3/V2/V1/v1 [2]),
    .ZN(\V3/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M1/M1/_1_  (.A(\V3/V2/V1/s1 [0]),
    .B(\V3/V2/V1/v1 [2]),
    .Z(\V3/V2/V1/A2/M1/s1 ));
 AND2_X1 \V3/V2/V1/A2/M1/M2/_0_  (.A1(\V3/V2/V1/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M1/M2/_1_  (.A(\V3/V2/V1/A2/M1/s1 ),
    .B(net5),
    .Z(\V3/v2 [2]));
 OR2_X1 \V3/V2/V1/A2/M1/_0_  (.A1(\V3/V2/V1/A2/M1/c1 ),
    .A2(\V3/V2/V1/A2/M1/c2 ),
    .ZN(\V3/V2/V1/A2/c1 ));
 AND2_X1 \V3/V2/V1/A2/M2/M1/_0_  (.A1(\V3/V2/V1/s1 [1]),
    .A2(\V3/V2/V1/v1 [3]),
    .ZN(\V3/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M2/M1/_1_  (.A(\V3/V2/V1/s1 [1]),
    .B(\V3/V2/V1/v1 [3]),
    .Z(\V3/V2/V1/A2/M2/s1 ));
 AND2_X1 \V3/V2/V1/A2/M2/M2/_0_  (.A1(\V3/V2/V1/A2/M2/s1 ),
    .A2(\V3/V2/V1/A2/c1 ),
    .ZN(\V3/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M2/M2/_1_  (.A(\V3/V2/V1/A2/M2/s1 ),
    .B(\V3/V2/V1/A2/c1 ),
    .Z(\V3/v2 [3]));
 OR2_X1 \V3/V2/V1/A2/M2/_0_  (.A1(\V3/V2/V1/A2/M2/c1 ),
    .A2(\V3/V2/V1/A2/M2/c2 ),
    .ZN(\V3/V2/V1/A2/c2 ));
 AND2_X1 \V3/V2/V1/A2/M3/M1/_0_  (.A1(\V3/V2/V1/s1 [2]),
    .A2(net5),
    .ZN(\V3/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M3/M1/_1_  (.A(\V3/V2/V1/s1 [2]),
    .B(net5),
    .Z(\V3/V2/V1/A2/M3/s1 ));
 AND2_X1 \V3/V2/V1/A2/M3/M2/_0_  (.A1(\V3/V2/V1/A2/M3/s1 ),
    .A2(\V3/V2/V1/A2/c2 ),
    .ZN(\V3/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M3/M2/_1_  (.A(\V3/V2/V1/A2/M3/s1 ),
    .B(\V3/V2/V1/A2/c2 ),
    .Z(\V3/V2/V1/s2 [2]));
 OR2_X1 \V3/V2/V1/A2/M3/_0_  (.A1(\V3/V2/V1/A2/M3/c1 ),
    .A2(\V3/V2/V1/A2/M3/c2 ),
    .ZN(\V3/V2/V1/A2/c3 ));
 AND2_X1 \V3/V2/V1/A2/M4/M1/_0_  (.A1(\V3/V2/V1/s1 [3]),
    .A2(net5),
    .ZN(\V3/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A2/M4/M1/_1_  (.A(\V3/V2/V1/s1 [3]),
    .B(net5),
    .Z(\V3/V2/V1/A2/M4/s1 ));
 AND2_X1 \V3/V2/V1/A2/M4/M2/_0_  (.A1(\V3/V2/V1/A2/M4/s1 ),
    .A2(\V3/V2/V1/A2/c3 ),
    .ZN(\V3/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A2/M4/M2/_1_  (.A(\V3/V2/V1/A2/M4/s1 ),
    .B(\V3/V2/V1/A2/c3 ),
    .Z(\V3/V2/V1/s2 [3]));
 OR2_X1 \V3/V2/V1/A2/M4/_0_  (.A1(\V3/V2/V1/A2/M4/c1 ),
    .A2(\V3/V2/V1/A2/M4/c2 ),
    .ZN(\V3/V2/V1/c2 ));
 AND2_X1 \V3/V2/V1/A3/M1/M1/_0_  (.A1(\V3/V2/V1/v4 [0]),
    .A2(\V3/V2/V1/s2 [2]),
    .ZN(\V3/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M1/M1/_1_  (.A(\V3/V2/V1/v4 [0]),
    .B(\V3/V2/V1/s2 [2]),
    .Z(\V3/V2/V1/A3/M1/s1 ));
 AND2_X1 \V3/V2/V1/A3/M1/M2/_0_  (.A1(\V3/V2/V1/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M1/M2/_1_  (.A(\V3/V2/V1/A3/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/v1 [4]));
 OR2_X1 \V3/V2/V1/A3/M1/_0_  (.A1(\V3/V2/V1/A3/M1/c1 ),
    .A2(\V3/V2/V1/A3/M1/c2 ),
    .ZN(\V3/V2/V1/A3/c1 ));
 AND2_X1 \V3/V2/V1/A3/M2/M1/_0_  (.A1(\V3/V2/V1/v4 [1]),
    .A2(\V3/V2/V1/s2 [3]),
    .ZN(\V3/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M2/M1/_1_  (.A(\V3/V2/V1/v4 [1]),
    .B(\V3/V2/V1/s2 [3]),
    .Z(\V3/V2/V1/A3/M2/s1 ));
 AND2_X1 \V3/V2/V1/A3/M2/M2/_0_  (.A1(\V3/V2/V1/A3/M2/s1 ),
    .A2(\V3/V2/V1/A3/c1 ),
    .ZN(\V3/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M2/M2/_1_  (.A(\V3/V2/V1/A3/M2/s1 ),
    .B(\V3/V2/V1/A3/c1 ),
    .Z(\V3/V2/v1 [5]));
 OR2_X1 \V3/V2/V1/A3/M2/_0_  (.A1(\V3/V2/V1/A3/M2/c1 ),
    .A2(\V3/V2/V1/A3/M2/c2 ),
    .ZN(\V3/V2/V1/A3/c2 ));
 AND2_X1 \V3/V2/V1/A3/M3/M1/_0_  (.A1(\V3/V2/V1/v4 [2]),
    .A2(\V3/V2/V1/c3 ),
    .ZN(\V3/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M3/M1/_1_  (.A(\V3/V2/V1/v4 [2]),
    .B(\V3/V2/V1/c3 ),
    .Z(\V3/V2/V1/A3/M3/s1 ));
 AND2_X1 \V3/V2/V1/A3/M3/M2/_0_  (.A1(\V3/V2/V1/A3/M3/s1 ),
    .A2(\V3/V2/V1/A3/c2 ),
    .ZN(\V3/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M3/M2/_1_  (.A(\V3/V2/V1/A3/M3/s1 ),
    .B(\V3/V2/V1/A3/c2 ),
    .Z(\V3/V2/v1 [6]));
 OR2_X1 \V3/V2/V1/A3/M3/_0_  (.A1(\V3/V2/V1/A3/M3/c1 ),
    .A2(\V3/V2/V1/A3/M3/c2 ),
    .ZN(\V3/V2/V1/A3/c3 ));
 AND2_X1 \V3/V2/V1/A3/M4/M1/_0_  (.A1(\V3/V2/V1/v4 [3]),
    .A2(net5),
    .ZN(\V3/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V1/A3/M4/M1/_1_  (.A(\V3/V2/V1/v4 [3]),
    .B(net5),
    .Z(\V3/V2/V1/A3/M4/s1 ));
 AND2_X1 \V3/V2/V1/A3/M4/M2/_0_  (.A1(\V3/V2/V1/A3/M4/s1 ),
    .A2(\V3/V2/V1/A3/c3 ),
    .ZN(\V3/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V1/A3/M4/M2/_1_  (.A(\V3/V2/V1/A3/M4/s1 ),
    .B(\V3/V2/V1/A3/c3 ),
    .Z(\V3/V2/v1 [7]));
 OR2_X1 \V3/V2/V1/A3/M4/_0_  (.A1(\V3/V2/V1/A3/M4/c1 ),
    .A2(\V3/V2/V1/A3/M4/c2 ),
    .ZN(\V3/V2/V1/overflow ));
 AND2_X1 \V3/V2/V1/V1/HA1/_0_  (.A1(\V3/V2/V1/V1/w2 ),
    .A2(\V3/V2/V1/V1/w1 ),
    .ZN(\V3/V2/V1/V1/w4 ));
 XOR2_X2 \V3/V2/V1/V1/HA1/_1_  (.A(\V3/V2/V1/V1/w2 ),
    .B(\V3/V2/V1/V1/w1 ),
    .Z(\V3/v2 [1]));
 AND2_X1 \V3/V2/V1/V1/HA2/_0_  (.A1(\V3/V2/V1/V1/w4 ),
    .A2(\V3/V2/V1/V1/w3 ),
    .ZN(\V3/V2/V1/v1 [3]));
 XOR2_X2 \V3/V2/V1/V1/HA2/_1_  (.A(\V3/V2/V1/V1/w4 ),
    .B(\V3/V2/V1/V1/w3 ),
    .Z(\V3/V2/V1/v1 [2]));
 AND2_X1 \V3/V2/V1/V1/_0_  (.A1(net25),
    .A2(B[16]),
    .ZN(\V3/v2 [0]));
 AND2_X1 \V3/V2/V1/V1/_1_  (.A1(net25),
    .A2(net21),
    .ZN(\V3/V2/V1/V1/w1 ));
 AND2_X1 \V3/V2/V1/V1/_2_  (.A1(B[16]),
    .A2(net24),
    .ZN(\V3/V2/V1/V1/w2 ));
 AND2_X1 \V3/V2/V1/V1/_3_  (.A1(net21),
    .A2(net24),
    .ZN(\V3/V2/V1/V1/w3 ));
 AND2_X1 \V3/V2/V1/V2/HA1/_0_  (.A1(\V3/V2/V1/V2/w2 ),
    .A2(\V3/V2/V1/V2/w1 ),
    .ZN(\V3/V2/V1/V2/w4 ));
 XOR2_X2 \V3/V2/V1/V2/HA1/_1_  (.A(\V3/V2/V1/V2/w2 ),
    .B(\V3/V2/V1/V2/w1 ),
    .Z(\V3/V2/V1/v2 [1]));
 AND2_X1 \V3/V2/V1/V2/HA2/_0_  (.A1(\V3/V2/V1/V2/w4 ),
    .A2(\V3/V2/V1/V2/w3 ),
    .ZN(\V3/V2/V1/v2 [3]));
 XOR2_X2 \V3/V2/V1/V2/HA2/_1_  (.A(\V3/V2/V1/V2/w4 ),
    .B(\V3/V2/V1/V2/w3 ),
    .Z(\V3/V2/V1/v2 [2]));
 AND2_X1 \V3/V2/V1/V2/_0_  (.A1(net47),
    .A2(B[16]),
    .ZN(\V3/V2/V1/v2 [0]));
 AND2_X1 \V3/V2/V1/V2/_1_  (.A1(net47),
    .A2(net21),
    .ZN(\V3/V2/V1/V2/w1 ));
 AND2_X1 \V3/V2/V1/V2/_2_  (.A1(B[16]),
    .A2(net46),
    .ZN(\V3/V2/V1/V2/w2 ));
 AND2_X1 \V3/V2/V1/V2/_3_  (.A1(net21),
    .A2(net46),
    .ZN(\V3/V2/V1/V2/w3 ));
 AND2_X1 \V3/V2/V1/V3/HA1/_0_  (.A1(\V3/V2/V1/V3/w2 ),
    .A2(\V3/V2/V1/V3/w1 ),
    .ZN(\V3/V2/V1/V3/w4 ));
 XOR2_X2 \V3/V2/V1/V3/HA1/_1_  (.A(\V3/V2/V1/V3/w2 ),
    .B(\V3/V2/V1/V3/w1 ),
    .Z(\V3/V2/V1/v3 [1]));
 AND2_X1 \V3/V2/V1/V3/HA2/_0_  (.A1(\V3/V2/V1/V3/w4 ),
    .A2(\V3/V2/V1/V3/w3 ),
    .ZN(\V3/V2/V1/v3 [3]));
 XOR2_X2 \V3/V2/V1/V3/HA2/_1_  (.A(\V3/V2/V1/V3/w4 ),
    .B(\V3/V2/V1/V3/w3 ),
    .Z(\V3/V2/V1/v3 [2]));
 AND2_X1 \V3/V2/V1/V3/_0_  (.A1(net25),
    .A2(net20),
    .ZN(\V3/V2/V1/v3 [0]));
 AND2_X1 \V3/V2/V1/V3/_1_  (.A1(net25),
    .A2(net19),
    .ZN(\V3/V2/V1/V3/w1 ));
 AND2_X1 \V3/V2/V1/V3/_2_  (.A1(net20),
    .A2(net24),
    .ZN(\V3/V2/V1/V3/w2 ));
 AND2_X1 \V3/V2/V1/V3/_3_  (.A1(net19),
    .A2(net24),
    .ZN(\V3/V2/V1/V3/w3 ));
 AND2_X1 \V3/V2/V1/V4/HA1/_0_  (.A1(\V3/V2/V1/V4/w2 ),
    .A2(\V3/V2/V1/V4/w1 ),
    .ZN(\V3/V2/V1/V4/w4 ));
 XOR2_X2 \V3/V2/V1/V4/HA1/_1_  (.A(\V3/V2/V1/V4/w2 ),
    .B(\V3/V2/V1/V4/w1 ),
    .Z(\V3/V2/V1/v4 [1]));
 AND2_X1 \V3/V2/V1/V4/HA2/_0_  (.A1(\V3/V2/V1/V4/w4 ),
    .A2(\V3/V2/V1/V4/w3 ),
    .ZN(\V3/V2/V1/v4 [3]));
 XOR2_X2 \V3/V2/V1/V4/HA2/_1_  (.A(\V3/V2/V1/V4/w4 ),
    .B(\V3/V2/V1/V4/w3 ),
    .Z(\V3/V2/V1/v4 [2]));
 AND2_X1 \V3/V2/V1/V4/_0_  (.A1(net47),
    .A2(net20),
    .ZN(\V3/V2/V1/v4 [0]));
 AND2_X1 \V3/V2/V1/V4/_1_  (.A1(net47),
    .A2(net19),
    .ZN(\V3/V2/V1/V4/w1 ));
 AND2_X1 \V3/V2/V1/V4/_2_  (.A1(net20),
    .A2(net46),
    .ZN(\V3/V2/V1/V4/w2 ));
 AND2_X1 \V3/V2/V1/V4/_3_  (.A1(net19),
    .A2(net46),
    .ZN(\V3/V2/V1/V4/w3 ));
 OR2_X1 \V3/V2/V1/_0_  (.A1(\V3/V2/V1/c1 ),
    .A2(\V3/V2/V1/c2 ),
    .ZN(\V3/V2/V1/c3 ));
 AND2_X1 \V3/V2/V2/A1/M1/M1/_0_  (.A1(\V3/V2/V2/v2 [0]),
    .A2(\V3/V2/V2/v3 [0]),
    .ZN(\V3/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M1/M1/_1_  (.A(\V3/V2/V2/v2 [0]),
    .B(\V3/V2/V2/v3 [0]),
    .Z(\V3/V2/V2/A1/M1/s1 ));
 AND2_X1 \V3/V2/V2/A1/M1/M2/_0_  (.A1(\V3/V2/V2/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M1/M2/_1_  (.A(\V3/V2/V2/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/V2/V2/s1 [0]));
 OR2_X1 \V3/V2/V2/A1/M1/_0_  (.A1(\V3/V2/V2/A1/M1/c1 ),
    .A2(\V3/V2/V2/A1/M1/c2 ),
    .ZN(\V3/V2/V2/A1/c1 ));
 AND2_X1 \V3/V2/V2/A1/M2/M1/_0_  (.A1(\V3/V2/V2/v2 [1]),
    .A2(\V3/V2/V2/v3 [1]),
    .ZN(\V3/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M2/M1/_1_  (.A(\V3/V2/V2/v2 [1]),
    .B(\V3/V2/V2/v3 [1]),
    .Z(\V3/V2/V2/A1/M2/s1 ));
 AND2_X1 \V3/V2/V2/A1/M2/M2/_0_  (.A1(\V3/V2/V2/A1/M2/s1 ),
    .A2(\V3/V2/V2/A1/c1 ),
    .ZN(\V3/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M2/M2/_1_  (.A(\V3/V2/V2/A1/M2/s1 ),
    .B(\V3/V2/V2/A1/c1 ),
    .Z(\V3/V2/V2/s1 [1]));
 OR2_X1 \V3/V2/V2/A1/M2/_0_  (.A1(\V3/V2/V2/A1/M2/c1 ),
    .A2(\V3/V2/V2/A1/M2/c2 ),
    .ZN(\V3/V2/V2/A1/c2 ));
 AND2_X1 \V3/V2/V2/A1/M3/M1/_0_  (.A1(\V3/V2/V2/v2 [2]),
    .A2(\V3/V2/V2/v3 [2]),
    .ZN(\V3/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M3/M1/_1_  (.A(\V3/V2/V2/v2 [2]),
    .B(\V3/V2/V2/v3 [2]),
    .Z(\V3/V2/V2/A1/M3/s1 ));
 AND2_X1 \V3/V2/V2/A1/M3/M2/_0_  (.A1(\V3/V2/V2/A1/M3/s1 ),
    .A2(\V3/V2/V2/A1/c2 ),
    .ZN(\V3/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M3/M2/_1_  (.A(\V3/V2/V2/A1/M3/s1 ),
    .B(\V3/V2/V2/A1/c2 ),
    .Z(\V3/V2/V2/s1 [2]));
 OR2_X1 \V3/V2/V2/A1/M3/_0_  (.A1(\V3/V2/V2/A1/M3/c1 ),
    .A2(\V3/V2/V2/A1/M3/c2 ),
    .ZN(\V3/V2/V2/A1/c3 ));
 AND2_X1 \V3/V2/V2/A1/M4/M1/_0_  (.A1(\V3/V2/V2/v2 [3]),
    .A2(\V3/V2/V2/v3 [3]),
    .ZN(\V3/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A1/M4/M1/_1_  (.A(\V3/V2/V2/v2 [3]),
    .B(\V3/V2/V2/v3 [3]),
    .Z(\V3/V2/V2/A1/M4/s1 ));
 AND2_X1 \V3/V2/V2/A1/M4/M2/_0_  (.A1(\V3/V2/V2/A1/M4/s1 ),
    .A2(\V3/V2/V2/A1/c3 ),
    .ZN(\V3/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A1/M4/M2/_1_  (.A(\V3/V2/V2/A1/M4/s1 ),
    .B(\V3/V2/V2/A1/c3 ),
    .Z(\V3/V2/V2/s1 [3]));
 OR2_X1 \V3/V2/V2/A1/M4/_0_  (.A1(\V3/V2/V2/A1/M4/c1 ),
    .A2(\V3/V2/V2/A1/M4/c2 ),
    .ZN(\V3/V2/V2/c1 ));
 AND2_X1 \V3/V2/V2/A2/M1/M1/_0_  (.A1(\V3/V2/V2/s1 [0]),
    .A2(\V3/V2/V2/v1 [2]),
    .ZN(\V3/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M1/M1/_1_  (.A(\V3/V2/V2/s1 [0]),
    .B(\V3/V2/V2/v1 [2]),
    .Z(\V3/V2/V2/A2/M1/s1 ));
 AND2_X1 \V3/V2/V2/A2/M1/M2/_0_  (.A1(\V3/V2/V2/A2/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M1/M2/_1_  (.A(\V3/V2/V2/A2/M1/s1 ),
    .B(net6),
    .Z(\V3/V2/v2 [2]));
 OR2_X1 \V3/V2/V2/A2/M1/_0_  (.A1(\V3/V2/V2/A2/M1/c1 ),
    .A2(\V3/V2/V2/A2/M1/c2 ),
    .ZN(\V3/V2/V2/A2/c1 ));
 AND2_X1 \V3/V2/V2/A2/M2/M1/_0_  (.A1(\V3/V2/V2/s1 [1]),
    .A2(\V3/V2/V2/v1 [3]),
    .ZN(\V3/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M2/M1/_1_  (.A(\V3/V2/V2/s1 [1]),
    .B(\V3/V2/V2/v1 [3]),
    .Z(\V3/V2/V2/A2/M2/s1 ));
 AND2_X1 \V3/V2/V2/A2/M2/M2/_0_  (.A1(\V3/V2/V2/A2/M2/s1 ),
    .A2(\V3/V2/V2/A2/c1 ),
    .ZN(\V3/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M2/M2/_1_  (.A(\V3/V2/V2/A2/M2/s1 ),
    .B(\V3/V2/V2/A2/c1 ),
    .Z(\V3/V2/v2 [3]));
 OR2_X1 \V3/V2/V2/A2/M2/_0_  (.A1(\V3/V2/V2/A2/M2/c1 ),
    .A2(\V3/V2/V2/A2/M2/c2 ),
    .ZN(\V3/V2/V2/A2/c2 ));
 AND2_X1 \V3/V2/V2/A2/M3/M1/_0_  (.A1(\V3/V2/V2/s1 [2]),
    .A2(net6),
    .ZN(\V3/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M3/M1/_1_  (.A(\V3/V2/V2/s1 [2]),
    .B(net6),
    .Z(\V3/V2/V2/A2/M3/s1 ));
 AND2_X1 \V3/V2/V2/A2/M3/M2/_0_  (.A1(\V3/V2/V2/A2/M3/s1 ),
    .A2(\V3/V2/V2/A2/c2 ),
    .ZN(\V3/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M3/M2/_1_  (.A(\V3/V2/V2/A2/M3/s1 ),
    .B(\V3/V2/V2/A2/c2 ),
    .Z(\V3/V2/V2/s2 [2]));
 OR2_X1 \V3/V2/V2/A2/M3/_0_  (.A1(\V3/V2/V2/A2/M3/c1 ),
    .A2(\V3/V2/V2/A2/M3/c2 ),
    .ZN(\V3/V2/V2/A2/c3 ));
 AND2_X1 \V3/V2/V2/A2/M4/M1/_0_  (.A1(\V3/V2/V2/s1 [3]),
    .A2(net6),
    .ZN(\V3/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A2/M4/M1/_1_  (.A(\V3/V2/V2/s1 [3]),
    .B(net6),
    .Z(\V3/V2/V2/A2/M4/s1 ));
 AND2_X1 \V3/V2/V2/A2/M4/M2/_0_  (.A1(\V3/V2/V2/A2/M4/s1 ),
    .A2(\V3/V2/V2/A2/c3 ),
    .ZN(\V3/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A2/M4/M2/_1_  (.A(\V3/V2/V2/A2/M4/s1 ),
    .B(\V3/V2/V2/A2/c3 ),
    .Z(\V3/V2/V2/s2 [3]));
 OR2_X1 \V3/V2/V2/A2/M4/_0_  (.A1(\V3/V2/V2/A2/M4/c1 ),
    .A2(\V3/V2/V2/A2/M4/c2 ),
    .ZN(\V3/V2/V2/c2 ));
 AND2_X1 \V3/V2/V2/A3/M1/M1/_0_  (.A1(\V3/V2/V2/v4 [0]),
    .A2(\V3/V2/V2/s2 [2]),
    .ZN(\V3/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M1/M1/_1_  (.A(\V3/V2/V2/v4 [0]),
    .B(\V3/V2/V2/s2 [2]),
    .Z(\V3/V2/V2/A3/M1/s1 ));
 AND2_X1 \V3/V2/V2/A3/M1/M2/_0_  (.A1(\V3/V2/V2/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M1/M2/_1_  (.A(\V3/V2/V2/A3/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/v2 [4]));
 OR2_X1 \V3/V2/V2/A3/M1/_0_  (.A1(\V3/V2/V2/A3/M1/c1 ),
    .A2(\V3/V2/V2/A3/M1/c2 ),
    .ZN(\V3/V2/V2/A3/c1 ));
 AND2_X1 \V3/V2/V2/A3/M2/M1/_0_  (.A1(\V3/V2/V2/v4 [1]),
    .A2(\V3/V2/V2/s2 [3]),
    .ZN(\V3/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M2/M1/_1_  (.A(\V3/V2/V2/v4 [1]),
    .B(\V3/V2/V2/s2 [3]),
    .Z(\V3/V2/V2/A3/M2/s1 ));
 AND2_X1 \V3/V2/V2/A3/M2/M2/_0_  (.A1(\V3/V2/V2/A3/M2/s1 ),
    .A2(\V3/V2/V2/A3/c1 ),
    .ZN(\V3/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M2/M2/_1_  (.A(\V3/V2/V2/A3/M2/s1 ),
    .B(\V3/V2/V2/A3/c1 ),
    .Z(\V3/V2/v2 [5]));
 OR2_X1 \V3/V2/V2/A3/M2/_0_  (.A1(\V3/V2/V2/A3/M2/c1 ),
    .A2(\V3/V2/V2/A3/M2/c2 ),
    .ZN(\V3/V2/V2/A3/c2 ));
 AND2_X1 \V3/V2/V2/A3/M3/M1/_0_  (.A1(\V3/V2/V2/v4 [2]),
    .A2(\V3/V2/V2/c3 ),
    .ZN(\V3/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M3/M1/_1_  (.A(\V3/V2/V2/v4 [2]),
    .B(\V3/V2/V2/c3 ),
    .Z(\V3/V2/V2/A3/M3/s1 ));
 AND2_X1 \V3/V2/V2/A3/M3/M2/_0_  (.A1(\V3/V2/V2/A3/M3/s1 ),
    .A2(\V3/V2/V2/A3/c2 ),
    .ZN(\V3/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M3/M2/_1_  (.A(\V3/V2/V2/A3/M3/s1 ),
    .B(\V3/V2/V2/A3/c2 ),
    .Z(\V3/V2/v2 [6]));
 OR2_X1 \V3/V2/V2/A3/M3/_0_  (.A1(\V3/V2/V2/A3/M3/c1 ),
    .A2(\V3/V2/V2/A3/M3/c2 ),
    .ZN(\V3/V2/V2/A3/c3 ));
 AND2_X1 \V3/V2/V2/A3/M4/M1/_0_  (.A1(\V3/V2/V2/v4 [3]),
    .A2(net6),
    .ZN(\V3/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V2/A3/M4/M1/_1_  (.A(\V3/V2/V2/v4 [3]),
    .B(net6),
    .Z(\V3/V2/V2/A3/M4/s1 ));
 AND2_X1 \V3/V2/V2/A3/M4/M2/_0_  (.A1(\V3/V2/V2/A3/M4/s1 ),
    .A2(\V3/V2/V2/A3/c3 ),
    .ZN(\V3/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V2/A3/M4/M2/_1_  (.A(\V3/V2/V2/A3/M4/s1 ),
    .B(\V3/V2/V2/A3/c3 ),
    .Z(\V3/V2/v2 [7]));
 OR2_X1 \V3/V2/V2/A3/M4/_0_  (.A1(\V3/V2/V2/A3/M4/c1 ),
    .A2(\V3/V2/V2/A3/M4/c2 ),
    .ZN(\V3/V2/V2/overflow ));
 AND2_X1 \V3/V2/V2/V1/HA1/_0_  (.A1(\V3/V2/V2/V1/w2 ),
    .A2(\V3/V2/V2/V1/w1 ),
    .ZN(\V3/V2/V2/V1/w4 ));
 XOR2_X2 \V3/V2/V2/V1/HA1/_1_  (.A(\V3/V2/V2/V1/w2 ),
    .B(\V3/V2/V2/V1/w1 ),
    .Z(\V3/V2/v2 [1]));
 AND2_X1 \V3/V2/V2/V1/HA2/_0_  (.A1(\V3/V2/V2/V1/w4 ),
    .A2(\V3/V2/V2/V1/w3 ),
    .ZN(\V3/V2/V2/v1 [3]));
 XOR2_X2 \V3/V2/V2/V1/HA2/_1_  (.A(\V3/V2/V2/V1/w4 ),
    .B(\V3/V2/V2/V1/w3 ),
    .Z(\V3/V2/V2/v1 [2]));
 AND2_X1 \V3/V2/V2/V1/_0_  (.A1(net45),
    .A2(B[16]),
    .ZN(\V3/V2/v2 [0]));
 AND2_X1 \V3/V2/V2/V1/_1_  (.A1(net45),
    .A2(net21),
    .ZN(\V3/V2/V2/V1/w1 ));
 AND2_X1 \V3/V2/V2/V1/_2_  (.A1(B[16]),
    .A2(net44),
    .ZN(\V3/V2/V2/V1/w2 ));
 AND2_X1 \V3/V2/V2/V1/_3_  (.A1(net21),
    .A2(net44),
    .ZN(\V3/V2/V2/V1/w3 ));
 AND2_X1 \V3/V2/V2/V2/HA1/_0_  (.A1(\V3/V2/V2/V2/w2 ),
    .A2(\V3/V2/V2/V2/w1 ),
    .ZN(\V3/V2/V2/V2/w4 ));
 XOR2_X2 \V3/V2/V2/V2/HA1/_1_  (.A(\V3/V2/V2/V2/w2 ),
    .B(\V3/V2/V2/V2/w1 ),
    .Z(\V3/V2/V2/v2 [1]));
 AND2_X1 \V3/V2/V2/V2/HA2/_0_  (.A1(\V3/V2/V2/V2/w4 ),
    .A2(\V3/V2/V2/V2/w3 ),
    .ZN(\V3/V2/V2/v2 [3]));
 XOR2_X2 \V3/V2/V2/V2/HA2/_1_  (.A(\V3/V2/V2/V2/w4 ),
    .B(\V3/V2/V2/V2/w3 ),
    .Z(\V3/V2/V2/v2 [2]));
 AND2_X1 \V3/V2/V2/V2/_0_  (.A1(net43),
    .A2(B[16]),
    .ZN(\V3/V2/V2/v2 [0]));
 AND2_X1 \V3/V2/V2/V2/_1_  (.A1(net43),
    .A2(net21),
    .ZN(\V3/V2/V2/V2/w1 ));
 AND2_X1 \V3/V2/V2/V2/_2_  (.A1(B[16]),
    .A2(net42),
    .ZN(\V3/V2/V2/V2/w2 ));
 AND2_X1 \V3/V2/V2/V2/_3_  (.A1(net21),
    .A2(net42),
    .ZN(\V3/V2/V2/V2/w3 ));
 AND2_X1 \V3/V2/V2/V3/HA1/_0_  (.A1(\V3/V2/V2/V3/w2 ),
    .A2(\V3/V2/V2/V3/w1 ),
    .ZN(\V3/V2/V2/V3/w4 ));
 XOR2_X2 \V3/V2/V2/V3/HA1/_1_  (.A(\V3/V2/V2/V3/w2 ),
    .B(\V3/V2/V2/V3/w1 ),
    .Z(\V3/V2/V2/v3 [1]));
 AND2_X1 \V3/V2/V2/V3/HA2/_0_  (.A1(\V3/V2/V2/V3/w4 ),
    .A2(\V3/V2/V2/V3/w3 ),
    .ZN(\V3/V2/V2/v3 [3]));
 XOR2_X2 \V3/V2/V2/V3/HA2/_1_  (.A(\V3/V2/V2/V3/w4 ),
    .B(\V3/V2/V2/V3/w3 ),
    .Z(\V3/V2/V2/v3 [2]));
 AND2_X1 \V3/V2/V2/V3/_0_  (.A1(net45),
    .A2(net20),
    .ZN(\V3/V2/V2/v3 [0]));
 AND2_X1 \V3/V2/V2/V3/_1_  (.A1(net45),
    .A2(net19),
    .ZN(\V3/V2/V2/V3/w1 ));
 AND2_X1 \V3/V2/V2/V3/_2_  (.A1(net20),
    .A2(net44),
    .ZN(\V3/V2/V2/V3/w2 ));
 AND2_X1 \V3/V2/V2/V3/_3_  (.A1(net19),
    .A2(net44),
    .ZN(\V3/V2/V2/V3/w3 ));
 AND2_X1 \V3/V2/V2/V4/HA1/_0_  (.A1(\V3/V2/V2/V4/w2 ),
    .A2(\V3/V2/V2/V4/w1 ),
    .ZN(\V3/V2/V2/V4/w4 ));
 XOR2_X2 \V3/V2/V2/V4/HA1/_1_  (.A(\V3/V2/V2/V4/w2 ),
    .B(\V3/V2/V2/V4/w1 ),
    .Z(\V3/V2/V2/v4 [1]));
 AND2_X1 \V3/V2/V2/V4/HA2/_0_  (.A1(\V3/V2/V2/V4/w4 ),
    .A2(\V3/V2/V2/V4/w3 ),
    .ZN(\V3/V2/V2/v4 [3]));
 XOR2_X2 \V3/V2/V2/V4/HA2/_1_  (.A(\V3/V2/V2/V4/w4 ),
    .B(\V3/V2/V2/V4/w3 ),
    .Z(\V3/V2/V2/v4 [2]));
 AND2_X1 \V3/V2/V2/V4/_0_  (.A1(net43),
    .A2(net20),
    .ZN(\V3/V2/V2/v4 [0]));
 AND2_X1 \V3/V2/V2/V4/_1_  (.A1(net43),
    .A2(net19),
    .ZN(\V3/V2/V2/V4/w1 ));
 AND2_X1 \V3/V2/V2/V4/_2_  (.A1(net20),
    .A2(net42),
    .ZN(\V3/V2/V2/V4/w2 ));
 AND2_X1 \V3/V2/V2/V4/_3_  (.A1(net19),
    .A2(net42),
    .ZN(\V3/V2/V2/V4/w3 ));
 OR2_X1 \V3/V2/V2/_0_  (.A1(\V3/V2/V2/c1 ),
    .A2(\V3/V2/V2/c2 ),
    .ZN(\V3/V2/V2/c3 ));
 AND2_X1 \V3/V2/V3/A1/M1/M1/_0_  (.A1(\V3/V2/V3/v2 [0]),
    .A2(\V3/V2/V3/v3 [0]),
    .ZN(\V3/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M1/M1/_1_  (.A(\V3/V2/V3/v2 [0]),
    .B(\V3/V2/V3/v3 [0]),
    .Z(\V3/V2/V3/A1/M1/s1 ));
 AND2_X1 \V3/V2/V3/A1/M1/M2/_0_  (.A1(\V3/V2/V3/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M1/M2/_1_  (.A(\V3/V2/V3/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/V3/s1 [0]));
 OR2_X1 \V3/V2/V3/A1/M1/_0_  (.A1(\V3/V2/V3/A1/M1/c1 ),
    .A2(\V3/V2/V3/A1/M1/c2 ),
    .ZN(\V3/V2/V3/A1/c1 ));
 AND2_X1 \V3/V2/V3/A1/M2/M1/_0_  (.A1(\V3/V2/V3/v2 [1]),
    .A2(\V3/V2/V3/v3 [1]),
    .ZN(\V3/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M2/M1/_1_  (.A(\V3/V2/V3/v2 [1]),
    .B(\V3/V2/V3/v3 [1]),
    .Z(\V3/V2/V3/A1/M2/s1 ));
 AND2_X1 \V3/V2/V3/A1/M2/M2/_0_  (.A1(\V3/V2/V3/A1/M2/s1 ),
    .A2(\V3/V2/V3/A1/c1 ),
    .ZN(\V3/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M2/M2/_1_  (.A(\V3/V2/V3/A1/M2/s1 ),
    .B(\V3/V2/V3/A1/c1 ),
    .Z(\V3/V2/V3/s1 [1]));
 OR2_X1 \V3/V2/V3/A1/M2/_0_  (.A1(\V3/V2/V3/A1/M2/c1 ),
    .A2(\V3/V2/V3/A1/M2/c2 ),
    .ZN(\V3/V2/V3/A1/c2 ));
 AND2_X1 \V3/V2/V3/A1/M3/M1/_0_  (.A1(\V3/V2/V3/v2 [2]),
    .A2(\V3/V2/V3/v3 [2]),
    .ZN(\V3/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M3/M1/_1_  (.A(\V3/V2/V3/v2 [2]),
    .B(\V3/V2/V3/v3 [2]),
    .Z(\V3/V2/V3/A1/M3/s1 ));
 AND2_X1 \V3/V2/V3/A1/M3/M2/_0_  (.A1(\V3/V2/V3/A1/M3/s1 ),
    .A2(\V3/V2/V3/A1/c2 ),
    .ZN(\V3/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M3/M2/_1_  (.A(\V3/V2/V3/A1/M3/s1 ),
    .B(\V3/V2/V3/A1/c2 ),
    .Z(\V3/V2/V3/s1 [2]));
 OR2_X1 \V3/V2/V3/A1/M3/_0_  (.A1(\V3/V2/V3/A1/M3/c1 ),
    .A2(\V3/V2/V3/A1/M3/c2 ),
    .ZN(\V3/V2/V3/A1/c3 ));
 AND2_X1 \V3/V2/V3/A1/M4/M1/_0_  (.A1(\V3/V2/V3/v2 [3]),
    .A2(\V3/V2/V3/v3 [3]),
    .ZN(\V3/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A1/M4/M1/_1_  (.A(\V3/V2/V3/v2 [3]),
    .B(\V3/V2/V3/v3 [3]),
    .Z(\V3/V2/V3/A1/M4/s1 ));
 AND2_X1 \V3/V2/V3/A1/M4/M2/_0_  (.A1(\V3/V2/V3/A1/M4/s1 ),
    .A2(\V3/V2/V3/A1/c3 ),
    .ZN(\V3/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A1/M4/M2/_1_  (.A(\V3/V2/V3/A1/M4/s1 ),
    .B(\V3/V2/V3/A1/c3 ),
    .Z(\V3/V2/V3/s1 [3]));
 OR2_X1 \V3/V2/V3/A1/M4/_0_  (.A1(\V3/V2/V3/A1/M4/c1 ),
    .A2(\V3/V2/V3/A1/M4/c2 ),
    .ZN(\V3/V2/V3/c1 ));
 AND2_X1 \V3/V2/V3/A2/M1/M1/_0_  (.A1(\V3/V2/V3/s1 [0]),
    .A2(\V3/V2/V3/v1 [2]),
    .ZN(\V3/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M1/M1/_1_  (.A(\V3/V2/V3/s1 [0]),
    .B(\V3/V2/V3/v1 [2]),
    .Z(\V3/V2/V3/A2/M1/s1 ));
 AND2_X1 \V3/V2/V3/A2/M1/M2/_0_  (.A1(\V3/V2/V3/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M1/M2/_1_  (.A(\V3/V2/V3/A2/M1/s1 ),
    .B(net6),
    .Z(\V3/V2/v3 [2]));
 OR2_X1 \V3/V2/V3/A2/M1/_0_  (.A1(\V3/V2/V3/A2/M1/c1 ),
    .A2(\V3/V2/V3/A2/M1/c2 ),
    .ZN(\V3/V2/V3/A2/c1 ));
 AND2_X1 \V3/V2/V3/A2/M2/M1/_0_  (.A1(\V3/V2/V3/s1 [1]),
    .A2(\V3/V2/V3/v1 [3]),
    .ZN(\V3/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M2/M1/_1_  (.A(\V3/V2/V3/s1 [1]),
    .B(\V3/V2/V3/v1 [3]),
    .Z(\V3/V2/V3/A2/M2/s1 ));
 AND2_X1 \V3/V2/V3/A2/M2/M2/_0_  (.A1(\V3/V2/V3/A2/M2/s1 ),
    .A2(\V3/V2/V3/A2/c1 ),
    .ZN(\V3/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M2/M2/_1_  (.A(\V3/V2/V3/A2/M2/s1 ),
    .B(\V3/V2/V3/A2/c1 ),
    .Z(\V3/V2/v3 [3]));
 OR2_X1 \V3/V2/V3/A2/M2/_0_  (.A1(\V3/V2/V3/A2/M2/c1 ),
    .A2(\V3/V2/V3/A2/M2/c2 ),
    .ZN(\V3/V2/V3/A2/c2 ));
 AND2_X1 \V3/V2/V3/A2/M3/M1/_0_  (.A1(\V3/V2/V3/s1 [2]),
    .A2(net5),
    .ZN(\V3/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M3/M1/_1_  (.A(\V3/V2/V3/s1 [2]),
    .B(net5),
    .Z(\V3/V2/V3/A2/M3/s1 ));
 AND2_X1 \V3/V2/V3/A2/M3/M2/_0_  (.A1(\V3/V2/V3/A2/M3/s1 ),
    .A2(\V3/V2/V3/A2/c2 ),
    .ZN(\V3/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M3/M2/_1_  (.A(\V3/V2/V3/A2/M3/s1 ),
    .B(\V3/V2/V3/A2/c2 ),
    .Z(\V3/V2/V3/s2 [2]));
 OR2_X1 \V3/V2/V3/A2/M3/_0_  (.A1(\V3/V2/V3/A2/M3/c1 ),
    .A2(\V3/V2/V3/A2/M3/c2 ),
    .ZN(\V3/V2/V3/A2/c3 ));
 AND2_X1 \V3/V2/V3/A2/M4/M1/_0_  (.A1(\V3/V2/V3/s1 [3]),
    .A2(net5),
    .ZN(\V3/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A2/M4/M1/_1_  (.A(\V3/V2/V3/s1 [3]),
    .B(net5),
    .Z(\V3/V2/V3/A2/M4/s1 ));
 AND2_X1 \V3/V2/V3/A2/M4/M2/_0_  (.A1(\V3/V2/V3/A2/M4/s1 ),
    .A2(\V3/V2/V3/A2/c3 ),
    .ZN(\V3/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A2/M4/M2/_1_  (.A(\V3/V2/V3/A2/M4/s1 ),
    .B(\V3/V2/V3/A2/c3 ),
    .Z(\V3/V2/V3/s2 [3]));
 OR2_X1 \V3/V2/V3/A2/M4/_0_  (.A1(\V3/V2/V3/A2/M4/c1 ),
    .A2(\V3/V2/V3/A2/M4/c2 ),
    .ZN(\V3/V2/V3/c2 ));
 AND2_X1 \V3/V2/V3/A3/M1/M1/_0_  (.A1(\V3/V2/V3/v4 [0]),
    .A2(\V3/V2/V3/s2 [2]),
    .ZN(\V3/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M1/M1/_1_  (.A(\V3/V2/V3/v4 [0]),
    .B(\V3/V2/V3/s2 [2]),
    .Z(\V3/V2/V3/A3/M1/s1 ));
 AND2_X1 \V3/V2/V3/A3/M1/M2/_0_  (.A1(\V3/V2/V3/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M1/M2/_1_  (.A(\V3/V2/V3/A3/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/v3 [4]));
 OR2_X1 \V3/V2/V3/A3/M1/_0_  (.A1(\V3/V2/V3/A3/M1/c1 ),
    .A2(\V3/V2/V3/A3/M1/c2 ),
    .ZN(\V3/V2/V3/A3/c1 ));
 AND2_X1 \V3/V2/V3/A3/M2/M1/_0_  (.A1(\V3/V2/V3/v4 [1]),
    .A2(\V3/V2/V3/s2 [3]),
    .ZN(\V3/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M2/M1/_1_  (.A(\V3/V2/V3/v4 [1]),
    .B(\V3/V2/V3/s2 [3]),
    .Z(\V3/V2/V3/A3/M2/s1 ));
 AND2_X1 \V3/V2/V3/A3/M2/M2/_0_  (.A1(\V3/V2/V3/A3/M2/s1 ),
    .A2(\V3/V2/V3/A3/c1 ),
    .ZN(\V3/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M2/M2/_1_  (.A(\V3/V2/V3/A3/M2/s1 ),
    .B(\V3/V2/V3/A3/c1 ),
    .Z(\V3/V2/v3 [5]));
 OR2_X1 \V3/V2/V3/A3/M2/_0_  (.A1(\V3/V2/V3/A3/M2/c1 ),
    .A2(\V3/V2/V3/A3/M2/c2 ),
    .ZN(\V3/V2/V3/A3/c2 ));
 AND2_X1 \V3/V2/V3/A3/M3/M1/_0_  (.A1(\V3/V2/V3/v4 [2]),
    .A2(\V3/V2/V3/c3 ),
    .ZN(\V3/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M3/M1/_1_  (.A(\V3/V2/V3/v4 [2]),
    .B(\V3/V2/V3/c3 ),
    .Z(\V3/V2/V3/A3/M3/s1 ));
 AND2_X1 \V3/V2/V3/A3/M3/M2/_0_  (.A1(\V3/V2/V3/A3/M3/s1 ),
    .A2(\V3/V2/V3/A3/c2 ),
    .ZN(\V3/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M3/M2/_1_  (.A(\V3/V2/V3/A3/M3/s1 ),
    .B(\V3/V2/V3/A3/c2 ),
    .Z(\V3/V2/v3 [6]));
 OR2_X1 \V3/V2/V3/A3/M3/_0_  (.A1(\V3/V2/V3/A3/M3/c1 ),
    .A2(\V3/V2/V3/A3/M3/c2 ),
    .ZN(\V3/V2/V3/A3/c3 ));
 AND2_X1 \V3/V2/V3/A3/M4/M1/_0_  (.A1(\V3/V2/V3/v4 [3]),
    .A2(net6),
    .ZN(\V3/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V3/A3/M4/M1/_1_  (.A(\V3/V2/V3/v4 [3]),
    .B(net6),
    .Z(\V3/V2/V3/A3/M4/s1 ));
 AND2_X1 \V3/V2/V3/A3/M4/M2/_0_  (.A1(\V3/V2/V3/A3/M4/s1 ),
    .A2(\V3/V2/V3/A3/c3 ),
    .ZN(\V3/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V3/A3/M4/M2/_1_  (.A(\V3/V2/V3/A3/M4/s1 ),
    .B(\V3/V2/V3/A3/c3 ),
    .Z(\V3/V2/v3 [7]));
 OR2_X1 \V3/V2/V3/A3/M4/_0_  (.A1(\V3/V2/V3/A3/M4/c1 ),
    .A2(\V3/V2/V3/A3/M4/c2 ),
    .ZN(\V3/V2/V3/overflow ));
 AND2_X1 \V3/V2/V3/V1/HA1/_0_  (.A1(\V3/V2/V3/V1/w2 ),
    .A2(\V3/V2/V3/V1/w1 ),
    .ZN(\V3/V2/V3/V1/w4 ));
 XOR2_X2 \V3/V2/V3/V1/HA1/_1_  (.A(\V3/V2/V3/V1/w2 ),
    .B(\V3/V2/V3/V1/w1 ),
    .Z(\V3/V2/v3 [1]));
 AND2_X1 \V3/V2/V3/V1/HA2/_0_  (.A1(\V3/V2/V3/V1/w4 ),
    .A2(\V3/V2/V3/V1/w3 ),
    .ZN(\V3/V2/V3/v1 [3]));
 XOR2_X2 \V3/V2/V3/V1/HA2/_1_  (.A(\V3/V2/V3/V1/w4 ),
    .B(\V3/V2/V3/V1/w3 ),
    .Z(\V3/V2/V3/v1 [2]));
 AND2_X1 \V3/V2/V3/V1/_0_  (.A1(net25),
    .A2(net18),
    .ZN(\V3/V2/v3 [0]));
 AND2_X1 \V3/V2/V3/V1/_1_  (.A1(net25),
    .A2(net17),
    .ZN(\V3/V2/V3/V1/w1 ));
 AND2_X1 \V3/V2/V3/V1/_2_  (.A1(net18),
    .A2(net24),
    .ZN(\V3/V2/V3/V1/w2 ));
 AND2_X1 \V3/V2/V3/V1/_3_  (.A1(net17),
    .A2(net24),
    .ZN(\V3/V2/V3/V1/w3 ));
 AND2_X1 \V3/V2/V3/V2/HA1/_0_  (.A1(\V3/V2/V3/V2/w2 ),
    .A2(\V3/V2/V3/V2/w1 ),
    .ZN(\V3/V2/V3/V2/w4 ));
 XOR2_X2 \V3/V2/V3/V2/HA1/_1_  (.A(\V3/V2/V3/V2/w2 ),
    .B(\V3/V2/V3/V2/w1 ),
    .Z(\V3/V2/V3/v2 [1]));
 AND2_X1 \V3/V2/V3/V2/HA2/_0_  (.A1(\V3/V2/V3/V2/w4 ),
    .A2(\V3/V2/V3/V2/w3 ),
    .ZN(\V3/V2/V3/v2 [3]));
 XOR2_X2 \V3/V2/V3/V2/HA2/_1_  (.A(\V3/V2/V3/V2/w4 ),
    .B(\V3/V2/V3/V2/w3 ),
    .Z(\V3/V2/V3/v2 [2]));
 AND2_X1 \V3/V2/V3/V2/_0_  (.A1(net47),
    .A2(net18),
    .ZN(\V3/V2/V3/v2 [0]));
 AND2_X1 \V3/V2/V3/V2/_1_  (.A1(net47),
    .A2(net17),
    .ZN(\V3/V2/V3/V2/w1 ));
 AND2_X1 \V3/V2/V3/V2/_2_  (.A1(net18),
    .A2(net46),
    .ZN(\V3/V2/V3/V2/w2 ));
 AND2_X1 \V3/V2/V3/V2/_3_  (.A1(net17),
    .A2(net46),
    .ZN(\V3/V2/V3/V2/w3 ));
 AND2_X1 \V3/V2/V3/V3/HA1/_0_  (.A1(\V3/V2/V3/V3/w2 ),
    .A2(\V3/V2/V3/V3/w1 ),
    .ZN(\V3/V2/V3/V3/w4 ));
 XOR2_X2 \V3/V2/V3/V3/HA1/_1_  (.A(\V3/V2/V3/V3/w2 ),
    .B(\V3/V2/V3/V3/w1 ),
    .Z(\V3/V2/V3/v3 [1]));
 AND2_X1 \V3/V2/V3/V3/HA2/_0_  (.A1(\V3/V2/V3/V3/w4 ),
    .A2(\V3/V2/V3/V3/w3 ),
    .ZN(\V3/V2/V3/v3 [3]));
 XOR2_X2 \V3/V2/V3/V3/HA2/_1_  (.A(\V3/V2/V3/V3/w4 ),
    .B(\V3/V2/V3/V3/w3 ),
    .Z(\V3/V2/V3/v3 [2]));
 AND2_X1 \V3/V2/V3/V3/_0_  (.A1(net25),
    .A2(net16),
    .ZN(\V3/V2/V3/v3 [0]));
 AND2_X1 \V3/V2/V3/V3/_1_  (.A1(net25),
    .A2(net15),
    .ZN(\V3/V2/V3/V3/w1 ));
 AND2_X1 \V3/V2/V3/V3/_2_  (.A1(net16),
    .A2(net24),
    .ZN(\V3/V2/V3/V3/w2 ));
 AND2_X1 \V3/V2/V3/V3/_3_  (.A1(net15),
    .A2(net24),
    .ZN(\V3/V2/V3/V3/w3 ));
 AND2_X1 \V3/V2/V3/V4/HA1/_0_  (.A1(\V3/V2/V3/V4/w2 ),
    .A2(\V3/V2/V3/V4/w1 ),
    .ZN(\V3/V2/V3/V4/w4 ));
 XOR2_X2 \V3/V2/V3/V4/HA1/_1_  (.A(\V3/V2/V3/V4/w2 ),
    .B(\V3/V2/V3/V4/w1 ),
    .Z(\V3/V2/V3/v4 [1]));
 AND2_X1 \V3/V2/V3/V4/HA2/_0_  (.A1(\V3/V2/V3/V4/w4 ),
    .A2(\V3/V2/V3/V4/w3 ),
    .ZN(\V3/V2/V3/v4 [3]));
 XOR2_X2 \V3/V2/V3/V4/HA2/_1_  (.A(\V3/V2/V3/V4/w4 ),
    .B(\V3/V2/V3/V4/w3 ),
    .Z(\V3/V2/V3/v4 [2]));
 AND2_X1 \V3/V2/V3/V4/_0_  (.A1(net47),
    .A2(net16),
    .ZN(\V3/V2/V3/v4 [0]));
 AND2_X1 \V3/V2/V3/V4/_1_  (.A1(net47),
    .A2(net15),
    .ZN(\V3/V2/V3/V4/w1 ));
 AND2_X1 \V3/V2/V3/V4/_2_  (.A1(net16),
    .A2(net46),
    .ZN(\V3/V2/V3/V4/w2 ));
 AND2_X1 \V3/V2/V3/V4/_3_  (.A1(net15),
    .A2(net46),
    .ZN(\V3/V2/V3/V4/w3 ));
 OR2_X1 \V3/V2/V3/_0_  (.A1(\V3/V2/V3/c1 ),
    .A2(\V3/V2/V3/c2 ),
    .ZN(\V3/V2/V3/c3 ));
 AND2_X1 \V3/V2/V4/A1/M1/M1/_0_  (.A1(\V3/V2/V4/v2 [0]),
    .A2(\V3/V2/V4/v3 [0]),
    .ZN(\V3/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M1/M1/_1_  (.A(\V3/V2/V4/v2 [0]),
    .B(\V3/V2/V4/v3 [0]),
    .Z(\V3/V2/V4/A1/M1/s1 ));
 AND2_X1 \V3/V2/V4/A1/M1/M2/_0_  (.A1(\V3/V2/V4/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M1/M2/_1_  (.A(\V3/V2/V4/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/V4/s1 [0]));
 OR2_X1 \V3/V2/V4/A1/M1/_0_  (.A1(\V3/V2/V4/A1/M1/c1 ),
    .A2(\V3/V2/V4/A1/M1/c2 ),
    .ZN(\V3/V2/V4/A1/c1 ));
 AND2_X1 \V3/V2/V4/A1/M2/M1/_0_  (.A1(\V3/V2/V4/v2 [1]),
    .A2(\V3/V2/V4/v3 [1]),
    .ZN(\V3/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M2/M1/_1_  (.A(\V3/V2/V4/v2 [1]),
    .B(\V3/V2/V4/v3 [1]),
    .Z(\V3/V2/V4/A1/M2/s1 ));
 AND2_X1 \V3/V2/V4/A1/M2/M2/_0_  (.A1(\V3/V2/V4/A1/M2/s1 ),
    .A2(\V3/V2/V4/A1/c1 ),
    .ZN(\V3/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M2/M2/_1_  (.A(\V3/V2/V4/A1/M2/s1 ),
    .B(\V3/V2/V4/A1/c1 ),
    .Z(\V3/V2/V4/s1 [1]));
 OR2_X1 \V3/V2/V4/A1/M2/_0_  (.A1(\V3/V2/V4/A1/M2/c1 ),
    .A2(\V3/V2/V4/A1/M2/c2 ),
    .ZN(\V3/V2/V4/A1/c2 ));
 AND2_X1 \V3/V2/V4/A1/M3/M1/_0_  (.A1(\V3/V2/V4/v2 [2]),
    .A2(\V3/V2/V4/v3 [2]),
    .ZN(\V3/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M3/M1/_1_  (.A(\V3/V2/V4/v2 [2]),
    .B(\V3/V2/V4/v3 [2]),
    .Z(\V3/V2/V4/A1/M3/s1 ));
 AND2_X1 \V3/V2/V4/A1/M3/M2/_0_  (.A1(\V3/V2/V4/A1/M3/s1 ),
    .A2(\V3/V2/V4/A1/c2 ),
    .ZN(\V3/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M3/M2/_1_  (.A(\V3/V2/V4/A1/M3/s1 ),
    .B(\V3/V2/V4/A1/c2 ),
    .Z(\V3/V2/V4/s1 [2]));
 OR2_X1 \V3/V2/V4/A1/M3/_0_  (.A1(\V3/V2/V4/A1/M3/c1 ),
    .A2(\V3/V2/V4/A1/M3/c2 ),
    .ZN(\V3/V2/V4/A1/c3 ));
 AND2_X1 \V3/V2/V4/A1/M4/M1/_0_  (.A1(\V3/V2/V4/v2 [3]),
    .A2(\V3/V2/V4/v3 [3]),
    .ZN(\V3/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A1/M4/M1/_1_  (.A(\V3/V2/V4/v2 [3]),
    .B(\V3/V2/V4/v3 [3]),
    .Z(\V3/V2/V4/A1/M4/s1 ));
 AND2_X1 \V3/V2/V4/A1/M4/M2/_0_  (.A1(\V3/V2/V4/A1/M4/s1 ),
    .A2(\V3/V2/V4/A1/c3 ),
    .ZN(\V3/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A1/M4/M2/_1_  (.A(\V3/V2/V4/A1/M4/s1 ),
    .B(\V3/V2/V4/A1/c3 ),
    .Z(\V3/V2/V4/s1 [3]));
 OR2_X1 \V3/V2/V4/A1/M4/_0_  (.A1(\V3/V2/V4/A1/M4/c1 ),
    .A2(\V3/V2/V4/A1/M4/c2 ),
    .ZN(\V3/V2/V4/c1 ));
 AND2_X1 \V3/V2/V4/A2/M1/M1/_0_  (.A1(\V3/V2/V4/s1 [0]),
    .A2(\V3/V2/V4/v1 [2]),
    .ZN(\V3/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M1/M1/_1_  (.A(\V3/V2/V4/s1 [0]),
    .B(\V3/V2/V4/v1 [2]),
    .Z(\V3/V2/V4/A2/M1/s1 ));
 AND2_X1 \V3/V2/V4/A2/M1/M2/_0_  (.A1(\V3/V2/V4/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M1/M2/_1_  (.A(\V3/V2/V4/A2/M1/s1 ),
    .B(net5),
    .Z(\V3/V2/v4 [2]));
 OR2_X1 \V3/V2/V4/A2/M1/_0_  (.A1(\V3/V2/V4/A2/M1/c1 ),
    .A2(\V3/V2/V4/A2/M1/c2 ),
    .ZN(\V3/V2/V4/A2/c1 ));
 AND2_X1 \V3/V2/V4/A2/M2/M1/_0_  (.A1(\V3/V2/V4/s1 [1]),
    .A2(\V3/V2/V4/v1 [3]),
    .ZN(\V3/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M2/M1/_1_  (.A(\V3/V2/V4/s1 [1]),
    .B(\V3/V2/V4/v1 [3]),
    .Z(\V3/V2/V4/A2/M2/s1 ));
 AND2_X1 \V3/V2/V4/A2/M2/M2/_0_  (.A1(\V3/V2/V4/A2/M2/s1 ),
    .A2(\V3/V2/V4/A2/c1 ),
    .ZN(\V3/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M2/M2/_1_  (.A(\V3/V2/V4/A2/M2/s1 ),
    .B(\V3/V2/V4/A2/c1 ),
    .Z(\V3/V2/v4 [3]));
 OR2_X1 \V3/V2/V4/A2/M2/_0_  (.A1(\V3/V2/V4/A2/M2/c1 ),
    .A2(\V3/V2/V4/A2/M2/c2 ),
    .ZN(\V3/V2/V4/A2/c2 ));
 AND2_X1 \V3/V2/V4/A2/M3/M1/_0_  (.A1(\V3/V2/V4/s1 [2]),
    .A2(net5),
    .ZN(\V3/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M3/M1/_1_  (.A(\V3/V2/V4/s1 [2]),
    .B(net5),
    .Z(\V3/V2/V4/A2/M3/s1 ));
 AND2_X1 \V3/V2/V4/A2/M3/M2/_0_  (.A1(\V3/V2/V4/A2/M3/s1 ),
    .A2(\V3/V2/V4/A2/c2 ),
    .ZN(\V3/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M3/M2/_1_  (.A(\V3/V2/V4/A2/M3/s1 ),
    .B(\V3/V2/V4/A2/c2 ),
    .Z(\V3/V2/V4/s2 [2]));
 OR2_X1 \V3/V2/V4/A2/M3/_0_  (.A1(\V3/V2/V4/A2/M3/c1 ),
    .A2(\V3/V2/V4/A2/M3/c2 ),
    .ZN(\V3/V2/V4/A2/c3 ));
 AND2_X1 \V3/V2/V4/A2/M4/M1/_0_  (.A1(\V3/V2/V4/s1 [3]),
    .A2(net8),
    .ZN(\V3/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A2/M4/M1/_1_  (.A(\V3/V2/V4/s1 [3]),
    .B(net8),
    .Z(\V3/V2/V4/A2/M4/s1 ));
 AND2_X1 \V3/V2/V4/A2/M4/M2/_0_  (.A1(\V3/V2/V4/A2/M4/s1 ),
    .A2(\V3/V2/V4/A2/c3 ),
    .ZN(\V3/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A2/M4/M2/_1_  (.A(\V3/V2/V4/A2/M4/s1 ),
    .B(\V3/V2/V4/A2/c3 ),
    .Z(\V3/V2/V4/s2 [3]));
 OR2_X1 \V3/V2/V4/A2/M4/_0_  (.A1(\V3/V2/V4/A2/M4/c1 ),
    .A2(\V3/V2/V4/A2/M4/c2 ),
    .ZN(\V3/V2/V4/c2 ));
 AND2_X1 \V3/V2/V4/A3/M1/M1/_0_  (.A1(\V3/V2/V4/v4 [0]),
    .A2(\V3/V2/V4/s2 [2]),
    .ZN(\V3/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M1/M1/_1_  (.A(\V3/V2/V4/v4 [0]),
    .B(\V3/V2/V4/s2 [2]),
    .Z(\V3/V2/V4/A3/M1/s1 ));
 AND2_X1 \V3/V2/V4/A3/M1/M2/_0_  (.A1(\V3/V2/V4/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M1/M2/_1_  (.A(\V3/V2/V4/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V2/v4 [4]));
 OR2_X1 \V3/V2/V4/A3/M1/_0_  (.A1(\V3/V2/V4/A3/M1/c1 ),
    .A2(\V3/V2/V4/A3/M1/c2 ),
    .ZN(\V3/V2/V4/A3/c1 ));
 AND2_X1 \V3/V2/V4/A3/M2/M1/_0_  (.A1(\V3/V2/V4/v4 [1]),
    .A2(\V3/V2/V4/s2 [3]),
    .ZN(\V3/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M2/M1/_1_  (.A(\V3/V2/V4/v4 [1]),
    .B(\V3/V2/V4/s2 [3]),
    .Z(\V3/V2/V4/A3/M2/s1 ));
 AND2_X1 \V3/V2/V4/A3/M2/M2/_0_  (.A1(\V3/V2/V4/A3/M2/s1 ),
    .A2(\V3/V2/V4/A3/c1 ),
    .ZN(\V3/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M2/M2/_1_  (.A(\V3/V2/V4/A3/M2/s1 ),
    .B(\V3/V2/V4/A3/c1 ),
    .Z(\V3/V2/v4 [5]));
 OR2_X1 \V3/V2/V4/A3/M2/_0_  (.A1(\V3/V2/V4/A3/M2/c1 ),
    .A2(\V3/V2/V4/A3/M2/c2 ),
    .ZN(\V3/V2/V4/A3/c2 ));
 AND2_X1 \V3/V2/V4/A3/M3/M1/_0_  (.A1(\V3/V2/V4/v4 [2]),
    .A2(\V3/V2/V4/c3 ),
    .ZN(\V3/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M3/M1/_1_  (.A(\V3/V2/V4/v4 [2]),
    .B(\V3/V2/V4/c3 ),
    .Z(\V3/V2/V4/A3/M3/s1 ));
 AND2_X1 \V3/V2/V4/A3/M3/M2/_0_  (.A1(\V3/V2/V4/A3/M3/s1 ),
    .A2(\V3/V2/V4/A3/c2 ),
    .ZN(\V3/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M3/M2/_1_  (.A(\V3/V2/V4/A3/M3/s1 ),
    .B(\V3/V2/V4/A3/c2 ),
    .Z(\V3/V2/v4 [6]));
 OR2_X1 \V3/V2/V4/A3/M3/_0_  (.A1(\V3/V2/V4/A3/M3/c1 ),
    .A2(\V3/V2/V4/A3/M3/c2 ),
    .ZN(\V3/V2/V4/A3/c3 ));
 AND2_X1 \V3/V2/V4/A3/M4/M1/_0_  (.A1(\V3/V2/V4/v4 [3]),
    .A2(net8),
    .ZN(\V3/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V2/V4/A3/M4/M1/_1_  (.A(\V3/V2/V4/v4 [3]),
    .B(net8),
    .Z(\V3/V2/V4/A3/M4/s1 ));
 AND2_X1 \V3/V2/V4/A3/M4/M2/_0_  (.A1(\V3/V2/V4/A3/M4/s1 ),
    .A2(\V3/V2/V4/A3/c3 ),
    .ZN(\V3/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V2/V4/A3/M4/M2/_1_  (.A(\V3/V2/V4/A3/M4/s1 ),
    .B(\V3/V2/V4/A3/c3 ),
    .Z(\V3/V2/v4 [7]));
 OR2_X1 \V3/V2/V4/A3/M4/_0_  (.A1(\V3/V2/V4/A3/M4/c1 ),
    .A2(\V3/V2/V4/A3/M4/c2 ),
    .ZN(\V3/V2/V4/overflow ));
 AND2_X1 \V3/V2/V4/V1/HA1/_0_  (.A1(\V3/V2/V4/V1/w2 ),
    .A2(\V3/V2/V4/V1/w1 ),
    .ZN(\V3/V2/V4/V1/w4 ));
 XOR2_X2 \V3/V2/V4/V1/HA1/_1_  (.A(\V3/V2/V4/V1/w2 ),
    .B(\V3/V2/V4/V1/w1 ),
    .Z(\V3/V2/v4 [1]));
 AND2_X1 \V3/V2/V4/V1/HA2/_0_  (.A1(\V3/V2/V4/V1/w4 ),
    .A2(\V3/V2/V4/V1/w3 ),
    .ZN(\V3/V2/V4/v1 [3]));
 XOR2_X2 \V3/V2/V4/V1/HA2/_1_  (.A(\V3/V2/V4/V1/w4 ),
    .B(\V3/V2/V4/V1/w3 ),
    .Z(\V3/V2/V4/v1 [2]));
 AND2_X1 \V3/V2/V4/V1/_0_  (.A1(net45),
    .A2(net18),
    .ZN(\V3/V2/v4 [0]));
 AND2_X1 \V3/V2/V4/V1/_1_  (.A1(net45),
    .A2(net17),
    .ZN(\V3/V2/V4/V1/w1 ));
 AND2_X1 \V3/V2/V4/V1/_2_  (.A1(net18),
    .A2(net44),
    .ZN(\V3/V2/V4/V1/w2 ));
 AND2_X1 \V3/V2/V4/V1/_3_  (.A1(net17),
    .A2(net44),
    .ZN(\V3/V2/V4/V1/w3 ));
 AND2_X1 \V3/V2/V4/V2/HA1/_0_  (.A1(\V3/V2/V4/V2/w2 ),
    .A2(\V3/V2/V4/V2/w1 ),
    .ZN(\V3/V2/V4/V2/w4 ));
 XOR2_X2 \V3/V2/V4/V2/HA1/_1_  (.A(\V3/V2/V4/V2/w2 ),
    .B(\V3/V2/V4/V2/w1 ),
    .Z(\V3/V2/V4/v2 [1]));
 AND2_X1 \V3/V2/V4/V2/HA2/_0_  (.A1(\V3/V2/V4/V2/w4 ),
    .A2(\V3/V2/V4/V2/w3 ),
    .ZN(\V3/V2/V4/v2 [3]));
 XOR2_X2 \V3/V2/V4/V2/HA2/_1_  (.A(\V3/V2/V4/V2/w4 ),
    .B(\V3/V2/V4/V2/w3 ),
    .Z(\V3/V2/V4/v2 [2]));
 AND2_X1 \V3/V2/V4/V2/_0_  (.A1(net43),
    .A2(net18),
    .ZN(\V3/V2/V4/v2 [0]));
 AND2_X1 \V3/V2/V4/V2/_1_  (.A1(net43),
    .A2(net17),
    .ZN(\V3/V2/V4/V2/w1 ));
 AND2_X1 \V3/V2/V4/V2/_2_  (.A1(net18),
    .A2(net42),
    .ZN(\V3/V2/V4/V2/w2 ));
 AND2_X1 \V3/V2/V4/V2/_3_  (.A1(net17),
    .A2(net42),
    .ZN(\V3/V2/V4/V2/w3 ));
 AND2_X1 \V3/V2/V4/V3/HA1/_0_  (.A1(\V3/V2/V4/V3/w2 ),
    .A2(\V3/V2/V4/V3/w1 ),
    .ZN(\V3/V2/V4/V3/w4 ));
 XOR2_X2 \V3/V2/V4/V3/HA1/_1_  (.A(\V3/V2/V4/V3/w2 ),
    .B(\V3/V2/V4/V3/w1 ),
    .Z(\V3/V2/V4/v3 [1]));
 AND2_X1 \V3/V2/V4/V3/HA2/_0_  (.A1(\V3/V2/V4/V3/w4 ),
    .A2(\V3/V2/V4/V3/w3 ),
    .ZN(\V3/V2/V4/v3 [3]));
 XOR2_X2 \V3/V2/V4/V3/HA2/_1_  (.A(\V3/V2/V4/V3/w4 ),
    .B(\V3/V2/V4/V3/w3 ),
    .Z(\V3/V2/V4/v3 [2]));
 AND2_X1 \V3/V2/V4/V3/_0_  (.A1(net45),
    .A2(net16),
    .ZN(\V3/V2/V4/v3 [0]));
 AND2_X1 \V3/V2/V4/V3/_1_  (.A1(net45),
    .A2(net15),
    .ZN(\V3/V2/V4/V3/w1 ));
 AND2_X1 \V3/V2/V4/V3/_2_  (.A1(net16),
    .A2(net44),
    .ZN(\V3/V2/V4/V3/w2 ));
 AND2_X1 \V3/V2/V4/V3/_3_  (.A1(net15),
    .A2(net44),
    .ZN(\V3/V2/V4/V3/w3 ));
 AND2_X1 \V3/V2/V4/V4/HA1/_0_  (.A1(\V3/V2/V4/V4/w2 ),
    .A2(\V3/V2/V4/V4/w1 ),
    .ZN(\V3/V2/V4/V4/w4 ));
 XOR2_X2 \V3/V2/V4/V4/HA1/_1_  (.A(\V3/V2/V4/V4/w2 ),
    .B(\V3/V2/V4/V4/w1 ),
    .Z(\V3/V2/V4/v4 [1]));
 AND2_X1 \V3/V2/V4/V4/HA2/_0_  (.A1(\V3/V2/V4/V4/w4 ),
    .A2(\V3/V2/V4/V4/w3 ),
    .ZN(\V3/V2/V4/v4 [3]));
 XOR2_X2 \V3/V2/V4/V4/HA2/_1_  (.A(\V3/V2/V4/V4/w4 ),
    .B(\V3/V2/V4/V4/w3 ),
    .Z(\V3/V2/V4/v4 [2]));
 AND2_X1 \V3/V2/V4/V4/_0_  (.A1(net43),
    .A2(net16),
    .ZN(\V3/V2/V4/v4 [0]));
 AND2_X1 \V3/V2/V4/V4/_1_  (.A1(net43),
    .A2(net15),
    .ZN(\V3/V2/V4/V4/w1 ));
 AND2_X1 \V3/V2/V4/V4/_2_  (.A1(net16),
    .A2(net42),
    .ZN(\V3/V2/V4/V4/w2 ));
 AND2_X1 \V3/V2/V4/V4/_3_  (.A1(net15),
    .A2(net42),
    .ZN(\V3/V2/V4/V4/w3 ));
 OR2_X1 \V3/V2/V4/_0_  (.A1(\V3/V2/V4/c1 ),
    .A2(\V3/V2/V4/c2 ),
    .ZN(\V3/V2/V4/c3 ));
 OR2_X1 \V3/V2/_0_  (.A1(\V3/V2/c1 ),
    .A2(\V3/V2/c2 ),
    .ZN(\V3/V2/c3 ));
 AND2_X1 \V3/V3/A1/A1/M1/M1/_0_  (.A1(\V3/V3/v2 [0]),
    .A2(\V3/V3/v3 [0]),
    .ZN(\V3/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M1/M1/_1_  (.A(\V3/V3/v2 [0]),
    .B(\V3/V3/v3 [0]),
    .Z(\V3/V3/A1/A1/M1/s1 ));
 AND2_X1 \V3/V3/A1/A1/M1/M2/_0_  (.A1(\V3/V3/A1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M1/M2/_1_  (.A(\V3/V3/A1/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V3/s1 [0]));
 OR2_X1 \V3/V3/A1/A1/M1/_0_  (.A1(\V3/V3/A1/A1/M1/c1 ),
    .A2(\V3/V3/A1/A1/M1/c2 ),
    .ZN(\V3/V3/A1/A1/c1 ));
 AND2_X1 \V3/V3/A1/A1/M2/M1/_0_  (.A1(\V3/V3/v2 [1]),
    .A2(\V3/V3/v3 [1]),
    .ZN(\V3/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M2/M1/_1_  (.A(\V3/V3/v2 [1]),
    .B(\V3/V3/v3 [1]),
    .Z(\V3/V3/A1/A1/M2/s1 ));
 AND2_X1 \V3/V3/A1/A1/M2/M2/_0_  (.A1(\V3/V3/A1/A1/M2/s1 ),
    .A2(\V3/V3/A1/A1/c1 ),
    .ZN(\V3/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M2/M2/_1_  (.A(\V3/V3/A1/A1/M2/s1 ),
    .B(\V3/V3/A1/A1/c1 ),
    .Z(\V3/V3/s1 [1]));
 OR2_X1 \V3/V3/A1/A1/M2/_0_  (.A1(\V3/V3/A1/A1/M2/c1 ),
    .A2(\V3/V3/A1/A1/M2/c2 ),
    .ZN(\V3/V3/A1/A1/c2 ));
 AND2_X1 \V3/V3/A1/A1/M3/M1/_0_  (.A1(\V3/V3/v2 [2]),
    .A2(\V3/V3/v3 [2]),
    .ZN(\V3/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M3/M1/_1_  (.A(\V3/V3/v2 [2]),
    .B(\V3/V3/v3 [2]),
    .Z(\V3/V3/A1/A1/M3/s1 ));
 AND2_X1 \V3/V3/A1/A1/M3/M2/_0_  (.A1(\V3/V3/A1/A1/M3/s1 ),
    .A2(\V3/V3/A1/A1/c2 ),
    .ZN(\V3/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M3/M2/_1_  (.A(\V3/V3/A1/A1/M3/s1 ),
    .B(\V3/V3/A1/A1/c2 ),
    .Z(\V3/V3/s1 [2]));
 OR2_X1 \V3/V3/A1/A1/M3/_0_  (.A1(\V3/V3/A1/A1/M3/c1 ),
    .A2(\V3/V3/A1/A1/M3/c2 ),
    .ZN(\V3/V3/A1/A1/c3 ));
 AND2_X1 \V3/V3/A1/A1/M4/M1/_0_  (.A1(\V3/V3/v2 [3]),
    .A2(\V3/V3/v3 [3]),
    .ZN(\V3/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A1/A1/M4/M1/_1_  (.A(\V3/V3/v2 [3]),
    .B(\V3/V3/v3 [3]),
    .Z(\V3/V3/A1/A1/M4/s1 ));
 AND2_X1 \V3/V3/A1/A1/M4/M2/_0_  (.A1(\V3/V3/A1/A1/M4/s1 ),
    .A2(\V3/V3/A1/A1/c3 ),
    .ZN(\V3/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A1/A1/M4/M2/_1_  (.A(\V3/V3/A1/A1/M4/s1 ),
    .B(\V3/V3/A1/A1/c3 ),
    .Z(\V3/V3/s1 [3]));
 OR2_X1 \V3/V3/A1/A1/M4/_0_  (.A1(\V3/V3/A1/A1/M4/c1 ),
    .A2(\V3/V3/A1/A1/M4/c2 ),
    .ZN(\V3/V3/A1/c1 ));
 AND2_X1 \V3/V3/A1/A2/M1/M1/_0_  (.A1(\V3/V3/v2 [4]),
    .A2(\V3/V3/v3 [4]),
    .ZN(\V3/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M1/M1/_1_  (.A(\V3/V3/v2 [4]),
    .B(\V3/V3/v3 [4]),
    .Z(\V3/V3/A1/A2/M1/s1 ));
 AND2_X1 \V3/V3/A1/A2/M1/M2/_0_  (.A1(\V3/V3/A1/A2/M1/s1 ),
    .A2(\V3/V3/A1/c1 ),
    .ZN(\V3/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M1/M2/_1_  (.A(\V3/V3/A1/A2/M1/s1 ),
    .B(\V3/V3/A1/c1 ),
    .Z(\V3/V3/s1 [4]));
 OR2_X1 \V3/V3/A1/A2/M1/_0_  (.A1(\V3/V3/A1/A2/M1/c1 ),
    .A2(\V3/V3/A1/A2/M1/c2 ),
    .ZN(\V3/V3/A1/A2/c1 ));
 AND2_X1 \V3/V3/A1/A2/M2/M1/_0_  (.A1(\V3/V3/v2 [5]),
    .A2(\V3/V3/v3 [5]),
    .ZN(\V3/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M2/M1/_1_  (.A(\V3/V3/v2 [5]),
    .B(\V3/V3/v3 [5]),
    .Z(\V3/V3/A1/A2/M2/s1 ));
 AND2_X1 \V3/V3/A1/A2/M2/M2/_0_  (.A1(\V3/V3/A1/A2/M2/s1 ),
    .A2(\V3/V3/A1/A2/c1 ),
    .ZN(\V3/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M2/M2/_1_  (.A(\V3/V3/A1/A2/M2/s1 ),
    .B(\V3/V3/A1/A2/c1 ),
    .Z(\V3/V3/s1 [5]));
 OR2_X1 \V3/V3/A1/A2/M2/_0_  (.A1(\V3/V3/A1/A2/M2/c1 ),
    .A2(\V3/V3/A1/A2/M2/c2 ),
    .ZN(\V3/V3/A1/A2/c2 ));
 AND2_X1 \V3/V3/A1/A2/M3/M1/_0_  (.A1(\V3/V3/v2 [6]),
    .A2(\V3/V3/v3 [6]),
    .ZN(\V3/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M3/M1/_1_  (.A(\V3/V3/v2 [6]),
    .B(\V3/V3/v3 [6]),
    .Z(\V3/V3/A1/A2/M3/s1 ));
 AND2_X1 \V3/V3/A1/A2/M3/M2/_0_  (.A1(\V3/V3/A1/A2/M3/s1 ),
    .A2(\V3/V3/A1/A2/c2 ),
    .ZN(\V3/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M3/M2/_1_  (.A(\V3/V3/A1/A2/M3/s1 ),
    .B(\V3/V3/A1/A2/c2 ),
    .Z(\V3/V3/s1 [6]));
 OR2_X1 \V3/V3/A1/A2/M3/_0_  (.A1(\V3/V3/A1/A2/M3/c1 ),
    .A2(\V3/V3/A1/A2/M3/c2 ),
    .ZN(\V3/V3/A1/A2/c3 ));
 AND2_X1 \V3/V3/A1/A2/M4/M1/_0_  (.A1(\V3/V3/v2 [7]),
    .A2(\V3/V3/v3 [7]),
    .ZN(\V3/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A1/A2/M4/M1/_1_  (.A(\V3/V3/v2 [7]),
    .B(\V3/V3/v3 [7]),
    .Z(\V3/V3/A1/A2/M4/s1 ));
 AND2_X1 \V3/V3/A1/A2/M4/M2/_0_  (.A1(\V3/V3/A1/A2/M4/s1 ),
    .A2(\V3/V3/A1/A2/c3 ),
    .ZN(\V3/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A1/A2/M4/M2/_1_  (.A(\V3/V3/A1/A2/M4/s1 ),
    .B(\V3/V3/A1/A2/c3 ),
    .Z(\V3/V3/s1 [7]));
 OR2_X1 \V3/V3/A1/A2/M4/_0_  (.A1(\V3/V3/A1/A2/M4/c1 ),
    .A2(\V3/V3/A1/A2/M4/c2 ),
    .ZN(\V3/V3/c1 ));
 AND2_X1 \V3/V3/A2/A1/M1/M1/_0_  (.A1(\V3/V3/s1 [0]),
    .A2(\V3/V3/v1 [4]),
    .ZN(\V3/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M1/M1/_1_  (.A(\V3/V3/s1 [0]),
    .B(\V3/V3/v1 [4]),
    .Z(\V3/V3/A2/A1/M1/s1 ));
 AND2_X1 \V3/V3/A2/A1/M1/M2/_0_  (.A1(\V3/V3/A2/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M1/M2/_1_  (.A(\V3/V3/A2/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/v3 [4]));
 OR2_X1 \V3/V3/A2/A1/M1/_0_  (.A1(\V3/V3/A2/A1/M1/c1 ),
    .A2(\V3/V3/A2/A1/M1/c2 ),
    .ZN(\V3/V3/A2/A1/c1 ));
 AND2_X1 \V3/V3/A2/A1/M2/M1/_0_  (.A1(\V3/V3/s1 [1]),
    .A2(\V3/V3/v1 [5]),
    .ZN(\V3/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M2/M1/_1_  (.A(\V3/V3/s1 [1]),
    .B(\V3/V3/v1 [5]),
    .Z(\V3/V3/A2/A1/M2/s1 ));
 AND2_X1 \V3/V3/A2/A1/M2/M2/_0_  (.A1(\V3/V3/A2/A1/M2/s1 ),
    .A2(\V3/V3/A2/A1/c1 ),
    .ZN(\V3/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M2/M2/_1_  (.A(\V3/V3/A2/A1/M2/s1 ),
    .B(\V3/V3/A2/A1/c1 ),
    .Z(\V3/v3 [5]));
 OR2_X1 \V3/V3/A2/A1/M2/_0_  (.A1(\V3/V3/A2/A1/M2/c1 ),
    .A2(\V3/V3/A2/A1/M2/c2 ),
    .ZN(\V3/V3/A2/A1/c2 ));
 AND2_X1 \V3/V3/A2/A1/M3/M1/_0_  (.A1(\V3/V3/s1 [2]),
    .A2(\V3/V3/v1 [6]),
    .ZN(\V3/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M3/M1/_1_  (.A(\V3/V3/s1 [2]),
    .B(\V3/V3/v1 [6]),
    .Z(\V3/V3/A2/A1/M3/s1 ));
 AND2_X1 \V3/V3/A2/A1/M3/M2/_0_  (.A1(\V3/V3/A2/A1/M3/s1 ),
    .A2(\V3/V3/A2/A1/c2 ),
    .ZN(\V3/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M3/M2/_1_  (.A(\V3/V3/A2/A1/M3/s1 ),
    .B(\V3/V3/A2/A1/c2 ),
    .Z(\V3/v3 [6]));
 OR2_X1 \V3/V3/A2/A1/M3/_0_  (.A1(\V3/V3/A2/A1/M3/c1 ),
    .A2(\V3/V3/A2/A1/M3/c2 ),
    .ZN(\V3/V3/A2/A1/c3 ));
 AND2_X1 \V3/V3/A2/A1/M4/M1/_0_  (.A1(\V3/V3/s1 [3]),
    .A2(\V3/V3/v1 [7]),
    .ZN(\V3/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A2/A1/M4/M1/_1_  (.A(\V3/V3/s1 [3]),
    .B(\V3/V3/v1 [7]),
    .Z(\V3/V3/A2/A1/M4/s1 ));
 AND2_X1 \V3/V3/A2/A1/M4/M2/_0_  (.A1(\V3/V3/A2/A1/M4/s1 ),
    .A2(\V3/V3/A2/A1/c3 ),
    .ZN(\V3/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A2/A1/M4/M2/_1_  (.A(\V3/V3/A2/A1/M4/s1 ),
    .B(\V3/V3/A2/A1/c3 ),
    .Z(\V3/v3 [7]));
 OR2_X1 \V3/V3/A2/A1/M4/_0_  (.A1(\V3/V3/A2/A1/M4/c1 ),
    .A2(\V3/V3/A2/A1/M4/c2 ),
    .ZN(\V3/V3/A2/c1 ));
 AND2_X1 \V3/V3/A2/A2/M1/M1/_0_  (.A1(\V3/V3/s1 [4]),
    .A2(net8),
    .ZN(\V3/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M1/M1/_1_  (.A(\V3/V3/s1 [4]),
    .B(net8),
    .Z(\V3/V3/A2/A2/M1/s1 ));
 AND2_X1 \V3/V3/A2/A2/M1/M2/_0_  (.A1(\V3/V3/A2/A2/M1/s1 ),
    .A2(\V3/V3/A2/c1 ),
    .ZN(\V3/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M1/M2/_1_  (.A(\V3/V3/A2/A2/M1/s1 ),
    .B(\V3/V3/A2/c1 ),
    .Z(\V3/V3/s2 [4]));
 OR2_X1 \V3/V3/A2/A2/M1/_0_  (.A1(\V3/V3/A2/A2/M1/c1 ),
    .A2(\V3/V3/A2/A2/M1/c2 ),
    .ZN(\V3/V3/A2/A2/c1 ));
 AND2_X1 \V3/V3/A2/A2/M2/M1/_0_  (.A1(\V3/V3/s1 [5]),
    .A2(net8),
    .ZN(\V3/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M2/M1/_1_  (.A(\V3/V3/s1 [5]),
    .B(net8),
    .Z(\V3/V3/A2/A2/M2/s1 ));
 AND2_X1 \V3/V3/A2/A2/M2/M2/_0_  (.A1(\V3/V3/A2/A2/M2/s1 ),
    .A2(\V3/V3/A2/A2/c1 ),
    .ZN(\V3/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M2/M2/_1_  (.A(\V3/V3/A2/A2/M2/s1 ),
    .B(\V3/V3/A2/A2/c1 ),
    .Z(\V3/V3/s2 [5]));
 OR2_X1 \V3/V3/A2/A2/M2/_0_  (.A1(\V3/V3/A2/A2/M2/c1 ),
    .A2(\V3/V3/A2/A2/M2/c2 ),
    .ZN(\V3/V3/A2/A2/c2 ));
 AND2_X1 \V3/V3/A2/A2/M3/M1/_0_  (.A1(\V3/V3/s1 [6]),
    .A2(net8),
    .ZN(\V3/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M3/M1/_1_  (.A(\V3/V3/s1 [6]),
    .B(net8),
    .Z(\V3/V3/A2/A2/M3/s1 ));
 AND2_X1 \V3/V3/A2/A2/M3/M2/_0_  (.A1(\V3/V3/A2/A2/M3/s1 ),
    .A2(\V3/V3/A2/A2/c2 ),
    .ZN(\V3/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M3/M2/_1_  (.A(\V3/V3/A2/A2/M3/s1 ),
    .B(\V3/V3/A2/A2/c2 ),
    .Z(\V3/V3/s2 [6]));
 OR2_X1 \V3/V3/A2/A2/M3/_0_  (.A1(\V3/V3/A2/A2/M3/c1 ),
    .A2(\V3/V3/A2/A2/M3/c2 ),
    .ZN(\V3/V3/A2/A2/c3 ));
 AND2_X1 \V3/V3/A2/A2/M4/M1/_0_  (.A1(\V3/V3/s1 [7]),
    .A2(net8),
    .ZN(\V3/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A2/A2/M4/M1/_1_  (.A(\V3/V3/s1 [7]),
    .B(net8),
    .Z(\V3/V3/A2/A2/M4/s1 ));
 AND2_X1 \V3/V3/A2/A2/M4/M2/_0_  (.A1(\V3/V3/A2/A2/M4/s1 ),
    .A2(\V3/V3/A2/A2/c3 ),
    .ZN(\V3/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A2/A2/M4/M2/_1_  (.A(\V3/V3/A2/A2/M4/s1 ),
    .B(\V3/V3/A2/A2/c3 ),
    .Z(\V3/V3/s2 [7]));
 OR2_X1 \V3/V3/A2/A2/M4/_0_  (.A1(\V3/V3/A2/A2/M4/c1 ),
    .A2(\V3/V3/A2/A2/M4/c2 ),
    .ZN(\V3/V3/c2 ));
 AND2_X1 \V3/V3/A3/A1/M1/M1/_0_  (.A1(\V3/V3/v4 [0]),
    .A2(\V3/V3/s2 [4]),
    .ZN(\V3/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M1/M1/_1_  (.A(\V3/V3/v4 [0]),
    .B(\V3/V3/s2 [4]),
    .Z(\V3/V3/A3/A1/M1/s1 ));
 AND2_X1 \V3/V3/A3/A1/M1/M2/_0_  (.A1(\V3/V3/A3/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M1/M2/_1_  (.A(\V3/V3/A3/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/v3 [8]));
 OR2_X1 \V3/V3/A3/A1/M1/_0_  (.A1(\V3/V3/A3/A1/M1/c1 ),
    .A2(\V3/V3/A3/A1/M1/c2 ),
    .ZN(\V3/V3/A3/A1/c1 ));
 AND2_X1 \V3/V3/A3/A1/M2/M1/_0_  (.A1(\V3/V3/v4 [1]),
    .A2(\V3/V3/s2 [5]),
    .ZN(\V3/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M2/M1/_1_  (.A(\V3/V3/v4 [1]),
    .B(\V3/V3/s2 [5]),
    .Z(\V3/V3/A3/A1/M2/s1 ));
 AND2_X1 \V3/V3/A3/A1/M2/M2/_0_  (.A1(\V3/V3/A3/A1/M2/s1 ),
    .A2(\V3/V3/A3/A1/c1 ),
    .ZN(\V3/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M2/M2/_1_  (.A(\V3/V3/A3/A1/M2/s1 ),
    .B(\V3/V3/A3/A1/c1 ),
    .Z(\V3/v3 [9]));
 OR2_X1 \V3/V3/A3/A1/M2/_0_  (.A1(\V3/V3/A3/A1/M2/c1 ),
    .A2(\V3/V3/A3/A1/M2/c2 ),
    .ZN(\V3/V3/A3/A1/c2 ));
 AND2_X1 \V3/V3/A3/A1/M3/M1/_0_  (.A1(\V3/V3/v4 [2]),
    .A2(\V3/V3/s2 [6]),
    .ZN(\V3/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M3/M1/_1_  (.A(\V3/V3/v4 [2]),
    .B(\V3/V3/s2 [6]),
    .Z(\V3/V3/A3/A1/M3/s1 ));
 AND2_X1 \V3/V3/A3/A1/M3/M2/_0_  (.A1(\V3/V3/A3/A1/M3/s1 ),
    .A2(\V3/V3/A3/A1/c2 ),
    .ZN(\V3/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M3/M2/_1_  (.A(\V3/V3/A3/A1/M3/s1 ),
    .B(\V3/V3/A3/A1/c2 ),
    .Z(\V3/v3 [10]));
 OR2_X1 \V3/V3/A3/A1/M3/_0_  (.A1(\V3/V3/A3/A1/M3/c1 ),
    .A2(\V3/V3/A3/A1/M3/c2 ),
    .ZN(\V3/V3/A3/A1/c3 ));
 AND2_X1 \V3/V3/A3/A1/M4/M1/_0_  (.A1(\V3/V3/v4 [3]),
    .A2(\V3/V3/s2 [7]),
    .ZN(\V3/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V3/A3/A1/M4/M1/_1_  (.A(\V3/V3/v4 [3]),
    .B(\V3/V3/s2 [7]),
    .Z(\V3/V3/A3/A1/M4/s1 ));
 AND2_X1 \V3/V3/A3/A1/M4/M2/_0_  (.A1(\V3/V3/A3/A1/M4/s1 ),
    .A2(\V3/V3/A3/A1/c3 ),
    .ZN(\V3/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V3/A3/A1/M4/M2/_1_  (.A(\V3/V3/A3/A1/M4/s1 ),
    .B(\V3/V3/A3/A1/c3 ),
    .Z(\V3/v3 [11]));
 OR2_X1 \V3/V3/A3/A1/M4/_0_  (.A1(\V3/V3/A3/A1/M4/c1 ),
    .A2(\V3/V3/A3/A1/M4/c2 ),
    .ZN(\V3/V3/A3/c1 ));
 AND2_X1 \V3/V3/A3/A2/M1/M1/_0_  (.A1(\V3/V3/v4 [4]),
    .A2(\V3/V3/c3 ),
    .ZN(\V3/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M1/M1/_1_  (.A(\V3/V3/v4 [4]),
    .B(\V3/V3/c3 ),
    .Z(\V3/V3/A3/A2/M1/s1 ));
 AND2_X1 \V3/V3/A3/A2/M1/M2/_0_  (.A1(\V3/V3/A3/A2/M1/s1 ),
    .A2(\V3/V3/A3/c1 ),
    .ZN(\V3/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M1/M2/_1_  (.A(\V3/V3/A3/A2/M1/s1 ),
    .B(\V3/V3/A3/c1 ),
    .Z(\V3/v3 [12]));
 OR2_X1 \V3/V3/A3/A2/M1/_0_  (.A1(\V3/V3/A3/A2/M1/c1 ),
    .A2(\V3/V3/A3/A2/M1/c2 ),
    .ZN(\V3/V3/A3/A2/c1 ));
 AND2_X1 \V3/V3/A3/A2/M2/M1/_0_  (.A1(\V3/V3/v4 [5]),
    .A2(net8),
    .ZN(\V3/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M2/M1/_1_  (.A(\V3/V3/v4 [5]),
    .B(net8),
    .Z(\V3/V3/A3/A2/M2/s1 ));
 AND2_X1 \V3/V3/A3/A2/M2/M2/_0_  (.A1(\V3/V3/A3/A2/M2/s1 ),
    .A2(\V3/V3/A3/A2/c1 ),
    .ZN(\V3/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M2/M2/_1_  (.A(\V3/V3/A3/A2/M2/s1 ),
    .B(\V3/V3/A3/A2/c1 ),
    .Z(\V3/v3 [13]));
 OR2_X1 \V3/V3/A3/A2/M2/_0_  (.A1(\V3/V3/A3/A2/M2/c1 ),
    .A2(\V3/V3/A3/A2/M2/c2 ),
    .ZN(\V3/V3/A3/A2/c2 ));
 AND2_X1 \V3/V3/A3/A2/M3/M1/_0_  (.A1(\V3/V3/v4 [6]),
    .A2(net8),
    .ZN(\V3/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M3/M1/_1_  (.A(\V3/V3/v4 [6]),
    .B(net8),
    .Z(\V3/V3/A3/A2/M3/s1 ));
 AND2_X1 \V3/V3/A3/A2/M3/M2/_0_  (.A1(\V3/V3/A3/A2/M3/s1 ),
    .A2(\V3/V3/A3/A2/c2 ),
    .ZN(\V3/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M3/M2/_1_  (.A(\V3/V3/A3/A2/M3/s1 ),
    .B(\V3/V3/A3/A2/c2 ),
    .Z(\V3/v3 [14]));
 OR2_X1 \V3/V3/A3/A2/M3/_0_  (.A1(\V3/V3/A3/A2/M3/c1 ),
    .A2(\V3/V3/A3/A2/M3/c2 ),
    .ZN(\V3/V3/A3/A2/c3 ));
 AND2_X1 \V3/V3/A3/A2/M4/M1/_0_  (.A1(\V3/V3/v4 [7]),
    .A2(net8),
    .ZN(\V3/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V3/A3/A2/M4/M1/_1_  (.A(\V3/V3/v4 [7]),
    .B(net8),
    .Z(\V3/V3/A3/A2/M4/s1 ));
 AND2_X1 \V3/V3/A3/A2/M4/M2/_0_  (.A1(\V3/V3/A3/A2/M4/s1 ),
    .A2(\V3/V3/A3/A2/c3 ),
    .ZN(\V3/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V3/A3/A2/M4/M2/_1_  (.A(\V3/V3/A3/A2/M4/s1 ),
    .B(\V3/V3/A3/A2/c3 ),
    .Z(\V3/v3 [15]));
 OR2_X1 \V3/V3/A3/A2/M4/_0_  (.A1(\V3/V3/A3/A2/M4/c1 ),
    .A2(\V3/V3/A3/A2/M4/c2 ),
    .ZN(\V3/V3/overflow ));
 AND2_X1 \V3/V3/V1/A1/M1/M1/_0_  (.A1(\V3/V3/V1/v2 [0]),
    .A2(\V3/V3/V1/v3 [0]),
    .ZN(\V3/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M1/M1/_1_  (.A(\V3/V3/V1/v2 [0]),
    .B(\V3/V3/V1/v3 [0]),
    .Z(\V3/V3/V1/A1/M1/s1 ));
 AND2_X1 \V3/V3/V1/A1/M1/M2/_0_  (.A1(\V3/V3/V1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M1/M2/_1_  (.A(\V3/V3/V1/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V3/V1/s1 [0]));
 OR2_X1 \V3/V3/V1/A1/M1/_0_  (.A1(\V3/V3/V1/A1/M1/c1 ),
    .A2(\V3/V3/V1/A1/M1/c2 ),
    .ZN(\V3/V3/V1/A1/c1 ));
 AND2_X1 \V3/V3/V1/A1/M2/M1/_0_  (.A1(\V3/V3/V1/v2 [1]),
    .A2(\V3/V3/V1/v3 [1]),
    .ZN(\V3/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M2/M1/_1_  (.A(\V3/V3/V1/v2 [1]),
    .B(\V3/V3/V1/v3 [1]),
    .Z(\V3/V3/V1/A1/M2/s1 ));
 AND2_X1 \V3/V3/V1/A1/M2/M2/_0_  (.A1(\V3/V3/V1/A1/M2/s1 ),
    .A2(\V3/V3/V1/A1/c1 ),
    .ZN(\V3/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M2/M2/_1_  (.A(\V3/V3/V1/A1/M2/s1 ),
    .B(\V3/V3/V1/A1/c1 ),
    .Z(\V3/V3/V1/s1 [1]));
 OR2_X1 \V3/V3/V1/A1/M2/_0_  (.A1(\V3/V3/V1/A1/M2/c1 ),
    .A2(\V3/V3/V1/A1/M2/c2 ),
    .ZN(\V3/V3/V1/A1/c2 ));
 AND2_X1 \V3/V3/V1/A1/M3/M1/_0_  (.A1(\V3/V3/V1/v2 [2]),
    .A2(\V3/V3/V1/v3 [2]),
    .ZN(\V3/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M3/M1/_1_  (.A(\V3/V3/V1/v2 [2]),
    .B(\V3/V3/V1/v3 [2]),
    .Z(\V3/V3/V1/A1/M3/s1 ));
 AND2_X1 \V3/V3/V1/A1/M3/M2/_0_  (.A1(\V3/V3/V1/A1/M3/s1 ),
    .A2(\V3/V3/V1/A1/c2 ),
    .ZN(\V3/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M3/M2/_1_  (.A(\V3/V3/V1/A1/M3/s1 ),
    .B(\V3/V3/V1/A1/c2 ),
    .Z(\V3/V3/V1/s1 [2]));
 OR2_X1 \V3/V3/V1/A1/M3/_0_  (.A1(\V3/V3/V1/A1/M3/c1 ),
    .A2(\V3/V3/V1/A1/M3/c2 ),
    .ZN(\V3/V3/V1/A1/c3 ));
 AND2_X1 \V3/V3/V1/A1/M4/M1/_0_  (.A1(\V3/V3/V1/v2 [3]),
    .A2(\V3/V3/V1/v3 [3]),
    .ZN(\V3/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A1/M4/M1/_1_  (.A(\V3/V3/V1/v2 [3]),
    .B(\V3/V3/V1/v3 [3]),
    .Z(\V3/V3/V1/A1/M4/s1 ));
 AND2_X1 \V3/V3/V1/A1/M4/M2/_0_  (.A1(\V3/V3/V1/A1/M4/s1 ),
    .A2(\V3/V3/V1/A1/c3 ),
    .ZN(\V3/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A1/M4/M2/_1_  (.A(\V3/V3/V1/A1/M4/s1 ),
    .B(\V3/V3/V1/A1/c3 ),
    .Z(\V3/V3/V1/s1 [3]));
 OR2_X1 \V3/V3/V1/A1/M4/_0_  (.A1(\V3/V3/V1/A1/M4/c1 ),
    .A2(\V3/V3/V1/A1/M4/c2 ),
    .ZN(\V3/V3/V1/c1 ));
 AND2_X1 \V3/V3/V1/A2/M1/M1/_0_  (.A1(\V3/V3/V1/s1 [0]),
    .A2(\V3/V3/V1/v1 [2]),
    .ZN(\V3/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M1/M1/_1_  (.A(\V3/V3/V1/s1 [0]),
    .B(\V3/V3/V1/v1 [2]),
    .Z(\V3/V3/V1/A2/M1/s1 ));
 AND2_X1 \V3/V3/V1/A2/M1/M2/_0_  (.A1(\V3/V3/V1/A2/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M1/M2/_1_  (.A(\V3/V3/V1/A2/M1/s1 ),
    .B(net5),
    .Z(\V3/v3 [2]));
 OR2_X1 \V3/V3/V1/A2/M1/_0_  (.A1(\V3/V3/V1/A2/M1/c1 ),
    .A2(\V3/V3/V1/A2/M1/c2 ),
    .ZN(\V3/V3/V1/A2/c1 ));
 AND2_X1 \V3/V3/V1/A2/M2/M1/_0_  (.A1(\V3/V3/V1/s1 [1]),
    .A2(\V3/V3/V1/v1 [3]),
    .ZN(\V3/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M2/M1/_1_  (.A(\V3/V3/V1/s1 [1]),
    .B(\V3/V3/V1/v1 [3]),
    .Z(\V3/V3/V1/A2/M2/s1 ));
 AND2_X1 \V3/V3/V1/A2/M2/M2/_0_  (.A1(\V3/V3/V1/A2/M2/s1 ),
    .A2(\V3/V3/V1/A2/c1 ),
    .ZN(\V3/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M2/M2/_1_  (.A(\V3/V3/V1/A2/M2/s1 ),
    .B(\V3/V3/V1/A2/c1 ),
    .Z(\V3/v3 [3]));
 OR2_X1 \V3/V3/V1/A2/M2/_0_  (.A1(\V3/V3/V1/A2/M2/c1 ),
    .A2(\V3/V3/V1/A2/M2/c2 ),
    .ZN(\V3/V3/V1/A2/c2 ));
 AND2_X1 \V3/V3/V1/A2/M3/M1/_0_  (.A1(\V3/V3/V1/s1 [2]),
    .A2(net5),
    .ZN(\V3/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M3/M1/_1_  (.A(\V3/V3/V1/s1 [2]),
    .B(net5),
    .Z(\V3/V3/V1/A2/M3/s1 ));
 AND2_X1 \V3/V3/V1/A2/M3/M2/_0_  (.A1(\V3/V3/V1/A2/M3/s1 ),
    .A2(\V3/V3/V1/A2/c2 ),
    .ZN(\V3/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M3/M2/_1_  (.A(\V3/V3/V1/A2/M3/s1 ),
    .B(\V3/V3/V1/A2/c2 ),
    .Z(\V3/V3/V1/s2 [2]));
 OR2_X1 \V3/V3/V1/A2/M3/_0_  (.A1(\V3/V3/V1/A2/M3/c1 ),
    .A2(\V3/V3/V1/A2/M3/c2 ),
    .ZN(\V3/V3/V1/A2/c3 ));
 AND2_X1 \V3/V3/V1/A2/M4/M1/_0_  (.A1(\V3/V3/V1/s1 [3]),
    .A2(net5),
    .ZN(\V3/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A2/M4/M1/_1_  (.A(\V3/V3/V1/s1 [3]),
    .B(net5),
    .Z(\V3/V3/V1/A2/M4/s1 ));
 AND2_X1 \V3/V3/V1/A2/M4/M2/_0_  (.A1(\V3/V3/V1/A2/M4/s1 ),
    .A2(\V3/V3/V1/A2/c3 ),
    .ZN(\V3/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A2/M4/M2/_1_  (.A(\V3/V3/V1/A2/M4/s1 ),
    .B(\V3/V3/V1/A2/c3 ),
    .Z(\V3/V3/V1/s2 [3]));
 OR2_X1 \V3/V3/V1/A2/M4/_0_  (.A1(\V3/V3/V1/A2/M4/c1 ),
    .A2(\V3/V3/V1/A2/M4/c2 ),
    .ZN(\V3/V3/V1/c2 ));
 AND2_X1 \V3/V3/V1/A3/M1/M1/_0_  (.A1(\V3/V3/V1/v4 [0]),
    .A2(\V3/V3/V1/s2 [2]),
    .ZN(\V3/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M1/M1/_1_  (.A(\V3/V3/V1/v4 [0]),
    .B(\V3/V3/V1/s2 [2]),
    .Z(\V3/V3/V1/A3/M1/s1 ));
 AND2_X1 \V3/V3/V1/A3/M1/M2/_0_  (.A1(\V3/V3/V1/A3/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M1/M2/_1_  (.A(\V3/V3/V1/A3/M1/s1 ),
    .B(net5),
    .Z(\V3/V3/v1 [4]));
 OR2_X1 \V3/V3/V1/A3/M1/_0_  (.A1(\V3/V3/V1/A3/M1/c1 ),
    .A2(\V3/V3/V1/A3/M1/c2 ),
    .ZN(\V3/V3/V1/A3/c1 ));
 AND2_X1 \V3/V3/V1/A3/M2/M1/_0_  (.A1(\V3/V3/V1/v4 [1]),
    .A2(\V3/V3/V1/s2 [3]),
    .ZN(\V3/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M2/M1/_1_  (.A(\V3/V3/V1/v4 [1]),
    .B(\V3/V3/V1/s2 [3]),
    .Z(\V3/V3/V1/A3/M2/s1 ));
 AND2_X1 \V3/V3/V1/A3/M2/M2/_0_  (.A1(\V3/V3/V1/A3/M2/s1 ),
    .A2(\V3/V3/V1/A3/c1 ),
    .ZN(\V3/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M2/M2/_1_  (.A(\V3/V3/V1/A3/M2/s1 ),
    .B(\V3/V3/V1/A3/c1 ),
    .Z(\V3/V3/v1 [5]));
 OR2_X1 \V3/V3/V1/A3/M2/_0_  (.A1(\V3/V3/V1/A3/M2/c1 ),
    .A2(\V3/V3/V1/A3/M2/c2 ),
    .ZN(\V3/V3/V1/A3/c2 ));
 AND2_X1 \V3/V3/V1/A3/M3/M1/_0_  (.A1(\V3/V3/V1/v4 [2]),
    .A2(\V3/V3/V1/c3 ),
    .ZN(\V3/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M3/M1/_1_  (.A(\V3/V3/V1/v4 [2]),
    .B(\V3/V3/V1/c3 ),
    .Z(\V3/V3/V1/A3/M3/s1 ));
 AND2_X1 \V3/V3/V1/A3/M3/M2/_0_  (.A1(\V3/V3/V1/A3/M3/s1 ),
    .A2(\V3/V3/V1/A3/c2 ),
    .ZN(\V3/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M3/M2/_1_  (.A(\V3/V3/V1/A3/M3/s1 ),
    .B(\V3/V3/V1/A3/c2 ),
    .Z(\V3/V3/v1 [6]));
 OR2_X1 \V3/V3/V1/A3/M3/_0_  (.A1(\V3/V3/V1/A3/M3/c1 ),
    .A2(\V3/V3/V1/A3/M3/c2 ),
    .ZN(\V3/V3/V1/A3/c3 ));
 AND2_X1 \V3/V3/V1/A3/M4/M1/_0_  (.A1(\V3/V3/V1/v4 [3]),
    .A2(net8),
    .ZN(\V3/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V1/A3/M4/M1/_1_  (.A(\V3/V3/V1/v4 [3]),
    .B(net8),
    .Z(\V3/V3/V1/A3/M4/s1 ));
 AND2_X1 \V3/V3/V1/A3/M4/M2/_0_  (.A1(\V3/V3/V1/A3/M4/s1 ),
    .A2(\V3/V3/V1/A3/c3 ),
    .ZN(\V3/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V1/A3/M4/M2/_1_  (.A(\V3/V3/V1/A3/M4/s1 ),
    .B(\V3/V3/V1/A3/c3 ),
    .Z(\V3/V3/v1 [7]));
 OR2_X1 \V3/V3/V1/A3/M4/_0_  (.A1(\V3/V3/V1/A3/M4/c1 ),
    .A2(\V3/V3/V1/A3/M4/c2 ),
    .ZN(\V3/V3/V1/overflow ));
 AND2_X1 \V3/V3/V1/V1/HA1/_0_  (.A1(\V3/V3/V1/V1/w2 ),
    .A2(\V3/V3/V1/V1/w1 ),
    .ZN(\V3/V3/V1/V1/w4 ));
 XOR2_X2 \V3/V3/V1/V1/HA1/_1_  (.A(\V3/V3/V1/V1/w2 ),
    .B(\V3/V3/V1/V1/w1 ),
    .Z(\V3/v3 [1]));
 AND2_X1 \V3/V3/V1/V1/HA2/_0_  (.A1(\V3/V3/V1/V1/w4 ),
    .A2(\V3/V3/V1/V1/w3 ),
    .ZN(\V3/V3/V1/v1 [3]));
 XOR2_X2 \V3/V3/V1/V1/HA2/_1_  (.A(\V3/V3/V1/V1/w4 ),
    .B(\V3/V3/V1/V1/w3 ),
    .Z(\V3/V3/V1/v1 [2]));
 AND2_X1 \V3/V3/V1/V1/_0_  (.A1(net48),
    .A2(net14),
    .ZN(\V3/v3 [0]));
 AND2_X1 \V3/V3/V1/V1/_1_  (.A1(net48),
    .A2(B[25]),
    .ZN(\V3/V3/V1/V1/w1 ));
 AND2_X1 \V3/V3/V1/V1/_2_  (.A1(net14),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V1/w2 ));
 AND2_X1 \V3/V3/V1/V1/_3_  (.A1(B[25]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V1/w3 ));
 AND2_X1 \V3/V3/V1/V2/HA1/_0_  (.A1(\V3/V3/V1/V2/w2 ),
    .A2(\V3/V3/V1/V2/w1 ),
    .ZN(\V3/V3/V1/V2/w4 ));
 XOR2_X2 \V3/V3/V1/V2/HA1/_1_  (.A(\V3/V3/V1/V2/w2 ),
    .B(\V3/V3/V1/V2/w1 ),
    .Z(\V3/V3/V1/v2 [1]));
 AND2_X1 \V3/V3/V1/V2/HA2/_0_  (.A1(\V3/V3/V1/V2/w4 ),
    .A2(\V3/V3/V1/V2/w3 ),
    .ZN(\V3/V3/V1/v2 [3]));
 XOR2_X2 \V3/V3/V1/V2/HA2/_1_  (.A(\V3/V3/V1/V2/w4 ),
    .B(\V3/V3/V1/V2/w3 ),
    .Z(\V3/V3/V1/v2 [2]));
 AND2_X1 \V3/V3/V1/V2/_0_  (.A1(A[2]),
    .A2(net14),
    .ZN(\V3/V3/V1/v2 [0]));
 AND2_X1 \V3/V3/V1/V2/_1_  (.A1(A[2]),
    .A2(B[25]),
    .ZN(\V3/V3/V1/V2/w1 ));
 AND2_X1 \V3/V3/V1/V2/_2_  (.A1(net14),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V2/w2 ));
 AND2_X1 \V3/V3/V1/V2/_3_  (.A1(B[25]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V2/w3 ));
 AND2_X1 \V3/V3/V1/V3/HA1/_0_  (.A1(\V3/V3/V1/V3/w2 ),
    .A2(\V3/V3/V1/V3/w1 ),
    .ZN(\V3/V3/V1/V3/w4 ));
 XOR2_X2 \V3/V3/V1/V3/HA1/_1_  (.A(\V3/V3/V1/V3/w2 ),
    .B(\V3/V3/V1/V3/w1 ),
    .Z(\V3/V3/V1/v3 [1]));
 AND2_X1 \V3/V3/V1/V3/HA2/_0_  (.A1(\V3/V3/V1/V3/w4 ),
    .A2(\V3/V3/V1/V3/w3 ),
    .ZN(\V3/V3/V1/v3 [3]));
 XOR2_X2 \V3/V3/V1/V3/HA2/_1_  (.A(\V3/V3/V1/V3/w4 ),
    .B(\V3/V3/V1/V3/w3 ),
    .Z(\V3/V3/V1/v3 [2]));
 AND2_X1 \V3/V3/V1/V3/_0_  (.A1(net48),
    .A2(net13),
    .ZN(\V3/V3/V1/v3 [0]));
 AND2_X1 \V3/V3/V1/V3/_1_  (.A1(net48),
    .A2(B[27]),
    .ZN(\V3/V3/V1/V3/w1 ));
 AND2_X1 \V3/V3/V1/V3/_2_  (.A1(net13),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V3/w2 ));
 AND2_X1 \V3/V3/V1/V3/_3_  (.A1(B[27]),
    .A2(A[1]),
    .ZN(\V3/V3/V1/V3/w3 ));
 AND2_X1 \V3/V3/V1/V4/HA1/_0_  (.A1(\V3/V3/V1/V4/w2 ),
    .A2(\V3/V3/V1/V4/w1 ),
    .ZN(\V3/V3/V1/V4/w4 ));
 XOR2_X2 \V3/V3/V1/V4/HA1/_1_  (.A(\V3/V3/V1/V4/w2 ),
    .B(\V3/V3/V1/V4/w1 ),
    .Z(\V3/V3/V1/v4 [1]));
 AND2_X1 \V3/V3/V1/V4/HA2/_0_  (.A1(\V3/V3/V1/V4/w4 ),
    .A2(\V3/V3/V1/V4/w3 ),
    .ZN(\V3/V3/V1/v4 [3]));
 XOR2_X2 \V3/V3/V1/V4/HA2/_1_  (.A(\V3/V3/V1/V4/w4 ),
    .B(\V3/V3/V1/V4/w3 ),
    .Z(\V3/V3/V1/v4 [2]));
 AND2_X1 \V3/V3/V1/V4/_0_  (.A1(A[2]),
    .A2(net13),
    .ZN(\V3/V3/V1/v4 [0]));
 AND2_X1 \V3/V3/V1/V4/_1_  (.A1(A[2]),
    .A2(B[27]),
    .ZN(\V3/V3/V1/V4/w1 ));
 AND2_X1 \V3/V3/V1/V4/_2_  (.A1(net13),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V4/w2 ));
 AND2_X1 \V3/V3/V1/V4/_3_  (.A1(B[27]),
    .A2(A[3]),
    .ZN(\V3/V3/V1/V4/w3 ));
 OR2_X1 \V3/V3/V1/_0_  (.A1(\V3/V3/V1/c1 ),
    .A2(\V3/V3/V1/c2 ),
    .ZN(\V3/V3/V1/c3 ));
 AND2_X1 \V3/V3/V2/A1/M1/M1/_0_  (.A1(\V3/V3/V2/v2 [0]),
    .A2(\V3/V3/V2/v3 [0]),
    .ZN(\V3/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M1/M1/_1_  (.A(\V3/V3/V2/v2 [0]),
    .B(\V3/V3/V2/v3 [0]),
    .Z(\V3/V3/V2/A1/M1/s1 ));
 AND2_X1 \V3/V3/V2/A1/M1/M2/_0_  (.A1(\V3/V3/V2/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M1/M2/_1_  (.A(\V3/V3/V2/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/V2/s1 [0]));
 OR2_X1 \V3/V3/V2/A1/M1/_0_  (.A1(\V3/V3/V2/A1/M1/c1 ),
    .A2(\V3/V3/V2/A1/M1/c2 ),
    .ZN(\V3/V3/V2/A1/c1 ));
 AND2_X1 \V3/V3/V2/A1/M2/M1/_0_  (.A1(\V3/V3/V2/v2 [1]),
    .A2(\V3/V3/V2/v3 [1]),
    .ZN(\V3/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M2/M1/_1_  (.A(\V3/V3/V2/v2 [1]),
    .B(\V3/V3/V2/v3 [1]),
    .Z(\V3/V3/V2/A1/M2/s1 ));
 AND2_X1 \V3/V3/V2/A1/M2/M2/_0_  (.A1(\V3/V3/V2/A1/M2/s1 ),
    .A2(\V3/V3/V2/A1/c1 ),
    .ZN(\V3/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M2/M2/_1_  (.A(\V3/V3/V2/A1/M2/s1 ),
    .B(\V3/V3/V2/A1/c1 ),
    .Z(\V3/V3/V2/s1 [1]));
 OR2_X1 \V3/V3/V2/A1/M2/_0_  (.A1(\V3/V3/V2/A1/M2/c1 ),
    .A2(\V3/V3/V2/A1/M2/c2 ),
    .ZN(\V3/V3/V2/A1/c2 ));
 AND2_X1 \V3/V3/V2/A1/M3/M1/_0_  (.A1(\V3/V3/V2/v2 [2]),
    .A2(\V3/V3/V2/v3 [2]),
    .ZN(\V3/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M3/M1/_1_  (.A(\V3/V3/V2/v2 [2]),
    .B(\V3/V3/V2/v3 [2]),
    .Z(\V3/V3/V2/A1/M3/s1 ));
 AND2_X1 \V3/V3/V2/A1/M3/M2/_0_  (.A1(\V3/V3/V2/A1/M3/s1 ),
    .A2(\V3/V3/V2/A1/c2 ),
    .ZN(\V3/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M3/M2/_1_  (.A(\V3/V3/V2/A1/M3/s1 ),
    .B(\V3/V3/V2/A1/c2 ),
    .Z(\V3/V3/V2/s1 [2]));
 OR2_X1 \V3/V3/V2/A1/M3/_0_  (.A1(\V3/V3/V2/A1/M3/c1 ),
    .A2(\V3/V3/V2/A1/M3/c2 ),
    .ZN(\V3/V3/V2/A1/c3 ));
 AND2_X1 \V3/V3/V2/A1/M4/M1/_0_  (.A1(\V3/V3/V2/v2 [3]),
    .A2(\V3/V3/V2/v3 [3]),
    .ZN(\V3/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A1/M4/M1/_1_  (.A(\V3/V3/V2/v2 [3]),
    .B(\V3/V3/V2/v3 [3]),
    .Z(\V3/V3/V2/A1/M4/s1 ));
 AND2_X1 \V3/V3/V2/A1/M4/M2/_0_  (.A1(\V3/V3/V2/A1/M4/s1 ),
    .A2(\V3/V3/V2/A1/c3 ),
    .ZN(\V3/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A1/M4/M2/_1_  (.A(\V3/V3/V2/A1/M4/s1 ),
    .B(\V3/V3/V2/A1/c3 ),
    .Z(\V3/V3/V2/s1 [3]));
 OR2_X1 \V3/V3/V2/A1/M4/_0_  (.A1(\V3/V3/V2/A1/M4/c1 ),
    .A2(\V3/V3/V2/A1/M4/c2 ),
    .ZN(\V3/V3/V2/c1 ));
 AND2_X1 \V3/V3/V2/A2/M1/M1/_0_  (.A1(\V3/V3/V2/s1 [0]),
    .A2(\V3/V3/V2/v1 [2]),
    .ZN(\V3/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M1/M1/_1_  (.A(\V3/V3/V2/s1 [0]),
    .B(\V3/V3/V2/v1 [2]),
    .Z(\V3/V3/V2/A2/M1/s1 ));
 AND2_X1 \V3/V3/V2/A2/M1/M2/_0_  (.A1(\V3/V3/V2/A2/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M1/M2/_1_  (.A(\V3/V3/V2/A2/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v2 [2]));
 OR2_X1 \V3/V3/V2/A2/M1/_0_  (.A1(\V3/V3/V2/A2/M1/c1 ),
    .A2(\V3/V3/V2/A2/M1/c2 ),
    .ZN(\V3/V3/V2/A2/c1 ));
 AND2_X1 \V3/V3/V2/A2/M2/M1/_0_  (.A1(\V3/V3/V2/s1 [1]),
    .A2(\V3/V3/V2/v1 [3]),
    .ZN(\V3/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M2/M1/_1_  (.A(\V3/V3/V2/s1 [1]),
    .B(\V3/V3/V2/v1 [3]),
    .Z(\V3/V3/V2/A2/M2/s1 ));
 AND2_X1 \V3/V3/V2/A2/M2/M2/_0_  (.A1(\V3/V3/V2/A2/M2/s1 ),
    .A2(\V3/V3/V2/A2/c1 ),
    .ZN(\V3/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M2/M2/_1_  (.A(\V3/V3/V2/A2/M2/s1 ),
    .B(\V3/V3/V2/A2/c1 ),
    .Z(\V3/V3/v2 [3]));
 OR2_X1 \V3/V3/V2/A2/M2/_0_  (.A1(\V3/V3/V2/A2/M2/c1 ),
    .A2(\V3/V3/V2/A2/M2/c2 ),
    .ZN(\V3/V3/V2/A2/c2 ));
 AND2_X1 \V3/V3/V2/A2/M3/M1/_0_  (.A1(\V3/V3/V2/s1 [2]),
    .A2(net8),
    .ZN(\V3/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M3/M1/_1_  (.A(\V3/V3/V2/s1 [2]),
    .B(net8),
    .Z(\V3/V3/V2/A2/M3/s1 ));
 AND2_X1 \V3/V3/V2/A2/M3/M2/_0_  (.A1(\V3/V3/V2/A2/M3/s1 ),
    .A2(\V3/V3/V2/A2/c2 ),
    .ZN(\V3/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M3/M2/_1_  (.A(\V3/V3/V2/A2/M3/s1 ),
    .B(\V3/V3/V2/A2/c2 ),
    .Z(\V3/V3/V2/s2 [2]));
 OR2_X1 \V3/V3/V2/A2/M3/_0_  (.A1(\V3/V3/V2/A2/M3/c1 ),
    .A2(\V3/V3/V2/A2/M3/c2 ),
    .ZN(\V3/V3/V2/A2/c3 ));
 AND2_X1 \V3/V3/V2/A2/M4/M1/_0_  (.A1(\V3/V3/V2/s1 [3]),
    .A2(net8),
    .ZN(\V3/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A2/M4/M1/_1_  (.A(\V3/V3/V2/s1 [3]),
    .B(net8),
    .Z(\V3/V3/V2/A2/M4/s1 ));
 AND2_X1 \V3/V3/V2/A2/M4/M2/_0_  (.A1(\V3/V3/V2/A2/M4/s1 ),
    .A2(\V3/V3/V2/A2/c3 ),
    .ZN(\V3/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A2/M4/M2/_1_  (.A(\V3/V3/V2/A2/M4/s1 ),
    .B(\V3/V3/V2/A2/c3 ),
    .Z(\V3/V3/V2/s2 [3]));
 OR2_X1 \V3/V3/V2/A2/M4/_0_  (.A1(\V3/V3/V2/A2/M4/c1 ),
    .A2(\V3/V3/V2/A2/M4/c2 ),
    .ZN(\V3/V3/V2/c2 ));
 AND2_X1 \V3/V3/V2/A3/M1/M1/_0_  (.A1(\V3/V3/V2/v4 [0]),
    .A2(\V3/V3/V2/s2 [2]),
    .ZN(\V3/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M1/M1/_1_  (.A(\V3/V3/V2/v4 [0]),
    .B(\V3/V3/V2/s2 [2]),
    .Z(\V3/V3/V2/A3/M1/s1 ));
 AND2_X1 \V3/V3/V2/A3/M1/M2/_0_  (.A1(\V3/V3/V2/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M1/M2/_1_  (.A(\V3/V3/V2/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v2 [4]));
 OR2_X1 \V3/V3/V2/A3/M1/_0_  (.A1(\V3/V3/V2/A3/M1/c1 ),
    .A2(\V3/V3/V2/A3/M1/c2 ),
    .ZN(\V3/V3/V2/A3/c1 ));
 AND2_X1 \V3/V3/V2/A3/M2/M1/_0_  (.A1(\V3/V3/V2/v4 [1]),
    .A2(\V3/V3/V2/s2 [3]),
    .ZN(\V3/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M2/M1/_1_  (.A(\V3/V3/V2/v4 [1]),
    .B(\V3/V3/V2/s2 [3]),
    .Z(\V3/V3/V2/A3/M2/s1 ));
 AND2_X1 \V3/V3/V2/A3/M2/M2/_0_  (.A1(\V3/V3/V2/A3/M2/s1 ),
    .A2(\V3/V3/V2/A3/c1 ),
    .ZN(\V3/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M2/M2/_1_  (.A(\V3/V3/V2/A3/M2/s1 ),
    .B(\V3/V3/V2/A3/c1 ),
    .Z(\V3/V3/v2 [5]));
 OR2_X1 \V3/V3/V2/A3/M2/_0_  (.A1(\V3/V3/V2/A3/M2/c1 ),
    .A2(\V3/V3/V2/A3/M2/c2 ),
    .ZN(\V3/V3/V2/A3/c2 ));
 AND2_X1 \V3/V3/V2/A3/M3/M1/_0_  (.A1(\V3/V3/V2/v4 [2]),
    .A2(\V3/V3/V2/c3 ),
    .ZN(\V3/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M3/M1/_1_  (.A(\V3/V3/V2/v4 [2]),
    .B(\V3/V3/V2/c3 ),
    .Z(\V3/V3/V2/A3/M3/s1 ));
 AND2_X1 \V3/V3/V2/A3/M3/M2/_0_  (.A1(\V3/V3/V2/A3/M3/s1 ),
    .A2(\V3/V3/V2/A3/c2 ),
    .ZN(\V3/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M3/M2/_1_  (.A(\V3/V3/V2/A3/M3/s1 ),
    .B(\V3/V3/V2/A3/c2 ),
    .Z(\V3/V3/v2 [6]));
 OR2_X1 \V3/V3/V2/A3/M3/_0_  (.A1(\V3/V3/V2/A3/M3/c1 ),
    .A2(\V3/V3/V2/A3/M3/c2 ),
    .ZN(\V3/V3/V2/A3/c3 ));
 AND2_X1 \V3/V3/V2/A3/M4/M1/_0_  (.A1(\V3/V3/V2/v4 [3]),
    .A2(net8),
    .ZN(\V3/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V2/A3/M4/M1/_1_  (.A(\V3/V3/V2/v4 [3]),
    .B(net8),
    .Z(\V3/V3/V2/A3/M4/s1 ));
 AND2_X1 \V3/V3/V2/A3/M4/M2/_0_  (.A1(\V3/V3/V2/A3/M4/s1 ),
    .A2(\V3/V3/V2/A3/c3 ),
    .ZN(\V3/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V2/A3/M4/M2/_1_  (.A(\V3/V3/V2/A3/M4/s1 ),
    .B(\V3/V3/V2/A3/c3 ),
    .Z(\V3/V3/v2 [7]));
 OR2_X1 \V3/V3/V2/A3/M4/_0_  (.A1(\V3/V3/V2/A3/M4/c1 ),
    .A2(\V3/V3/V2/A3/M4/c2 ),
    .ZN(\V3/V3/V2/overflow ));
 AND2_X1 \V3/V3/V2/V1/HA1/_0_  (.A1(\V3/V3/V2/V1/w2 ),
    .A2(\V3/V3/V2/V1/w1 ),
    .ZN(\V3/V3/V2/V1/w4 ));
 XOR2_X2 \V3/V3/V2/V1/HA1/_1_  (.A(\V3/V3/V2/V1/w2 ),
    .B(\V3/V3/V2/V1/w1 ),
    .Z(\V3/V3/v2 [1]));
 AND2_X1 \V3/V3/V2/V1/HA2/_0_  (.A1(\V3/V3/V2/V1/w4 ),
    .A2(\V3/V3/V2/V1/w3 ),
    .ZN(\V3/V3/V2/v1 [3]));
 XOR2_X2 \V3/V3/V2/V1/HA2/_1_  (.A(\V3/V3/V2/V1/w4 ),
    .B(\V3/V3/V2/V1/w3 ),
    .Z(\V3/V3/V2/v1 [2]));
 AND2_X1 \V3/V3/V2/V1/_0_  (.A1(A[4]),
    .A2(net14),
    .ZN(\V3/V3/v2 [0]));
 AND2_X1 \V3/V3/V2/V1/_1_  (.A1(A[4]),
    .A2(B[25]),
    .ZN(\V3/V3/V2/V1/w1 ));
 AND2_X1 \V3/V3/V2/V1/_2_  (.A1(net14),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V1/w2 ));
 AND2_X1 \V3/V3/V2/V1/_3_  (.A1(B[25]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V1/w3 ));
 AND2_X1 \V3/V3/V2/V2/HA1/_0_  (.A1(\V3/V3/V2/V2/w2 ),
    .A2(\V3/V3/V2/V2/w1 ),
    .ZN(\V3/V3/V2/V2/w4 ));
 XOR2_X2 \V3/V3/V2/V2/HA1/_1_  (.A(\V3/V3/V2/V2/w2 ),
    .B(\V3/V3/V2/V2/w1 ),
    .Z(\V3/V3/V2/v2 [1]));
 AND2_X1 \V3/V3/V2/V2/HA2/_0_  (.A1(\V3/V3/V2/V2/w4 ),
    .A2(\V3/V3/V2/V2/w3 ),
    .ZN(\V3/V3/V2/v2 [3]));
 XOR2_X2 \V3/V3/V2/V2/HA2/_1_  (.A(\V3/V3/V2/V2/w4 ),
    .B(\V3/V3/V2/V2/w3 ),
    .Z(\V3/V3/V2/v2 [2]));
 AND2_X1 \V3/V3/V2/V2/_0_  (.A1(A[6]),
    .A2(net14),
    .ZN(\V3/V3/V2/v2 [0]));
 AND2_X1 \V3/V3/V2/V2/_1_  (.A1(A[6]),
    .A2(B[25]),
    .ZN(\V3/V3/V2/V2/w1 ));
 AND2_X1 \V3/V3/V2/V2/_2_  (.A1(net14),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V2/w2 ));
 AND2_X1 \V3/V3/V2/V2/_3_  (.A1(B[25]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V2/w3 ));
 AND2_X1 \V3/V3/V2/V3/HA1/_0_  (.A1(\V3/V3/V2/V3/w2 ),
    .A2(\V3/V3/V2/V3/w1 ),
    .ZN(\V3/V3/V2/V3/w4 ));
 XOR2_X2 \V3/V3/V2/V3/HA1/_1_  (.A(\V3/V3/V2/V3/w2 ),
    .B(\V3/V3/V2/V3/w1 ),
    .Z(\V3/V3/V2/v3 [1]));
 AND2_X1 \V3/V3/V2/V3/HA2/_0_  (.A1(\V3/V3/V2/V3/w4 ),
    .A2(\V3/V3/V2/V3/w3 ),
    .ZN(\V3/V3/V2/v3 [3]));
 XOR2_X2 \V3/V3/V2/V3/HA2/_1_  (.A(\V3/V3/V2/V3/w4 ),
    .B(\V3/V3/V2/V3/w3 ),
    .Z(\V3/V3/V2/v3 [2]));
 AND2_X1 \V3/V3/V2/V3/_0_  (.A1(A[4]),
    .A2(net13),
    .ZN(\V3/V3/V2/v3 [0]));
 AND2_X1 \V3/V3/V2/V3/_1_  (.A1(A[4]),
    .A2(B[27]),
    .ZN(\V3/V3/V2/V3/w1 ));
 AND2_X1 \V3/V3/V2/V3/_2_  (.A1(net13),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V3/w2 ));
 AND2_X1 \V3/V3/V2/V3/_3_  (.A1(B[27]),
    .A2(A[5]),
    .ZN(\V3/V3/V2/V3/w3 ));
 AND2_X1 \V3/V3/V2/V4/HA1/_0_  (.A1(\V3/V3/V2/V4/w2 ),
    .A2(\V3/V3/V2/V4/w1 ),
    .ZN(\V3/V3/V2/V4/w4 ));
 XOR2_X2 \V3/V3/V2/V4/HA1/_1_  (.A(\V3/V3/V2/V4/w2 ),
    .B(\V3/V3/V2/V4/w1 ),
    .Z(\V3/V3/V2/v4 [1]));
 AND2_X1 \V3/V3/V2/V4/HA2/_0_  (.A1(\V3/V3/V2/V4/w4 ),
    .A2(\V3/V3/V2/V4/w3 ),
    .ZN(\V3/V3/V2/v4 [3]));
 XOR2_X2 \V3/V3/V2/V4/HA2/_1_  (.A(\V3/V3/V2/V4/w4 ),
    .B(\V3/V3/V2/V4/w3 ),
    .Z(\V3/V3/V2/v4 [2]));
 AND2_X1 \V3/V3/V2/V4/_0_  (.A1(A[6]),
    .A2(net13),
    .ZN(\V3/V3/V2/v4 [0]));
 AND2_X1 \V3/V3/V2/V4/_1_  (.A1(A[6]),
    .A2(B[27]),
    .ZN(\V3/V3/V2/V4/w1 ));
 AND2_X1 \V3/V3/V2/V4/_2_  (.A1(net13),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V4/w2 ));
 AND2_X1 \V3/V3/V2/V4/_3_  (.A1(B[27]),
    .A2(A[7]),
    .ZN(\V3/V3/V2/V4/w3 ));
 OR2_X1 \V3/V3/V2/_0_  (.A1(\V3/V3/V2/c1 ),
    .A2(\V3/V3/V2/c2 ),
    .ZN(\V3/V3/V2/c3 ));
 AND2_X1 \V3/V3/V3/A1/M1/M1/_0_  (.A1(\V3/V3/V3/v2 [0]),
    .A2(\V3/V3/V3/v3 [0]),
    .ZN(\V3/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M1/M1/_1_  (.A(\V3/V3/V3/v2 [0]),
    .B(\V3/V3/V3/v3 [0]),
    .Z(\V3/V3/V3/A1/M1/s1 ));
 AND2_X1 \V3/V3/V3/A1/M1/M2/_0_  (.A1(\V3/V3/V3/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M1/M2/_1_  (.A(\V3/V3/V3/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/V3/s1 [0]));
 OR2_X1 \V3/V3/V3/A1/M1/_0_  (.A1(\V3/V3/V3/A1/M1/c1 ),
    .A2(\V3/V3/V3/A1/M1/c2 ),
    .ZN(\V3/V3/V3/A1/c1 ));
 AND2_X1 \V3/V3/V3/A1/M2/M1/_0_  (.A1(\V3/V3/V3/v2 [1]),
    .A2(\V3/V3/V3/v3 [1]),
    .ZN(\V3/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M2/M1/_1_  (.A(\V3/V3/V3/v2 [1]),
    .B(\V3/V3/V3/v3 [1]),
    .Z(\V3/V3/V3/A1/M2/s1 ));
 AND2_X1 \V3/V3/V3/A1/M2/M2/_0_  (.A1(\V3/V3/V3/A1/M2/s1 ),
    .A2(\V3/V3/V3/A1/c1 ),
    .ZN(\V3/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M2/M2/_1_  (.A(\V3/V3/V3/A1/M2/s1 ),
    .B(\V3/V3/V3/A1/c1 ),
    .Z(\V3/V3/V3/s1 [1]));
 OR2_X1 \V3/V3/V3/A1/M2/_0_  (.A1(\V3/V3/V3/A1/M2/c1 ),
    .A2(\V3/V3/V3/A1/M2/c2 ),
    .ZN(\V3/V3/V3/A1/c2 ));
 AND2_X1 \V3/V3/V3/A1/M3/M1/_0_  (.A1(\V3/V3/V3/v2 [2]),
    .A2(\V3/V3/V3/v3 [2]),
    .ZN(\V3/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M3/M1/_1_  (.A(\V3/V3/V3/v2 [2]),
    .B(\V3/V3/V3/v3 [2]),
    .Z(\V3/V3/V3/A1/M3/s1 ));
 AND2_X1 \V3/V3/V3/A1/M3/M2/_0_  (.A1(\V3/V3/V3/A1/M3/s1 ),
    .A2(\V3/V3/V3/A1/c2 ),
    .ZN(\V3/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M3/M2/_1_  (.A(\V3/V3/V3/A1/M3/s1 ),
    .B(\V3/V3/V3/A1/c2 ),
    .Z(\V3/V3/V3/s1 [2]));
 OR2_X1 \V3/V3/V3/A1/M3/_0_  (.A1(\V3/V3/V3/A1/M3/c1 ),
    .A2(\V3/V3/V3/A1/M3/c2 ),
    .ZN(\V3/V3/V3/A1/c3 ));
 AND2_X1 \V3/V3/V3/A1/M4/M1/_0_  (.A1(\V3/V3/V3/v2 [3]),
    .A2(\V3/V3/V3/v3 [3]),
    .ZN(\V3/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A1/M4/M1/_1_  (.A(\V3/V3/V3/v2 [3]),
    .B(\V3/V3/V3/v3 [3]),
    .Z(\V3/V3/V3/A1/M4/s1 ));
 AND2_X1 \V3/V3/V3/A1/M4/M2/_0_  (.A1(\V3/V3/V3/A1/M4/s1 ),
    .A2(\V3/V3/V3/A1/c3 ),
    .ZN(\V3/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A1/M4/M2/_1_  (.A(\V3/V3/V3/A1/M4/s1 ),
    .B(\V3/V3/V3/A1/c3 ),
    .Z(\V3/V3/V3/s1 [3]));
 OR2_X1 \V3/V3/V3/A1/M4/_0_  (.A1(\V3/V3/V3/A1/M4/c1 ),
    .A2(\V3/V3/V3/A1/M4/c2 ),
    .ZN(\V3/V3/V3/c1 ));
 AND2_X1 \V3/V3/V3/A2/M1/M1/_0_  (.A1(\V3/V3/V3/s1 [0]),
    .A2(\V3/V3/V3/v1 [2]),
    .ZN(\V3/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M1/M1/_1_  (.A(\V3/V3/V3/s1 [0]),
    .B(\V3/V3/V3/v1 [2]),
    .Z(\V3/V3/V3/A2/M1/s1 ));
 AND2_X1 \V3/V3/V3/A2/M1/M2/_0_  (.A1(\V3/V3/V3/A2/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M1/M2/_1_  (.A(\V3/V3/V3/A2/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v3 [2]));
 OR2_X1 \V3/V3/V3/A2/M1/_0_  (.A1(\V3/V3/V3/A2/M1/c1 ),
    .A2(\V3/V3/V3/A2/M1/c2 ),
    .ZN(\V3/V3/V3/A2/c1 ));
 AND2_X1 \V3/V3/V3/A2/M2/M1/_0_  (.A1(\V3/V3/V3/s1 [1]),
    .A2(\V3/V3/V3/v1 [3]),
    .ZN(\V3/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M2/M1/_1_  (.A(\V3/V3/V3/s1 [1]),
    .B(\V3/V3/V3/v1 [3]),
    .Z(\V3/V3/V3/A2/M2/s1 ));
 AND2_X1 \V3/V3/V3/A2/M2/M2/_0_  (.A1(\V3/V3/V3/A2/M2/s1 ),
    .A2(\V3/V3/V3/A2/c1 ),
    .ZN(\V3/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M2/M2/_1_  (.A(\V3/V3/V3/A2/M2/s1 ),
    .B(\V3/V3/V3/A2/c1 ),
    .Z(\V3/V3/v3 [3]));
 OR2_X1 \V3/V3/V3/A2/M2/_0_  (.A1(\V3/V3/V3/A2/M2/c1 ),
    .A2(\V3/V3/V3/A2/M2/c2 ),
    .ZN(\V3/V3/V3/A2/c2 ));
 AND2_X1 \V3/V3/V3/A2/M3/M1/_0_  (.A1(\V3/V3/V3/s1 [2]),
    .A2(net8),
    .ZN(\V3/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M3/M1/_1_  (.A(\V3/V3/V3/s1 [2]),
    .B(net8),
    .Z(\V3/V3/V3/A2/M3/s1 ));
 AND2_X1 \V3/V3/V3/A2/M3/M2/_0_  (.A1(\V3/V3/V3/A2/M3/s1 ),
    .A2(\V3/V3/V3/A2/c2 ),
    .ZN(\V3/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M3/M2/_1_  (.A(\V3/V3/V3/A2/M3/s1 ),
    .B(\V3/V3/V3/A2/c2 ),
    .Z(\V3/V3/V3/s2 [2]));
 OR2_X1 \V3/V3/V3/A2/M3/_0_  (.A1(\V3/V3/V3/A2/M3/c1 ),
    .A2(\V3/V3/V3/A2/M3/c2 ),
    .ZN(\V3/V3/V3/A2/c3 ));
 AND2_X1 \V3/V3/V3/A2/M4/M1/_0_  (.A1(\V3/V3/V3/s1 [3]),
    .A2(net8),
    .ZN(\V3/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A2/M4/M1/_1_  (.A(\V3/V3/V3/s1 [3]),
    .B(net8),
    .Z(\V3/V3/V3/A2/M4/s1 ));
 AND2_X1 \V3/V3/V3/A2/M4/M2/_0_  (.A1(\V3/V3/V3/A2/M4/s1 ),
    .A2(\V3/V3/V3/A2/c3 ),
    .ZN(\V3/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A2/M4/M2/_1_  (.A(\V3/V3/V3/A2/M4/s1 ),
    .B(\V3/V3/V3/A2/c3 ),
    .Z(\V3/V3/V3/s2 [3]));
 OR2_X1 \V3/V3/V3/A2/M4/_0_  (.A1(\V3/V3/V3/A2/M4/c1 ),
    .A2(\V3/V3/V3/A2/M4/c2 ),
    .ZN(\V3/V3/V3/c2 ));
 AND2_X1 \V3/V3/V3/A3/M1/M1/_0_  (.A1(\V3/V3/V3/v4 [0]),
    .A2(\V3/V3/V3/s2 [2]),
    .ZN(\V3/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M1/M1/_1_  (.A(\V3/V3/V3/v4 [0]),
    .B(\V3/V3/V3/s2 [2]),
    .Z(\V3/V3/V3/A3/M1/s1 ));
 AND2_X1 \V3/V3/V3/A3/M1/M2/_0_  (.A1(\V3/V3/V3/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M1/M2/_1_  (.A(\V3/V3/V3/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v3 [4]));
 OR2_X1 \V3/V3/V3/A3/M1/_0_  (.A1(\V3/V3/V3/A3/M1/c1 ),
    .A2(\V3/V3/V3/A3/M1/c2 ),
    .ZN(\V3/V3/V3/A3/c1 ));
 AND2_X1 \V3/V3/V3/A3/M2/M1/_0_  (.A1(\V3/V3/V3/v4 [1]),
    .A2(\V3/V3/V3/s2 [3]),
    .ZN(\V3/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M2/M1/_1_  (.A(\V3/V3/V3/v4 [1]),
    .B(\V3/V3/V3/s2 [3]),
    .Z(\V3/V3/V3/A3/M2/s1 ));
 AND2_X1 \V3/V3/V3/A3/M2/M2/_0_  (.A1(\V3/V3/V3/A3/M2/s1 ),
    .A2(\V3/V3/V3/A3/c1 ),
    .ZN(\V3/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M2/M2/_1_  (.A(\V3/V3/V3/A3/M2/s1 ),
    .B(\V3/V3/V3/A3/c1 ),
    .Z(\V3/V3/v3 [5]));
 OR2_X1 \V3/V3/V3/A3/M2/_0_  (.A1(\V3/V3/V3/A3/M2/c1 ),
    .A2(\V3/V3/V3/A3/M2/c2 ),
    .ZN(\V3/V3/V3/A3/c2 ));
 AND2_X1 \V3/V3/V3/A3/M3/M1/_0_  (.A1(\V3/V3/V3/v4 [2]),
    .A2(\V3/V3/V3/c3 ),
    .ZN(\V3/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M3/M1/_1_  (.A(\V3/V3/V3/v4 [2]),
    .B(\V3/V3/V3/c3 ),
    .Z(\V3/V3/V3/A3/M3/s1 ));
 AND2_X1 \V3/V3/V3/A3/M3/M2/_0_  (.A1(\V3/V3/V3/A3/M3/s1 ),
    .A2(\V3/V3/V3/A3/c2 ),
    .ZN(\V3/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M3/M2/_1_  (.A(\V3/V3/V3/A3/M3/s1 ),
    .B(\V3/V3/V3/A3/c2 ),
    .Z(\V3/V3/v3 [6]));
 OR2_X1 \V3/V3/V3/A3/M3/_0_  (.A1(\V3/V3/V3/A3/M3/c1 ),
    .A2(\V3/V3/V3/A3/M3/c2 ),
    .ZN(\V3/V3/V3/A3/c3 ));
 AND2_X1 \V3/V3/V3/A3/M4/M1/_0_  (.A1(\V3/V3/V3/v4 [3]),
    .A2(net8),
    .ZN(\V3/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V3/A3/M4/M1/_1_  (.A(\V3/V3/V3/v4 [3]),
    .B(net8),
    .Z(\V3/V3/V3/A3/M4/s1 ));
 AND2_X1 \V3/V3/V3/A3/M4/M2/_0_  (.A1(\V3/V3/V3/A3/M4/s1 ),
    .A2(\V3/V3/V3/A3/c3 ),
    .ZN(\V3/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V3/A3/M4/M2/_1_  (.A(\V3/V3/V3/A3/M4/s1 ),
    .B(\V3/V3/V3/A3/c3 ),
    .Z(\V3/V3/v3 [7]));
 OR2_X1 \V3/V3/V3/A3/M4/_0_  (.A1(\V3/V3/V3/A3/M4/c1 ),
    .A2(\V3/V3/V3/A3/M4/c2 ),
    .ZN(\V3/V3/V3/overflow ));
 AND2_X1 \V3/V3/V3/V1/HA1/_0_  (.A1(\V3/V3/V3/V1/w2 ),
    .A2(\V3/V3/V3/V1/w1 ),
    .ZN(\V3/V3/V3/V1/w4 ));
 XOR2_X2 \V3/V3/V3/V1/HA1/_1_  (.A(\V3/V3/V3/V1/w2 ),
    .B(\V3/V3/V3/V1/w1 ),
    .Z(\V3/V3/v3 [1]));
 AND2_X1 \V3/V3/V3/V1/HA2/_0_  (.A1(\V3/V3/V3/V1/w4 ),
    .A2(\V3/V3/V3/V1/w3 ),
    .ZN(\V3/V3/V3/v1 [3]));
 XOR2_X2 \V3/V3/V3/V1/HA2/_1_  (.A(\V3/V3/V3/V1/w4 ),
    .B(\V3/V3/V3/V1/w3 ),
    .Z(\V3/V3/V3/v1 [2]));
 AND2_X1 \V3/V3/V3/V1/_0_  (.A1(net48),
    .A2(B[28]),
    .ZN(\V3/V3/v3 [0]));
 AND2_X1 \V3/V3/V3/V1/_1_  (.A1(net48),
    .A2(B[29]),
    .ZN(\V3/V3/V3/V1/w1 ));
 AND2_X1 \V3/V3/V3/V1/_2_  (.A1(B[28]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V1/w2 ));
 AND2_X1 \V3/V3/V3/V1/_3_  (.A1(B[29]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V1/w3 ));
 AND2_X1 \V3/V3/V3/V2/HA1/_0_  (.A1(\V3/V3/V3/V2/w2 ),
    .A2(\V3/V3/V3/V2/w1 ),
    .ZN(\V3/V3/V3/V2/w4 ));
 XOR2_X2 \V3/V3/V3/V2/HA1/_1_  (.A(\V3/V3/V3/V2/w2 ),
    .B(\V3/V3/V3/V2/w1 ),
    .Z(\V3/V3/V3/v2 [1]));
 AND2_X1 \V3/V3/V3/V2/HA2/_0_  (.A1(\V3/V3/V3/V2/w4 ),
    .A2(\V3/V3/V3/V2/w3 ),
    .ZN(\V3/V3/V3/v2 [3]));
 XOR2_X2 \V3/V3/V3/V2/HA2/_1_  (.A(\V3/V3/V3/V2/w4 ),
    .B(\V3/V3/V3/V2/w3 ),
    .Z(\V3/V3/V3/v2 [2]));
 AND2_X1 \V3/V3/V3/V2/_0_  (.A1(A[2]),
    .A2(B[28]),
    .ZN(\V3/V3/V3/v2 [0]));
 AND2_X1 \V3/V3/V3/V2/_1_  (.A1(A[2]),
    .A2(B[29]),
    .ZN(\V3/V3/V3/V2/w1 ));
 AND2_X1 \V3/V3/V3/V2/_2_  (.A1(B[28]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V2/w2 ));
 AND2_X1 \V3/V3/V3/V2/_3_  (.A1(B[29]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V2/w3 ));
 AND2_X1 \V3/V3/V3/V3/HA1/_0_  (.A1(\V3/V3/V3/V3/w2 ),
    .A2(\V3/V3/V3/V3/w1 ),
    .ZN(\V3/V3/V3/V3/w4 ));
 XOR2_X2 \V3/V3/V3/V3/HA1/_1_  (.A(\V3/V3/V3/V3/w2 ),
    .B(\V3/V3/V3/V3/w1 ),
    .Z(\V3/V3/V3/v3 [1]));
 AND2_X1 \V3/V3/V3/V3/HA2/_0_  (.A1(\V3/V3/V3/V3/w4 ),
    .A2(\V3/V3/V3/V3/w3 ),
    .ZN(\V3/V3/V3/v3 [3]));
 XOR2_X2 \V3/V3/V3/V3/HA2/_1_  (.A(\V3/V3/V3/V3/w4 ),
    .B(\V3/V3/V3/V3/w3 ),
    .Z(\V3/V3/V3/v3 [2]));
 AND2_X1 \V3/V3/V3/V3/_0_  (.A1(net48),
    .A2(B[30]),
    .ZN(\V3/V3/V3/v3 [0]));
 AND2_X1 \V3/V3/V3/V3/_1_  (.A1(net48),
    .A2(B[31]),
    .ZN(\V3/V3/V3/V3/w1 ));
 AND2_X1 \V3/V3/V3/V3/_2_  (.A1(B[30]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V3/w2 ));
 AND2_X1 \V3/V3/V3/V3/_3_  (.A1(B[31]),
    .A2(A[1]),
    .ZN(\V3/V3/V3/V3/w3 ));
 AND2_X1 \V3/V3/V3/V4/HA1/_0_  (.A1(\V3/V3/V3/V4/w2 ),
    .A2(\V3/V3/V3/V4/w1 ),
    .ZN(\V3/V3/V3/V4/w4 ));
 XOR2_X2 \V3/V3/V3/V4/HA1/_1_  (.A(\V3/V3/V3/V4/w2 ),
    .B(\V3/V3/V3/V4/w1 ),
    .Z(\V3/V3/V3/v4 [1]));
 AND2_X1 \V3/V3/V3/V4/HA2/_0_  (.A1(\V3/V3/V3/V4/w4 ),
    .A2(\V3/V3/V3/V4/w3 ),
    .ZN(\V3/V3/V3/v4 [3]));
 XOR2_X2 \V3/V3/V3/V4/HA2/_1_  (.A(\V3/V3/V3/V4/w4 ),
    .B(\V3/V3/V3/V4/w3 ),
    .Z(\V3/V3/V3/v4 [2]));
 AND2_X1 \V3/V3/V3/V4/_0_  (.A1(A[2]),
    .A2(B[30]),
    .ZN(\V3/V3/V3/v4 [0]));
 AND2_X1 \V3/V3/V3/V4/_1_  (.A1(A[2]),
    .A2(B[31]),
    .ZN(\V3/V3/V3/V4/w1 ));
 AND2_X1 \V3/V3/V3/V4/_2_  (.A1(B[30]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V4/w2 ));
 AND2_X1 \V3/V3/V3/V4/_3_  (.A1(B[31]),
    .A2(A[3]),
    .ZN(\V3/V3/V3/V4/w3 ));
 OR2_X1 \V3/V3/V3/_0_  (.A1(\V3/V3/V3/c1 ),
    .A2(\V3/V3/V3/c2 ),
    .ZN(\V3/V3/V3/c3 ));
 AND2_X1 \V3/V3/V4/A1/M1/M1/_0_  (.A1(\V3/V3/V4/v2 [0]),
    .A2(\V3/V3/V4/v3 [0]),
    .ZN(\V3/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M1/M1/_1_  (.A(\V3/V3/V4/v2 [0]),
    .B(\V3/V3/V4/v3 [0]),
    .Z(\V3/V3/V4/A1/M1/s1 ));
 AND2_X1 \V3/V3/V4/A1/M1/M2/_0_  (.A1(\V3/V3/V4/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M1/M2/_1_  (.A(\V3/V3/V4/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/V4/s1 [0]));
 OR2_X1 \V3/V3/V4/A1/M1/_0_  (.A1(\V3/V3/V4/A1/M1/c1 ),
    .A2(\V3/V3/V4/A1/M1/c2 ),
    .ZN(\V3/V3/V4/A1/c1 ));
 AND2_X1 \V3/V3/V4/A1/M2/M1/_0_  (.A1(\V3/V3/V4/v2 [1]),
    .A2(\V3/V3/V4/v3 [1]),
    .ZN(\V3/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M2/M1/_1_  (.A(\V3/V3/V4/v2 [1]),
    .B(\V3/V3/V4/v3 [1]),
    .Z(\V3/V3/V4/A1/M2/s1 ));
 AND2_X1 \V3/V3/V4/A1/M2/M2/_0_  (.A1(\V3/V3/V4/A1/M2/s1 ),
    .A2(\V3/V3/V4/A1/c1 ),
    .ZN(\V3/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M2/M2/_1_  (.A(\V3/V3/V4/A1/M2/s1 ),
    .B(\V3/V3/V4/A1/c1 ),
    .Z(\V3/V3/V4/s1 [1]));
 OR2_X1 \V3/V3/V4/A1/M2/_0_  (.A1(\V3/V3/V4/A1/M2/c1 ),
    .A2(\V3/V3/V4/A1/M2/c2 ),
    .ZN(\V3/V3/V4/A1/c2 ));
 AND2_X1 \V3/V3/V4/A1/M3/M1/_0_  (.A1(\V3/V3/V4/v2 [2]),
    .A2(\V3/V3/V4/v3 [2]),
    .ZN(\V3/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M3/M1/_1_  (.A(\V3/V3/V4/v2 [2]),
    .B(\V3/V3/V4/v3 [2]),
    .Z(\V3/V3/V4/A1/M3/s1 ));
 AND2_X1 \V3/V3/V4/A1/M3/M2/_0_  (.A1(\V3/V3/V4/A1/M3/s1 ),
    .A2(\V3/V3/V4/A1/c2 ),
    .ZN(\V3/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M3/M2/_1_  (.A(\V3/V3/V4/A1/M3/s1 ),
    .B(\V3/V3/V4/A1/c2 ),
    .Z(\V3/V3/V4/s1 [2]));
 OR2_X1 \V3/V3/V4/A1/M3/_0_  (.A1(\V3/V3/V4/A1/M3/c1 ),
    .A2(\V3/V3/V4/A1/M3/c2 ),
    .ZN(\V3/V3/V4/A1/c3 ));
 AND2_X1 \V3/V3/V4/A1/M4/M1/_0_  (.A1(\V3/V3/V4/v2 [3]),
    .A2(\V3/V3/V4/v3 [3]),
    .ZN(\V3/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A1/M4/M1/_1_  (.A(\V3/V3/V4/v2 [3]),
    .B(\V3/V3/V4/v3 [3]),
    .Z(\V3/V3/V4/A1/M4/s1 ));
 AND2_X1 \V3/V3/V4/A1/M4/M2/_0_  (.A1(\V3/V3/V4/A1/M4/s1 ),
    .A2(\V3/V3/V4/A1/c3 ),
    .ZN(\V3/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A1/M4/M2/_1_  (.A(\V3/V3/V4/A1/M4/s1 ),
    .B(\V3/V3/V4/A1/c3 ),
    .Z(\V3/V3/V4/s1 [3]));
 OR2_X1 \V3/V3/V4/A1/M4/_0_  (.A1(\V3/V3/V4/A1/M4/c1 ),
    .A2(\V3/V3/V4/A1/M4/c2 ),
    .ZN(\V3/V3/V4/c1 ));
 AND2_X1 \V3/V3/V4/A2/M1/M1/_0_  (.A1(\V3/V3/V4/s1 [0]),
    .A2(\V3/V3/V4/v1 [2]),
    .ZN(\V3/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M1/M1/_1_  (.A(\V3/V3/V4/s1 [0]),
    .B(\V3/V3/V4/v1 [2]),
    .Z(\V3/V3/V4/A2/M1/s1 ));
 AND2_X1 \V3/V3/V4/A2/M1/M2/_0_  (.A1(\V3/V3/V4/A2/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M1/M2/_1_  (.A(\V3/V3/V4/A2/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v4 [2]));
 OR2_X1 \V3/V3/V4/A2/M1/_0_  (.A1(\V3/V3/V4/A2/M1/c1 ),
    .A2(\V3/V3/V4/A2/M1/c2 ),
    .ZN(\V3/V3/V4/A2/c1 ));
 AND2_X1 \V3/V3/V4/A2/M2/M1/_0_  (.A1(\V3/V3/V4/s1 [1]),
    .A2(\V3/V3/V4/v1 [3]),
    .ZN(\V3/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M2/M1/_1_  (.A(\V3/V3/V4/s1 [1]),
    .B(\V3/V3/V4/v1 [3]),
    .Z(\V3/V3/V4/A2/M2/s1 ));
 AND2_X1 \V3/V3/V4/A2/M2/M2/_0_  (.A1(\V3/V3/V4/A2/M2/s1 ),
    .A2(\V3/V3/V4/A2/c1 ),
    .ZN(\V3/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M2/M2/_1_  (.A(\V3/V3/V4/A2/M2/s1 ),
    .B(\V3/V3/V4/A2/c1 ),
    .Z(\V3/V3/v4 [3]));
 OR2_X1 \V3/V3/V4/A2/M2/_0_  (.A1(\V3/V3/V4/A2/M2/c1 ),
    .A2(\V3/V3/V4/A2/M2/c2 ),
    .ZN(\V3/V3/V4/A2/c2 ));
 AND2_X1 \V3/V3/V4/A2/M3/M1/_0_  (.A1(\V3/V3/V4/s1 [2]),
    .A2(net8),
    .ZN(\V3/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M3/M1/_1_  (.A(\V3/V3/V4/s1 [2]),
    .B(net8),
    .Z(\V3/V3/V4/A2/M3/s1 ));
 AND2_X1 \V3/V3/V4/A2/M3/M2/_0_  (.A1(\V3/V3/V4/A2/M3/s1 ),
    .A2(\V3/V3/V4/A2/c2 ),
    .ZN(\V3/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M3/M2/_1_  (.A(\V3/V3/V4/A2/M3/s1 ),
    .B(\V3/V3/V4/A2/c2 ),
    .Z(\V3/V3/V4/s2 [2]));
 OR2_X1 \V3/V3/V4/A2/M3/_0_  (.A1(\V3/V3/V4/A2/M3/c1 ),
    .A2(\V3/V3/V4/A2/M3/c2 ),
    .ZN(\V3/V3/V4/A2/c3 ));
 AND2_X1 \V3/V3/V4/A2/M4/M1/_0_  (.A1(\V3/V3/V4/s1 [3]),
    .A2(net8),
    .ZN(\V3/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A2/M4/M1/_1_  (.A(\V3/V3/V4/s1 [3]),
    .B(net8),
    .Z(\V3/V3/V4/A2/M4/s1 ));
 AND2_X1 \V3/V3/V4/A2/M4/M2/_0_  (.A1(\V3/V3/V4/A2/M4/s1 ),
    .A2(\V3/V3/V4/A2/c3 ),
    .ZN(\V3/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A2/M4/M2/_1_  (.A(\V3/V3/V4/A2/M4/s1 ),
    .B(\V3/V3/V4/A2/c3 ),
    .Z(\V3/V3/V4/s2 [3]));
 OR2_X1 \V3/V3/V4/A2/M4/_0_  (.A1(\V3/V3/V4/A2/M4/c1 ),
    .A2(\V3/V3/V4/A2/M4/c2 ),
    .ZN(\V3/V3/V4/c2 ));
 AND2_X1 \V3/V3/V4/A3/M1/M1/_0_  (.A1(\V3/V3/V4/v4 [0]),
    .A2(\V3/V3/V4/s2 [2]),
    .ZN(\V3/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M1/M1/_1_  (.A(\V3/V3/V4/v4 [0]),
    .B(\V3/V3/V4/s2 [2]),
    .Z(\V3/V3/V4/A3/M1/s1 ));
 AND2_X1 \V3/V3/V4/A3/M1/M2/_0_  (.A1(\V3/V3/V4/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M1/M2/_1_  (.A(\V3/V3/V4/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V3/v4 [4]));
 OR2_X1 \V3/V3/V4/A3/M1/_0_  (.A1(\V3/V3/V4/A3/M1/c1 ),
    .A2(\V3/V3/V4/A3/M1/c2 ),
    .ZN(\V3/V3/V4/A3/c1 ));
 AND2_X1 \V3/V3/V4/A3/M2/M1/_0_  (.A1(\V3/V3/V4/v4 [1]),
    .A2(\V3/V3/V4/s2 [3]),
    .ZN(\V3/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M2/M1/_1_  (.A(\V3/V3/V4/v4 [1]),
    .B(\V3/V3/V4/s2 [3]),
    .Z(\V3/V3/V4/A3/M2/s1 ));
 AND2_X1 \V3/V3/V4/A3/M2/M2/_0_  (.A1(\V3/V3/V4/A3/M2/s1 ),
    .A2(\V3/V3/V4/A3/c1 ),
    .ZN(\V3/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M2/M2/_1_  (.A(\V3/V3/V4/A3/M2/s1 ),
    .B(\V3/V3/V4/A3/c1 ),
    .Z(\V3/V3/v4 [5]));
 OR2_X1 \V3/V3/V4/A3/M2/_0_  (.A1(\V3/V3/V4/A3/M2/c1 ),
    .A2(\V3/V3/V4/A3/M2/c2 ),
    .ZN(\V3/V3/V4/A3/c2 ));
 AND2_X1 \V3/V3/V4/A3/M3/M1/_0_  (.A1(\V3/V3/V4/v4 [2]),
    .A2(\V3/V3/V4/c3 ),
    .ZN(\V3/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M3/M1/_1_  (.A(\V3/V3/V4/v4 [2]),
    .B(\V3/V3/V4/c3 ),
    .Z(\V3/V3/V4/A3/M3/s1 ));
 AND2_X1 \V3/V3/V4/A3/M3/M2/_0_  (.A1(\V3/V3/V4/A3/M3/s1 ),
    .A2(\V3/V3/V4/A3/c2 ),
    .ZN(\V3/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M3/M2/_1_  (.A(\V3/V3/V4/A3/M3/s1 ),
    .B(\V3/V3/V4/A3/c2 ),
    .Z(\V3/V3/v4 [6]));
 OR2_X1 \V3/V3/V4/A3/M3/_0_  (.A1(\V3/V3/V4/A3/M3/c1 ),
    .A2(\V3/V3/V4/A3/M3/c2 ),
    .ZN(\V3/V3/V4/A3/c3 ));
 AND2_X1 \V3/V3/V4/A3/M4/M1/_0_  (.A1(\V3/V3/V4/v4 [3]),
    .A2(net8),
    .ZN(\V3/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V3/V4/A3/M4/M1/_1_  (.A(\V3/V3/V4/v4 [3]),
    .B(net8),
    .Z(\V3/V3/V4/A3/M4/s1 ));
 AND2_X1 \V3/V3/V4/A3/M4/M2/_0_  (.A1(\V3/V3/V4/A3/M4/s1 ),
    .A2(\V3/V3/V4/A3/c3 ),
    .ZN(\V3/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V3/V4/A3/M4/M2/_1_  (.A(\V3/V3/V4/A3/M4/s1 ),
    .B(\V3/V3/V4/A3/c3 ),
    .Z(\V3/V3/v4 [7]));
 OR2_X1 \V3/V3/V4/A3/M4/_0_  (.A1(\V3/V3/V4/A3/M4/c1 ),
    .A2(\V3/V3/V4/A3/M4/c2 ),
    .ZN(\V3/V3/V4/overflow ));
 AND2_X1 \V3/V3/V4/V1/HA1/_0_  (.A1(\V3/V3/V4/V1/w2 ),
    .A2(\V3/V3/V4/V1/w1 ),
    .ZN(\V3/V3/V4/V1/w4 ));
 XOR2_X2 \V3/V3/V4/V1/HA1/_1_  (.A(\V3/V3/V4/V1/w2 ),
    .B(\V3/V3/V4/V1/w1 ),
    .Z(\V3/V3/v4 [1]));
 AND2_X1 \V3/V3/V4/V1/HA2/_0_  (.A1(\V3/V3/V4/V1/w4 ),
    .A2(\V3/V3/V4/V1/w3 ),
    .ZN(\V3/V3/V4/v1 [3]));
 XOR2_X2 \V3/V3/V4/V1/HA2/_1_  (.A(\V3/V3/V4/V1/w4 ),
    .B(\V3/V3/V4/V1/w3 ),
    .Z(\V3/V3/V4/v1 [2]));
 AND2_X1 \V3/V3/V4/V1/_0_  (.A1(A[4]),
    .A2(B[28]),
    .ZN(\V3/V3/v4 [0]));
 AND2_X1 \V3/V3/V4/V1/_1_  (.A1(A[4]),
    .A2(B[29]),
    .ZN(\V3/V3/V4/V1/w1 ));
 AND2_X1 \V3/V3/V4/V1/_2_  (.A1(B[28]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V1/w2 ));
 AND2_X1 \V3/V3/V4/V1/_3_  (.A1(B[29]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V1/w3 ));
 AND2_X1 \V3/V3/V4/V2/HA1/_0_  (.A1(\V3/V3/V4/V2/w2 ),
    .A2(\V3/V3/V4/V2/w1 ),
    .ZN(\V3/V3/V4/V2/w4 ));
 XOR2_X2 \V3/V3/V4/V2/HA1/_1_  (.A(\V3/V3/V4/V2/w2 ),
    .B(\V3/V3/V4/V2/w1 ),
    .Z(\V3/V3/V4/v2 [1]));
 AND2_X1 \V3/V3/V4/V2/HA2/_0_  (.A1(\V3/V3/V4/V2/w4 ),
    .A2(\V3/V3/V4/V2/w3 ),
    .ZN(\V3/V3/V4/v2 [3]));
 XOR2_X2 \V3/V3/V4/V2/HA2/_1_  (.A(\V3/V3/V4/V2/w4 ),
    .B(\V3/V3/V4/V2/w3 ),
    .Z(\V3/V3/V4/v2 [2]));
 AND2_X1 \V3/V3/V4/V2/_0_  (.A1(A[6]),
    .A2(B[28]),
    .ZN(\V3/V3/V4/v2 [0]));
 AND2_X1 \V3/V3/V4/V2/_1_  (.A1(A[6]),
    .A2(B[29]),
    .ZN(\V3/V3/V4/V2/w1 ));
 AND2_X1 \V3/V3/V4/V2/_2_  (.A1(B[28]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V2/w2 ));
 AND2_X1 \V3/V3/V4/V2/_3_  (.A1(B[29]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V2/w3 ));
 AND2_X1 \V3/V3/V4/V3/HA1/_0_  (.A1(\V3/V3/V4/V3/w2 ),
    .A2(\V3/V3/V4/V3/w1 ),
    .ZN(\V3/V3/V4/V3/w4 ));
 XOR2_X2 \V3/V3/V4/V3/HA1/_1_  (.A(\V3/V3/V4/V3/w2 ),
    .B(\V3/V3/V4/V3/w1 ),
    .Z(\V3/V3/V4/v3 [1]));
 AND2_X1 \V3/V3/V4/V3/HA2/_0_  (.A1(\V3/V3/V4/V3/w4 ),
    .A2(\V3/V3/V4/V3/w3 ),
    .ZN(\V3/V3/V4/v3 [3]));
 XOR2_X2 \V3/V3/V4/V3/HA2/_1_  (.A(\V3/V3/V4/V3/w4 ),
    .B(\V3/V3/V4/V3/w3 ),
    .Z(\V3/V3/V4/v3 [2]));
 AND2_X1 \V3/V3/V4/V3/_0_  (.A1(A[4]),
    .A2(B[30]),
    .ZN(\V3/V3/V4/v3 [0]));
 AND2_X1 \V3/V3/V4/V3/_1_  (.A1(A[4]),
    .A2(B[31]),
    .ZN(\V3/V3/V4/V3/w1 ));
 AND2_X1 \V3/V3/V4/V3/_2_  (.A1(B[30]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V3/w2 ));
 AND2_X1 \V3/V3/V4/V3/_3_  (.A1(B[31]),
    .A2(A[5]),
    .ZN(\V3/V3/V4/V3/w3 ));
 AND2_X1 \V3/V3/V4/V4/HA1/_0_  (.A1(\V3/V3/V4/V4/w2 ),
    .A2(\V3/V3/V4/V4/w1 ),
    .ZN(\V3/V3/V4/V4/w4 ));
 XOR2_X2 \V3/V3/V4/V4/HA1/_1_  (.A(\V3/V3/V4/V4/w2 ),
    .B(\V3/V3/V4/V4/w1 ),
    .Z(\V3/V3/V4/v4 [1]));
 AND2_X1 \V3/V3/V4/V4/HA2/_0_  (.A1(\V3/V3/V4/V4/w4 ),
    .A2(\V3/V3/V4/V4/w3 ),
    .ZN(\V3/V3/V4/v4 [3]));
 XOR2_X2 \V3/V3/V4/V4/HA2/_1_  (.A(\V3/V3/V4/V4/w4 ),
    .B(\V3/V3/V4/V4/w3 ),
    .Z(\V3/V3/V4/v4 [2]));
 AND2_X1 \V3/V3/V4/V4/_0_  (.A1(A[6]),
    .A2(B[30]),
    .ZN(\V3/V3/V4/v4 [0]));
 AND2_X1 \V3/V3/V4/V4/_1_  (.A1(A[6]),
    .A2(B[31]),
    .ZN(\V3/V3/V4/V4/w1 ));
 AND2_X1 \V3/V3/V4/V4/_2_  (.A1(B[30]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V4/w2 ));
 AND2_X1 \V3/V3/V4/V4/_3_  (.A1(B[31]),
    .A2(A[7]),
    .ZN(\V3/V3/V4/V4/w3 ));
 OR2_X1 \V3/V3/V4/_0_  (.A1(\V3/V3/V4/c1 ),
    .A2(\V3/V3/V4/c2 ),
    .ZN(\V3/V3/V4/c3 ));
 OR2_X1 \V3/V3/_0_  (.A1(\V3/V3/c1 ),
    .A2(\V3/V3/c2 ),
    .ZN(\V3/V3/c3 ));
 AND2_X1 \V3/V4/A1/A1/M1/M1/_0_  (.A1(\V3/V4/v2 [0]),
    .A2(\V3/V4/v3 [0]),
    .ZN(\V3/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M1/M1/_1_  (.A(\V3/V4/v2 [0]),
    .B(\V3/V4/v3 [0]),
    .Z(\V3/V4/A1/A1/M1/s1 ));
 AND2_X1 \V3/V4/A1/A1/M1/M2/_0_  (.A1(\V3/V4/A1/A1/M1/s1 ),
    .A2(net5),
    .ZN(\V3/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M1/M2/_1_  (.A(\V3/V4/A1/A1/M1/s1 ),
    .B(net5),
    .Z(\V3/V4/s1 [0]));
 OR2_X1 \V3/V4/A1/A1/M1/_0_  (.A1(\V3/V4/A1/A1/M1/c1 ),
    .A2(\V3/V4/A1/A1/M1/c2 ),
    .ZN(\V3/V4/A1/A1/c1 ));
 AND2_X1 \V3/V4/A1/A1/M2/M1/_0_  (.A1(\V3/V4/v2 [1]),
    .A2(\V3/V4/v3 [1]),
    .ZN(\V3/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M2/M1/_1_  (.A(\V3/V4/v2 [1]),
    .B(\V3/V4/v3 [1]),
    .Z(\V3/V4/A1/A1/M2/s1 ));
 AND2_X1 \V3/V4/A1/A1/M2/M2/_0_  (.A1(\V3/V4/A1/A1/M2/s1 ),
    .A2(\V3/V4/A1/A1/c1 ),
    .ZN(\V3/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M2/M2/_1_  (.A(\V3/V4/A1/A1/M2/s1 ),
    .B(\V3/V4/A1/A1/c1 ),
    .Z(\V3/V4/s1 [1]));
 OR2_X1 \V3/V4/A1/A1/M2/_0_  (.A1(\V3/V4/A1/A1/M2/c1 ),
    .A2(\V3/V4/A1/A1/M2/c2 ),
    .ZN(\V3/V4/A1/A1/c2 ));
 AND2_X1 \V3/V4/A1/A1/M3/M1/_0_  (.A1(\V3/V4/v2 [2]),
    .A2(\V3/V4/v3 [2]),
    .ZN(\V3/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M3/M1/_1_  (.A(\V3/V4/v2 [2]),
    .B(\V3/V4/v3 [2]),
    .Z(\V3/V4/A1/A1/M3/s1 ));
 AND2_X1 \V3/V4/A1/A1/M3/M2/_0_  (.A1(\V3/V4/A1/A1/M3/s1 ),
    .A2(\V3/V4/A1/A1/c2 ),
    .ZN(\V3/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M3/M2/_1_  (.A(\V3/V4/A1/A1/M3/s1 ),
    .B(\V3/V4/A1/A1/c2 ),
    .Z(\V3/V4/s1 [2]));
 OR2_X1 \V3/V4/A1/A1/M3/_0_  (.A1(\V3/V4/A1/A1/M3/c1 ),
    .A2(\V3/V4/A1/A1/M3/c2 ),
    .ZN(\V3/V4/A1/A1/c3 ));
 AND2_X1 \V3/V4/A1/A1/M4/M1/_0_  (.A1(\V3/V4/v2 [3]),
    .A2(\V3/V4/v3 [3]),
    .ZN(\V3/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A1/A1/M4/M1/_1_  (.A(\V3/V4/v2 [3]),
    .B(\V3/V4/v3 [3]),
    .Z(\V3/V4/A1/A1/M4/s1 ));
 AND2_X1 \V3/V4/A1/A1/M4/M2/_0_  (.A1(\V3/V4/A1/A1/M4/s1 ),
    .A2(\V3/V4/A1/A1/c3 ),
    .ZN(\V3/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A1/A1/M4/M2/_1_  (.A(\V3/V4/A1/A1/M4/s1 ),
    .B(\V3/V4/A1/A1/c3 ),
    .Z(\V3/V4/s1 [3]));
 OR2_X1 \V3/V4/A1/A1/M4/_0_  (.A1(\V3/V4/A1/A1/M4/c1 ),
    .A2(\V3/V4/A1/A1/M4/c2 ),
    .ZN(\V3/V4/A1/c1 ));
 AND2_X1 \V3/V4/A1/A2/M1/M1/_0_  (.A1(\V3/V4/v2 [4]),
    .A2(\V3/V4/v3 [4]),
    .ZN(\V3/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M1/M1/_1_  (.A(\V3/V4/v2 [4]),
    .B(\V3/V4/v3 [4]),
    .Z(\V3/V4/A1/A2/M1/s1 ));
 AND2_X1 \V3/V4/A1/A2/M1/M2/_0_  (.A1(\V3/V4/A1/A2/M1/s1 ),
    .A2(\V3/V4/A1/c1 ),
    .ZN(\V3/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M1/M2/_1_  (.A(\V3/V4/A1/A2/M1/s1 ),
    .B(\V3/V4/A1/c1 ),
    .Z(\V3/V4/s1 [4]));
 OR2_X1 \V3/V4/A1/A2/M1/_0_  (.A1(\V3/V4/A1/A2/M1/c1 ),
    .A2(\V3/V4/A1/A2/M1/c2 ),
    .ZN(\V3/V4/A1/A2/c1 ));
 AND2_X1 \V3/V4/A1/A2/M2/M1/_0_  (.A1(\V3/V4/v2 [5]),
    .A2(\V3/V4/v3 [5]),
    .ZN(\V3/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M2/M1/_1_  (.A(\V3/V4/v2 [5]),
    .B(\V3/V4/v3 [5]),
    .Z(\V3/V4/A1/A2/M2/s1 ));
 AND2_X1 \V3/V4/A1/A2/M2/M2/_0_  (.A1(\V3/V4/A1/A2/M2/s1 ),
    .A2(\V3/V4/A1/A2/c1 ),
    .ZN(\V3/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M2/M2/_1_  (.A(\V3/V4/A1/A2/M2/s1 ),
    .B(\V3/V4/A1/A2/c1 ),
    .Z(\V3/V4/s1 [5]));
 OR2_X1 \V3/V4/A1/A2/M2/_0_  (.A1(\V3/V4/A1/A2/M2/c1 ),
    .A2(\V3/V4/A1/A2/M2/c2 ),
    .ZN(\V3/V4/A1/A2/c2 ));
 AND2_X1 \V3/V4/A1/A2/M3/M1/_0_  (.A1(\V3/V4/v2 [6]),
    .A2(\V3/V4/v3 [6]),
    .ZN(\V3/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M3/M1/_1_  (.A(\V3/V4/v2 [6]),
    .B(\V3/V4/v3 [6]),
    .Z(\V3/V4/A1/A2/M3/s1 ));
 AND2_X1 \V3/V4/A1/A2/M3/M2/_0_  (.A1(\V3/V4/A1/A2/M3/s1 ),
    .A2(\V3/V4/A1/A2/c2 ),
    .ZN(\V3/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M3/M2/_1_  (.A(\V3/V4/A1/A2/M3/s1 ),
    .B(\V3/V4/A1/A2/c2 ),
    .Z(\V3/V4/s1 [6]));
 OR2_X1 \V3/V4/A1/A2/M3/_0_  (.A1(\V3/V4/A1/A2/M3/c1 ),
    .A2(\V3/V4/A1/A2/M3/c2 ),
    .ZN(\V3/V4/A1/A2/c3 ));
 AND2_X1 \V3/V4/A1/A2/M4/M1/_0_  (.A1(\V3/V4/v2 [7]),
    .A2(\V3/V4/v3 [7]),
    .ZN(\V3/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A1/A2/M4/M1/_1_  (.A(\V3/V4/v2 [7]),
    .B(\V3/V4/v3 [7]),
    .Z(\V3/V4/A1/A2/M4/s1 ));
 AND2_X1 \V3/V4/A1/A2/M4/M2/_0_  (.A1(\V3/V4/A1/A2/M4/s1 ),
    .A2(\V3/V4/A1/A2/c3 ),
    .ZN(\V3/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A1/A2/M4/M2/_1_  (.A(\V3/V4/A1/A2/M4/s1 ),
    .B(\V3/V4/A1/A2/c3 ),
    .Z(\V3/V4/s1 [7]));
 OR2_X1 \V3/V4/A1/A2/M4/_0_  (.A1(\V3/V4/A1/A2/M4/c1 ),
    .A2(\V3/V4/A1/A2/M4/c2 ),
    .ZN(\V3/V4/c1 ));
 AND2_X1 \V3/V4/A2/A1/M1/M1/_0_  (.A1(\V3/V4/s1 [0]),
    .A2(\V3/V4/v1 [4]),
    .ZN(\V3/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M1/M1/_1_  (.A(\V3/V4/s1 [0]),
    .B(\V3/V4/v1 [4]),
    .Z(\V3/V4/A2/A1/M1/s1 ));
 AND2_X1 \V3/V4/A2/A1/M1/M2/_0_  (.A1(\V3/V4/A2/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M1/M2/_1_  (.A(\V3/V4/A2/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/v4 [4]));
 OR2_X1 \V3/V4/A2/A1/M1/_0_  (.A1(\V3/V4/A2/A1/M1/c1 ),
    .A2(\V3/V4/A2/A1/M1/c2 ),
    .ZN(\V3/V4/A2/A1/c1 ));
 AND2_X1 \V3/V4/A2/A1/M2/M1/_0_  (.A1(\V3/V4/s1 [1]),
    .A2(\V3/V4/v1 [5]),
    .ZN(\V3/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M2/M1/_1_  (.A(\V3/V4/s1 [1]),
    .B(\V3/V4/v1 [5]),
    .Z(\V3/V4/A2/A1/M2/s1 ));
 AND2_X1 \V3/V4/A2/A1/M2/M2/_0_  (.A1(\V3/V4/A2/A1/M2/s1 ),
    .A2(\V3/V4/A2/A1/c1 ),
    .ZN(\V3/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M2/M2/_1_  (.A(\V3/V4/A2/A1/M2/s1 ),
    .B(\V3/V4/A2/A1/c1 ),
    .Z(\V3/v4 [5]));
 OR2_X1 \V3/V4/A2/A1/M2/_0_  (.A1(\V3/V4/A2/A1/M2/c1 ),
    .A2(\V3/V4/A2/A1/M2/c2 ),
    .ZN(\V3/V4/A2/A1/c2 ));
 AND2_X1 \V3/V4/A2/A1/M3/M1/_0_  (.A1(\V3/V4/s1 [2]),
    .A2(\V3/V4/v1 [6]),
    .ZN(\V3/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M3/M1/_1_  (.A(\V3/V4/s1 [2]),
    .B(\V3/V4/v1 [6]),
    .Z(\V3/V4/A2/A1/M3/s1 ));
 AND2_X1 \V3/V4/A2/A1/M3/M2/_0_  (.A1(\V3/V4/A2/A1/M3/s1 ),
    .A2(\V3/V4/A2/A1/c2 ),
    .ZN(\V3/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M3/M2/_1_  (.A(\V3/V4/A2/A1/M3/s1 ),
    .B(\V3/V4/A2/A1/c2 ),
    .Z(\V3/v4 [6]));
 OR2_X1 \V3/V4/A2/A1/M3/_0_  (.A1(\V3/V4/A2/A1/M3/c1 ),
    .A2(\V3/V4/A2/A1/M3/c2 ),
    .ZN(\V3/V4/A2/A1/c3 ));
 AND2_X1 \V3/V4/A2/A1/M4/M1/_0_  (.A1(\V3/V4/s1 [3]),
    .A2(\V3/V4/v1 [7]),
    .ZN(\V3/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A2/A1/M4/M1/_1_  (.A(\V3/V4/s1 [3]),
    .B(\V3/V4/v1 [7]),
    .Z(\V3/V4/A2/A1/M4/s1 ));
 AND2_X1 \V3/V4/A2/A1/M4/M2/_0_  (.A1(\V3/V4/A2/A1/M4/s1 ),
    .A2(\V3/V4/A2/A1/c3 ),
    .ZN(\V3/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A2/A1/M4/M2/_1_  (.A(\V3/V4/A2/A1/M4/s1 ),
    .B(\V3/V4/A2/A1/c3 ),
    .Z(\V3/v4 [7]));
 OR2_X1 \V3/V4/A2/A1/M4/_0_  (.A1(\V3/V4/A2/A1/M4/c1 ),
    .A2(\V3/V4/A2/A1/M4/c2 ),
    .ZN(\V3/V4/A2/c1 ));
 AND2_X1 \V3/V4/A2/A2/M1/M1/_0_  (.A1(\V3/V4/s1 [4]),
    .A2(net8),
    .ZN(\V3/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M1/M1/_1_  (.A(\V3/V4/s1 [4]),
    .B(net8),
    .Z(\V3/V4/A2/A2/M1/s1 ));
 AND2_X1 \V3/V4/A2/A2/M1/M2/_0_  (.A1(\V3/V4/A2/A2/M1/s1 ),
    .A2(\V3/V4/A2/c1 ),
    .ZN(\V3/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M1/M2/_1_  (.A(\V3/V4/A2/A2/M1/s1 ),
    .B(\V3/V4/A2/c1 ),
    .Z(\V3/V4/s2 [4]));
 OR2_X1 \V3/V4/A2/A2/M1/_0_  (.A1(\V3/V4/A2/A2/M1/c1 ),
    .A2(\V3/V4/A2/A2/M1/c2 ),
    .ZN(\V3/V4/A2/A2/c1 ));
 AND2_X1 \V3/V4/A2/A2/M2/M1/_0_  (.A1(\V3/V4/s1 [5]),
    .A2(net8),
    .ZN(\V3/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M2/M1/_1_  (.A(\V3/V4/s1 [5]),
    .B(net8),
    .Z(\V3/V4/A2/A2/M2/s1 ));
 AND2_X1 \V3/V4/A2/A2/M2/M2/_0_  (.A1(\V3/V4/A2/A2/M2/s1 ),
    .A2(\V3/V4/A2/A2/c1 ),
    .ZN(\V3/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M2/M2/_1_  (.A(\V3/V4/A2/A2/M2/s1 ),
    .B(\V3/V4/A2/A2/c1 ),
    .Z(\V3/V4/s2 [5]));
 OR2_X1 \V3/V4/A2/A2/M2/_0_  (.A1(\V3/V4/A2/A2/M2/c1 ),
    .A2(\V3/V4/A2/A2/M2/c2 ),
    .ZN(\V3/V4/A2/A2/c2 ));
 AND2_X1 \V3/V4/A2/A2/M3/M1/_0_  (.A1(\V3/V4/s1 [6]),
    .A2(net8),
    .ZN(\V3/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M3/M1/_1_  (.A(\V3/V4/s1 [6]),
    .B(net8),
    .Z(\V3/V4/A2/A2/M3/s1 ));
 AND2_X1 \V3/V4/A2/A2/M3/M2/_0_  (.A1(\V3/V4/A2/A2/M3/s1 ),
    .A2(\V3/V4/A2/A2/c2 ),
    .ZN(\V3/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M3/M2/_1_  (.A(\V3/V4/A2/A2/M3/s1 ),
    .B(\V3/V4/A2/A2/c2 ),
    .Z(\V3/V4/s2 [6]));
 OR2_X1 \V3/V4/A2/A2/M3/_0_  (.A1(\V3/V4/A2/A2/M3/c1 ),
    .A2(\V3/V4/A2/A2/M3/c2 ),
    .ZN(\V3/V4/A2/A2/c3 ));
 AND2_X1 \V3/V4/A2/A2/M4/M1/_0_  (.A1(\V3/V4/s1 [7]),
    .A2(net8),
    .ZN(\V3/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A2/A2/M4/M1/_1_  (.A(\V3/V4/s1 [7]),
    .B(net8),
    .Z(\V3/V4/A2/A2/M4/s1 ));
 AND2_X1 \V3/V4/A2/A2/M4/M2/_0_  (.A1(\V3/V4/A2/A2/M4/s1 ),
    .A2(\V3/V4/A2/A2/c3 ),
    .ZN(\V3/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A2/A2/M4/M2/_1_  (.A(\V3/V4/A2/A2/M4/s1 ),
    .B(\V3/V4/A2/A2/c3 ),
    .Z(\V3/V4/s2 [7]));
 OR2_X1 \V3/V4/A2/A2/M4/_0_  (.A1(\V3/V4/A2/A2/M4/c1 ),
    .A2(\V3/V4/A2/A2/M4/c2 ),
    .ZN(\V3/V4/c2 ));
 AND2_X1 \V3/V4/A3/A1/M1/M1/_0_  (.A1(\V3/V4/v4 [0]),
    .A2(\V3/V4/s2 [4]),
    .ZN(\V3/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M1/M1/_1_  (.A(\V3/V4/v4 [0]),
    .B(\V3/V4/s2 [4]),
    .Z(\V3/V4/A3/A1/M1/s1 ));
 AND2_X1 \V3/V4/A3/A1/M1/M2/_0_  (.A1(\V3/V4/A3/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M1/M2/_1_  (.A(\V3/V4/A3/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/v4 [8]));
 OR2_X1 \V3/V4/A3/A1/M1/_0_  (.A1(\V3/V4/A3/A1/M1/c1 ),
    .A2(\V3/V4/A3/A1/M1/c2 ),
    .ZN(\V3/V4/A3/A1/c1 ));
 AND2_X1 \V3/V4/A3/A1/M2/M1/_0_  (.A1(\V3/V4/v4 [1]),
    .A2(\V3/V4/s2 [5]),
    .ZN(\V3/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M2/M1/_1_  (.A(\V3/V4/v4 [1]),
    .B(\V3/V4/s2 [5]),
    .Z(\V3/V4/A3/A1/M2/s1 ));
 AND2_X1 \V3/V4/A3/A1/M2/M2/_0_  (.A1(\V3/V4/A3/A1/M2/s1 ),
    .A2(\V3/V4/A3/A1/c1 ),
    .ZN(\V3/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M2/M2/_1_  (.A(\V3/V4/A3/A1/M2/s1 ),
    .B(\V3/V4/A3/A1/c1 ),
    .Z(\V3/v4 [9]));
 OR2_X1 \V3/V4/A3/A1/M2/_0_  (.A1(\V3/V4/A3/A1/M2/c1 ),
    .A2(\V3/V4/A3/A1/M2/c2 ),
    .ZN(\V3/V4/A3/A1/c2 ));
 AND2_X1 \V3/V4/A3/A1/M3/M1/_0_  (.A1(\V3/V4/v4 [2]),
    .A2(\V3/V4/s2 [6]),
    .ZN(\V3/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M3/M1/_1_  (.A(\V3/V4/v4 [2]),
    .B(\V3/V4/s2 [6]),
    .Z(\V3/V4/A3/A1/M3/s1 ));
 AND2_X1 \V3/V4/A3/A1/M3/M2/_0_  (.A1(\V3/V4/A3/A1/M3/s1 ),
    .A2(\V3/V4/A3/A1/c2 ),
    .ZN(\V3/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M3/M2/_1_  (.A(\V3/V4/A3/A1/M3/s1 ),
    .B(\V3/V4/A3/A1/c2 ),
    .Z(\V3/v4 [10]));
 OR2_X1 \V3/V4/A3/A1/M3/_0_  (.A1(\V3/V4/A3/A1/M3/c1 ),
    .A2(\V3/V4/A3/A1/M3/c2 ),
    .ZN(\V3/V4/A3/A1/c3 ));
 AND2_X1 \V3/V4/A3/A1/M4/M1/_0_  (.A1(\V3/V4/v4 [3]),
    .A2(\V3/V4/s2 [7]),
    .ZN(\V3/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V3/V4/A3/A1/M4/M1/_1_  (.A(\V3/V4/v4 [3]),
    .B(\V3/V4/s2 [7]),
    .Z(\V3/V4/A3/A1/M4/s1 ));
 AND2_X1 \V3/V4/A3/A1/M4/M2/_0_  (.A1(\V3/V4/A3/A1/M4/s1 ),
    .A2(\V3/V4/A3/A1/c3 ),
    .ZN(\V3/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V3/V4/A3/A1/M4/M2/_1_  (.A(\V3/V4/A3/A1/M4/s1 ),
    .B(\V3/V4/A3/A1/c3 ),
    .Z(\V3/v4 [11]));
 OR2_X1 \V3/V4/A3/A1/M4/_0_  (.A1(\V3/V4/A3/A1/M4/c1 ),
    .A2(\V3/V4/A3/A1/M4/c2 ),
    .ZN(\V3/V4/A3/c1 ));
 AND2_X1 \V3/V4/A3/A2/M1/M1/_0_  (.A1(\V3/V4/v4 [4]),
    .A2(\V3/V4/c3 ),
    .ZN(\V3/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M1/M1/_1_  (.A(\V3/V4/v4 [4]),
    .B(\V3/V4/c3 ),
    .Z(\V3/V4/A3/A2/M1/s1 ));
 AND2_X1 \V3/V4/A3/A2/M1/M2/_0_  (.A1(\V3/V4/A3/A2/M1/s1 ),
    .A2(\V3/V4/A3/c1 ),
    .ZN(\V3/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M1/M2/_1_  (.A(\V3/V4/A3/A2/M1/s1 ),
    .B(\V3/V4/A3/c1 ),
    .Z(\V3/v4 [12]));
 OR2_X1 \V3/V4/A3/A2/M1/_0_  (.A1(\V3/V4/A3/A2/M1/c1 ),
    .A2(\V3/V4/A3/A2/M1/c2 ),
    .ZN(\V3/V4/A3/A2/c1 ));
 AND2_X1 \V3/V4/A3/A2/M2/M1/_0_  (.A1(\V3/V4/v4 [5]),
    .A2(net7),
    .ZN(\V3/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M2/M1/_1_  (.A(\V3/V4/v4 [5]),
    .B(net7),
    .Z(\V3/V4/A3/A2/M2/s1 ));
 AND2_X1 \V3/V4/A3/A2/M2/M2/_0_  (.A1(\V3/V4/A3/A2/M2/s1 ),
    .A2(\V3/V4/A3/A2/c1 ),
    .ZN(\V3/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M2/M2/_1_  (.A(\V3/V4/A3/A2/M2/s1 ),
    .B(\V3/V4/A3/A2/c1 ),
    .Z(\V3/v4 [13]));
 OR2_X1 \V3/V4/A3/A2/M2/_0_  (.A1(\V3/V4/A3/A2/M2/c1 ),
    .A2(\V3/V4/A3/A2/M2/c2 ),
    .ZN(\V3/V4/A3/A2/c2 ));
 AND2_X1 \V3/V4/A3/A2/M3/M1/_0_  (.A1(\V3/V4/v4 [6]),
    .A2(net7),
    .ZN(\V3/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M3/M1/_1_  (.A(\V3/V4/v4 [6]),
    .B(net7),
    .Z(\V3/V4/A3/A2/M3/s1 ));
 AND2_X1 \V3/V4/A3/A2/M3/M2/_0_  (.A1(\V3/V4/A3/A2/M3/s1 ),
    .A2(\V3/V4/A3/A2/c2 ),
    .ZN(\V3/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M3/M2/_1_  (.A(\V3/V4/A3/A2/M3/s1 ),
    .B(\V3/V4/A3/A2/c2 ),
    .Z(\V3/v4 [14]));
 OR2_X1 \V3/V4/A3/A2/M3/_0_  (.A1(\V3/V4/A3/A2/M3/c1 ),
    .A2(\V3/V4/A3/A2/M3/c2 ),
    .ZN(\V3/V4/A3/A2/c3 ));
 AND2_X1 \V3/V4/A3/A2/M4/M1/_0_  (.A1(\V3/V4/v4 [7]),
    .A2(net7),
    .ZN(\V3/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V3/V4/A3/A2/M4/M1/_1_  (.A(\V3/V4/v4 [7]),
    .B(net7),
    .Z(\V3/V4/A3/A2/M4/s1 ));
 AND2_X1 \V3/V4/A3/A2/M4/M2/_0_  (.A1(\V3/V4/A3/A2/M4/s1 ),
    .A2(\V3/V4/A3/A2/c3 ),
    .ZN(\V3/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V3/V4/A3/A2/M4/M2/_1_  (.A(\V3/V4/A3/A2/M4/s1 ),
    .B(\V3/V4/A3/A2/c3 ),
    .Z(\V3/v4 [15]));
 OR2_X1 \V3/V4/A3/A2/M4/_0_  (.A1(\V3/V4/A3/A2/M4/c1 ),
    .A2(\V3/V4/A3/A2/M4/c2 ),
    .ZN(\V3/V4/overflow ));
 AND2_X1 \V3/V4/V1/A1/M1/M1/_0_  (.A1(\V3/V4/V1/v2 [0]),
    .A2(\V3/V4/V1/v3 [0]),
    .ZN(\V3/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M1/M1/_1_  (.A(\V3/V4/V1/v2 [0]),
    .B(\V3/V4/V1/v3 [0]),
    .Z(\V3/V4/V1/A1/M1/s1 ));
 AND2_X1 \V3/V4/V1/A1/M1/M2/_0_  (.A1(\V3/V4/V1/A1/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M1/M2/_1_  (.A(\V3/V4/V1/A1/M1/s1 ),
    .B(net6),
    .Z(\V3/V4/V1/s1 [0]));
 OR2_X1 \V3/V4/V1/A1/M1/_0_  (.A1(\V3/V4/V1/A1/M1/c1 ),
    .A2(\V3/V4/V1/A1/M1/c2 ),
    .ZN(\V3/V4/V1/A1/c1 ));
 AND2_X1 \V3/V4/V1/A1/M2/M1/_0_  (.A1(\V3/V4/V1/v2 [1]),
    .A2(\V3/V4/V1/v3 [1]),
    .ZN(\V3/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M2/M1/_1_  (.A(\V3/V4/V1/v2 [1]),
    .B(\V3/V4/V1/v3 [1]),
    .Z(\V3/V4/V1/A1/M2/s1 ));
 AND2_X1 \V3/V4/V1/A1/M2/M2/_0_  (.A1(\V3/V4/V1/A1/M2/s1 ),
    .A2(\V3/V4/V1/A1/c1 ),
    .ZN(\V3/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M2/M2/_1_  (.A(\V3/V4/V1/A1/M2/s1 ),
    .B(\V3/V4/V1/A1/c1 ),
    .Z(\V3/V4/V1/s1 [1]));
 OR2_X1 \V3/V4/V1/A1/M2/_0_  (.A1(\V3/V4/V1/A1/M2/c1 ),
    .A2(\V3/V4/V1/A1/M2/c2 ),
    .ZN(\V3/V4/V1/A1/c2 ));
 AND2_X1 \V3/V4/V1/A1/M3/M1/_0_  (.A1(\V3/V4/V1/v2 [2]),
    .A2(\V3/V4/V1/v3 [2]),
    .ZN(\V3/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M3/M1/_1_  (.A(\V3/V4/V1/v2 [2]),
    .B(\V3/V4/V1/v3 [2]),
    .Z(\V3/V4/V1/A1/M3/s1 ));
 AND2_X1 \V3/V4/V1/A1/M3/M2/_0_  (.A1(\V3/V4/V1/A1/M3/s1 ),
    .A2(\V3/V4/V1/A1/c2 ),
    .ZN(\V3/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M3/M2/_1_  (.A(\V3/V4/V1/A1/M3/s1 ),
    .B(\V3/V4/V1/A1/c2 ),
    .Z(\V3/V4/V1/s1 [2]));
 OR2_X1 \V3/V4/V1/A1/M3/_0_  (.A1(\V3/V4/V1/A1/M3/c1 ),
    .A2(\V3/V4/V1/A1/M3/c2 ),
    .ZN(\V3/V4/V1/A1/c3 ));
 AND2_X1 \V3/V4/V1/A1/M4/M1/_0_  (.A1(\V3/V4/V1/v2 [3]),
    .A2(\V3/V4/V1/v3 [3]),
    .ZN(\V3/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A1/M4/M1/_1_  (.A(\V3/V4/V1/v2 [3]),
    .B(\V3/V4/V1/v3 [3]),
    .Z(\V3/V4/V1/A1/M4/s1 ));
 AND2_X1 \V3/V4/V1/A1/M4/M2/_0_  (.A1(\V3/V4/V1/A1/M4/s1 ),
    .A2(\V3/V4/V1/A1/c3 ),
    .ZN(\V3/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A1/M4/M2/_1_  (.A(\V3/V4/V1/A1/M4/s1 ),
    .B(\V3/V4/V1/A1/c3 ),
    .Z(\V3/V4/V1/s1 [3]));
 OR2_X1 \V3/V4/V1/A1/M4/_0_  (.A1(\V3/V4/V1/A1/M4/c1 ),
    .A2(\V3/V4/V1/A1/M4/c2 ),
    .ZN(\V3/V4/V1/c1 ));
 AND2_X1 \V3/V4/V1/A2/M1/M1/_0_  (.A1(\V3/V4/V1/s1 [0]),
    .A2(\V3/V4/V1/v1 [2]),
    .ZN(\V3/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M1/M1/_1_  (.A(\V3/V4/V1/s1 [0]),
    .B(\V3/V4/V1/v1 [2]),
    .Z(\V3/V4/V1/A2/M1/s1 ));
 AND2_X1 \V3/V4/V1/A2/M1/M2/_0_  (.A1(\V3/V4/V1/A2/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M1/M2/_1_  (.A(\V3/V4/V1/A2/M1/s1 ),
    .B(net6),
    .Z(\V3/v4 [2]));
 OR2_X1 \V3/V4/V1/A2/M1/_0_  (.A1(\V3/V4/V1/A2/M1/c1 ),
    .A2(\V3/V4/V1/A2/M1/c2 ),
    .ZN(\V3/V4/V1/A2/c1 ));
 AND2_X1 \V3/V4/V1/A2/M2/M1/_0_  (.A1(\V3/V4/V1/s1 [1]),
    .A2(\V3/V4/V1/v1 [3]),
    .ZN(\V3/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M2/M1/_1_  (.A(\V3/V4/V1/s1 [1]),
    .B(\V3/V4/V1/v1 [3]),
    .Z(\V3/V4/V1/A2/M2/s1 ));
 AND2_X1 \V3/V4/V1/A2/M2/M2/_0_  (.A1(\V3/V4/V1/A2/M2/s1 ),
    .A2(\V3/V4/V1/A2/c1 ),
    .ZN(\V3/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M2/M2/_1_  (.A(\V3/V4/V1/A2/M2/s1 ),
    .B(\V3/V4/V1/A2/c1 ),
    .Z(\V3/v4 [3]));
 OR2_X1 \V3/V4/V1/A2/M2/_0_  (.A1(\V3/V4/V1/A2/M2/c1 ),
    .A2(\V3/V4/V1/A2/M2/c2 ),
    .ZN(\V3/V4/V1/A2/c2 ));
 AND2_X1 \V3/V4/V1/A2/M3/M1/_0_  (.A1(\V3/V4/V1/s1 [2]),
    .A2(net6),
    .ZN(\V3/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M3/M1/_1_  (.A(\V3/V4/V1/s1 [2]),
    .B(net6),
    .Z(\V3/V4/V1/A2/M3/s1 ));
 AND2_X1 \V3/V4/V1/A2/M3/M2/_0_  (.A1(\V3/V4/V1/A2/M3/s1 ),
    .A2(\V3/V4/V1/A2/c2 ),
    .ZN(\V3/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M3/M2/_1_  (.A(\V3/V4/V1/A2/M3/s1 ),
    .B(\V3/V4/V1/A2/c2 ),
    .Z(\V3/V4/V1/s2 [2]));
 OR2_X1 \V3/V4/V1/A2/M3/_0_  (.A1(\V3/V4/V1/A2/M3/c1 ),
    .A2(\V3/V4/V1/A2/M3/c2 ),
    .ZN(\V3/V4/V1/A2/c3 ));
 AND2_X1 \V3/V4/V1/A2/M4/M1/_0_  (.A1(\V3/V4/V1/s1 [3]),
    .A2(net6),
    .ZN(\V3/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A2/M4/M1/_1_  (.A(\V3/V4/V1/s1 [3]),
    .B(net6),
    .Z(\V3/V4/V1/A2/M4/s1 ));
 AND2_X1 \V3/V4/V1/A2/M4/M2/_0_  (.A1(\V3/V4/V1/A2/M4/s1 ),
    .A2(\V3/V4/V1/A2/c3 ),
    .ZN(\V3/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A2/M4/M2/_1_  (.A(\V3/V4/V1/A2/M4/s1 ),
    .B(\V3/V4/V1/A2/c3 ),
    .Z(\V3/V4/V1/s2 [3]));
 OR2_X1 \V3/V4/V1/A2/M4/_0_  (.A1(\V3/V4/V1/A2/M4/c1 ),
    .A2(\V3/V4/V1/A2/M4/c2 ),
    .ZN(\V3/V4/V1/c2 ));
 AND2_X1 \V3/V4/V1/A3/M1/M1/_0_  (.A1(\V3/V4/V1/v4 [0]),
    .A2(\V3/V4/V1/s2 [2]),
    .ZN(\V3/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M1/M1/_1_  (.A(\V3/V4/V1/v4 [0]),
    .B(\V3/V4/V1/s2 [2]),
    .Z(\V3/V4/V1/A3/M1/s1 ));
 AND2_X1 \V3/V4/V1/A3/M1/M2/_0_  (.A1(\V3/V4/V1/A3/M1/s1 ),
    .A2(net6),
    .ZN(\V3/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M1/M2/_1_  (.A(\V3/V4/V1/A3/M1/s1 ),
    .B(net6),
    .Z(\V3/V4/v1 [4]));
 OR2_X1 \V3/V4/V1/A3/M1/_0_  (.A1(\V3/V4/V1/A3/M1/c1 ),
    .A2(\V3/V4/V1/A3/M1/c2 ),
    .ZN(\V3/V4/V1/A3/c1 ));
 AND2_X1 \V3/V4/V1/A3/M2/M1/_0_  (.A1(\V3/V4/V1/v4 [1]),
    .A2(\V3/V4/V1/s2 [3]),
    .ZN(\V3/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M2/M1/_1_  (.A(\V3/V4/V1/v4 [1]),
    .B(\V3/V4/V1/s2 [3]),
    .Z(\V3/V4/V1/A3/M2/s1 ));
 AND2_X1 \V3/V4/V1/A3/M2/M2/_0_  (.A1(\V3/V4/V1/A3/M2/s1 ),
    .A2(\V3/V4/V1/A3/c1 ),
    .ZN(\V3/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M2/M2/_1_  (.A(\V3/V4/V1/A3/M2/s1 ),
    .B(\V3/V4/V1/A3/c1 ),
    .Z(\V3/V4/v1 [5]));
 OR2_X1 \V3/V4/V1/A3/M2/_0_  (.A1(\V3/V4/V1/A3/M2/c1 ),
    .A2(\V3/V4/V1/A3/M2/c2 ),
    .ZN(\V3/V4/V1/A3/c2 ));
 AND2_X1 \V3/V4/V1/A3/M3/M1/_0_  (.A1(\V3/V4/V1/v4 [2]),
    .A2(\V3/V4/V1/c3 ),
    .ZN(\V3/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M3/M1/_1_  (.A(\V3/V4/V1/v4 [2]),
    .B(\V3/V4/V1/c3 ),
    .Z(\V3/V4/V1/A3/M3/s1 ));
 AND2_X1 \V3/V4/V1/A3/M3/M2/_0_  (.A1(\V3/V4/V1/A3/M3/s1 ),
    .A2(\V3/V4/V1/A3/c2 ),
    .ZN(\V3/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M3/M2/_1_  (.A(\V3/V4/V1/A3/M3/s1 ),
    .B(\V3/V4/V1/A3/c2 ),
    .Z(\V3/V4/v1 [6]));
 OR2_X1 \V3/V4/V1/A3/M3/_0_  (.A1(\V3/V4/V1/A3/M3/c1 ),
    .A2(\V3/V4/V1/A3/M3/c2 ),
    .ZN(\V3/V4/V1/A3/c3 ));
 AND2_X1 \V3/V4/V1/A3/M4/M1/_0_  (.A1(\V3/V4/V1/v4 [3]),
    .A2(net6),
    .ZN(\V3/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V1/A3/M4/M1/_1_  (.A(\V3/V4/V1/v4 [3]),
    .B(net6),
    .Z(\V3/V4/V1/A3/M4/s1 ));
 AND2_X1 \V3/V4/V1/A3/M4/M2/_0_  (.A1(\V3/V4/V1/A3/M4/s1 ),
    .A2(\V3/V4/V1/A3/c3 ),
    .ZN(\V3/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V1/A3/M4/M2/_1_  (.A(\V3/V4/V1/A3/M4/s1 ),
    .B(\V3/V4/V1/A3/c3 ),
    .Z(\V3/V4/v1 [7]));
 OR2_X1 \V3/V4/V1/A3/M4/_0_  (.A1(\V3/V4/V1/A3/M4/c1 ),
    .A2(\V3/V4/V1/A3/M4/c2 ),
    .ZN(\V3/V4/V1/overflow ));
 AND2_X1 \V3/V4/V1/V1/HA1/_0_  (.A1(\V3/V4/V1/V1/w2 ),
    .A2(\V3/V4/V1/V1/w1 ),
    .ZN(\V3/V4/V1/V1/w4 ));
 XOR2_X2 \V3/V4/V1/V1/HA1/_1_  (.A(\V3/V4/V1/V1/w2 ),
    .B(\V3/V4/V1/V1/w1 ),
    .Z(\V3/v4 [1]));
 AND2_X1 \V3/V4/V1/V1/HA2/_0_  (.A1(\V3/V4/V1/V1/w4 ),
    .A2(\V3/V4/V1/V1/w3 ),
    .ZN(\V3/V4/V1/v1 [3]));
 XOR2_X2 \V3/V4/V1/V1/HA2/_1_  (.A(\V3/V4/V1/V1/w4 ),
    .B(\V3/V4/V1/V1/w3 ),
    .Z(\V3/V4/V1/v1 [2]));
 AND2_X1 \V3/V4/V1/V1/_0_  (.A1(net25),
    .A2(net14),
    .ZN(\V3/v4 [0]));
 AND2_X1 \V3/V4/V1/V1/_1_  (.A1(net25),
    .A2(B[25]),
    .ZN(\V3/V4/V1/V1/w1 ));
 AND2_X1 \V3/V4/V1/V1/_2_  (.A1(net14),
    .A2(net24),
    .ZN(\V3/V4/V1/V1/w2 ));
 AND2_X1 \V3/V4/V1/V1/_3_  (.A1(B[25]),
    .A2(net24),
    .ZN(\V3/V4/V1/V1/w3 ));
 AND2_X1 \V3/V4/V1/V2/HA1/_0_  (.A1(\V3/V4/V1/V2/w2 ),
    .A2(\V3/V4/V1/V2/w1 ),
    .ZN(\V3/V4/V1/V2/w4 ));
 XOR2_X2 \V3/V4/V1/V2/HA1/_1_  (.A(\V3/V4/V1/V2/w2 ),
    .B(\V3/V4/V1/V2/w1 ),
    .Z(\V3/V4/V1/v2 [1]));
 AND2_X1 \V3/V4/V1/V2/HA2/_0_  (.A1(\V3/V4/V1/V2/w4 ),
    .A2(\V3/V4/V1/V2/w3 ),
    .ZN(\V3/V4/V1/v2 [3]));
 XOR2_X2 \V3/V4/V1/V2/HA2/_1_  (.A(\V3/V4/V1/V2/w4 ),
    .B(\V3/V4/V1/V2/w3 ),
    .Z(\V3/V4/V1/v2 [2]));
 AND2_X1 \V3/V4/V1/V2/_0_  (.A1(net47),
    .A2(net14),
    .ZN(\V3/V4/V1/v2 [0]));
 AND2_X1 \V3/V4/V1/V2/_1_  (.A1(net47),
    .A2(B[25]),
    .ZN(\V3/V4/V1/V2/w1 ));
 AND2_X1 \V3/V4/V1/V2/_2_  (.A1(net14),
    .A2(net46),
    .ZN(\V3/V4/V1/V2/w2 ));
 AND2_X1 \V3/V4/V1/V2/_3_  (.A1(B[25]),
    .A2(net46),
    .ZN(\V3/V4/V1/V2/w3 ));
 AND2_X1 \V3/V4/V1/V3/HA1/_0_  (.A1(\V3/V4/V1/V3/w2 ),
    .A2(\V3/V4/V1/V3/w1 ),
    .ZN(\V3/V4/V1/V3/w4 ));
 XOR2_X2 \V3/V4/V1/V3/HA1/_1_  (.A(\V3/V4/V1/V3/w2 ),
    .B(\V3/V4/V1/V3/w1 ),
    .Z(\V3/V4/V1/v3 [1]));
 AND2_X1 \V3/V4/V1/V3/HA2/_0_  (.A1(\V3/V4/V1/V3/w4 ),
    .A2(\V3/V4/V1/V3/w3 ),
    .ZN(\V3/V4/V1/v3 [3]));
 XOR2_X2 \V3/V4/V1/V3/HA2/_1_  (.A(\V3/V4/V1/V3/w4 ),
    .B(\V3/V4/V1/V3/w3 ),
    .Z(\V3/V4/V1/v3 [2]));
 AND2_X1 \V3/V4/V1/V3/_0_  (.A1(net25),
    .A2(net13),
    .ZN(\V3/V4/V1/v3 [0]));
 AND2_X1 \V3/V4/V1/V3/_1_  (.A1(net25),
    .A2(B[27]),
    .ZN(\V3/V4/V1/V3/w1 ));
 AND2_X1 \V3/V4/V1/V3/_2_  (.A1(net13),
    .A2(net24),
    .ZN(\V3/V4/V1/V3/w2 ));
 AND2_X1 \V3/V4/V1/V3/_3_  (.A1(B[27]),
    .A2(net24),
    .ZN(\V3/V4/V1/V3/w3 ));
 AND2_X1 \V3/V4/V1/V4/HA1/_0_  (.A1(\V3/V4/V1/V4/w2 ),
    .A2(\V3/V4/V1/V4/w1 ),
    .ZN(\V3/V4/V1/V4/w4 ));
 XOR2_X2 \V3/V4/V1/V4/HA1/_1_  (.A(\V3/V4/V1/V4/w2 ),
    .B(\V3/V4/V1/V4/w1 ),
    .Z(\V3/V4/V1/v4 [1]));
 AND2_X1 \V3/V4/V1/V4/HA2/_0_  (.A1(\V3/V4/V1/V4/w4 ),
    .A2(\V3/V4/V1/V4/w3 ),
    .ZN(\V3/V4/V1/v4 [3]));
 XOR2_X2 \V3/V4/V1/V4/HA2/_1_  (.A(\V3/V4/V1/V4/w4 ),
    .B(\V3/V4/V1/V4/w3 ),
    .Z(\V3/V4/V1/v4 [2]));
 AND2_X1 \V3/V4/V1/V4/_0_  (.A1(net47),
    .A2(net13),
    .ZN(\V3/V4/V1/v4 [0]));
 AND2_X1 \V3/V4/V1/V4/_1_  (.A1(net47),
    .A2(B[27]),
    .ZN(\V3/V4/V1/V4/w1 ));
 AND2_X1 \V3/V4/V1/V4/_2_  (.A1(net13),
    .A2(net46),
    .ZN(\V3/V4/V1/V4/w2 ));
 AND2_X1 \V3/V4/V1/V4/_3_  (.A1(B[27]),
    .A2(net46),
    .ZN(\V3/V4/V1/V4/w3 ));
 OR2_X1 \V3/V4/V1/_0_  (.A1(\V3/V4/V1/c1 ),
    .A2(\V3/V4/V1/c2 ),
    .ZN(\V3/V4/V1/c3 ));
 AND2_X1 \V3/V4/V2/A1/M1/M1/_0_  (.A1(\V3/V4/V2/v2 [0]),
    .A2(\V3/V4/V2/v3 [0]),
    .ZN(\V3/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M1/M1/_1_  (.A(\V3/V4/V2/v2 [0]),
    .B(\V3/V4/V2/v3 [0]),
    .Z(\V3/V4/V2/A1/M1/s1 ));
 AND2_X1 \V3/V4/V2/A1/M1/M2/_0_  (.A1(\V3/V4/V2/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M1/M2/_1_  (.A(\V3/V4/V2/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/V2/s1 [0]));
 OR2_X1 \V3/V4/V2/A1/M1/_0_  (.A1(\V3/V4/V2/A1/M1/c1 ),
    .A2(\V3/V4/V2/A1/M1/c2 ),
    .ZN(\V3/V4/V2/A1/c1 ));
 AND2_X1 \V3/V4/V2/A1/M2/M1/_0_  (.A1(\V3/V4/V2/v2 [1]),
    .A2(\V3/V4/V2/v3 [1]),
    .ZN(\V3/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M2/M1/_1_  (.A(\V3/V4/V2/v2 [1]),
    .B(\V3/V4/V2/v3 [1]),
    .Z(\V3/V4/V2/A1/M2/s1 ));
 AND2_X1 \V3/V4/V2/A1/M2/M2/_0_  (.A1(\V3/V4/V2/A1/M2/s1 ),
    .A2(\V3/V4/V2/A1/c1 ),
    .ZN(\V3/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M2/M2/_1_  (.A(\V3/V4/V2/A1/M2/s1 ),
    .B(\V3/V4/V2/A1/c1 ),
    .Z(\V3/V4/V2/s1 [1]));
 OR2_X1 \V3/V4/V2/A1/M2/_0_  (.A1(\V3/V4/V2/A1/M2/c1 ),
    .A2(\V3/V4/V2/A1/M2/c2 ),
    .ZN(\V3/V4/V2/A1/c2 ));
 AND2_X1 \V3/V4/V2/A1/M3/M1/_0_  (.A1(\V3/V4/V2/v2 [2]),
    .A2(\V3/V4/V2/v3 [2]),
    .ZN(\V3/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M3/M1/_1_  (.A(\V3/V4/V2/v2 [2]),
    .B(\V3/V4/V2/v3 [2]),
    .Z(\V3/V4/V2/A1/M3/s1 ));
 AND2_X1 \V3/V4/V2/A1/M3/M2/_0_  (.A1(\V3/V4/V2/A1/M3/s1 ),
    .A2(\V3/V4/V2/A1/c2 ),
    .ZN(\V3/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M3/M2/_1_  (.A(\V3/V4/V2/A1/M3/s1 ),
    .B(\V3/V4/V2/A1/c2 ),
    .Z(\V3/V4/V2/s1 [2]));
 OR2_X1 \V3/V4/V2/A1/M3/_0_  (.A1(\V3/V4/V2/A1/M3/c1 ),
    .A2(\V3/V4/V2/A1/M3/c2 ),
    .ZN(\V3/V4/V2/A1/c3 ));
 AND2_X1 \V3/V4/V2/A1/M4/M1/_0_  (.A1(\V3/V4/V2/v2 [3]),
    .A2(\V3/V4/V2/v3 [3]),
    .ZN(\V3/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A1/M4/M1/_1_  (.A(\V3/V4/V2/v2 [3]),
    .B(\V3/V4/V2/v3 [3]),
    .Z(\V3/V4/V2/A1/M4/s1 ));
 AND2_X1 \V3/V4/V2/A1/M4/M2/_0_  (.A1(\V3/V4/V2/A1/M4/s1 ),
    .A2(\V3/V4/V2/A1/c3 ),
    .ZN(\V3/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A1/M4/M2/_1_  (.A(\V3/V4/V2/A1/M4/s1 ),
    .B(\V3/V4/V2/A1/c3 ),
    .Z(\V3/V4/V2/s1 [3]));
 OR2_X1 \V3/V4/V2/A1/M4/_0_  (.A1(\V3/V4/V2/A1/M4/c1 ),
    .A2(\V3/V4/V2/A1/M4/c2 ),
    .ZN(\V3/V4/V2/c1 ));
 AND2_X1 \V3/V4/V2/A2/M1/M1/_0_  (.A1(\V3/V4/V2/s1 [0]),
    .A2(\V3/V4/V2/v1 [2]),
    .ZN(\V3/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M1/M1/_1_  (.A(\V3/V4/V2/s1 [0]),
    .B(\V3/V4/V2/v1 [2]),
    .Z(\V3/V4/V2/A2/M1/s1 ));
 AND2_X1 \V3/V4/V2/A2/M1/M2/_0_  (.A1(\V3/V4/V2/A2/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M1/M2/_1_  (.A(\V3/V4/V2/A2/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/v2 [2]));
 OR2_X1 \V3/V4/V2/A2/M1/_0_  (.A1(\V3/V4/V2/A2/M1/c1 ),
    .A2(\V3/V4/V2/A2/M1/c2 ),
    .ZN(\V3/V4/V2/A2/c1 ));
 AND2_X1 \V3/V4/V2/A2/M2/M1/_0_  (.A1(\V3/V4/V2/s1 [1]),
    .A2(\V3/V4/V2/v1 [3]),
    .ZN(\V3/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M2/M1/_1_  (.A(\V3/V4/V2/s1 [1]),
    .B(\V3/V4/V2/v1 [3]),
    .Z(\V3/V4/V2/A2/M2/s1 ));
 AND2_X1 \V3/V4/V2/A2/M2/M2/_0_  (.A1(\V3/V4/V2/A2/M2/s1 ),
    .A2(\V3/V4/V2/A2/c1 ),
    .ZN(\V3/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M2/M2/_1_  (.A(\V3/V4/V2/A2/M2/s1 ),
    .B(\V3/V4/V2/A2/c1 ),
    .Z(\V3/V4/v2 [3]));
 OR2_X1 \V3/V4/V2/A2/M2/_0_  (.A1(\V3/V4/V2/A2/M2/c1 ),
    .A2(\V3/V4/V2/A2/M2/c2 ),
    .ZN(\V3/V4/V2/A2/c2 ));
 AND2_X1 \V3/V4/V2/A2/M3/M1/_0_  (.A1(\V3/V4/V2/s1 [2]),
    .A2(net8),
    .ZN(\V3/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M3/M1/_1_  (.A(\V3/V4/V2/s1 [2]),
    .B(net8),
    .Z(\V3/V4/V2/A2/M3/s1 ));
 AND2_X1 \V3/V4/V2/A2/M3/M2/_0_  (.A1(\V3/V4/V2/A2/M3/s1 ),
    .A2(\V3/V4/V2/A2/c2 ),
    .ZN(\V3/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M3/M2/_1_  (.A(\V3/V4/V2/A2/M3/s1 ),
    .B(\V3/V4/V2/A2/c2 ),
    .Z(\V3/V4/V2/s2 [2]));
 OR2_X1 \V3/V4/V2/A2/M3/_0_  (.A1(\V3/V4/V2/A2/M3/c1 ),
    .A2(\V3/V4/V2/A2/M3/c2 ),
    .ZN(\V3/V4/V2/A2/c3 ));
 AND2_X1 \V3/V4/V2/A2/M4/M1/_0_  (.A1(\V3/V4/V2/s1 [3]),
    .A2(net8),
    .ZN(\V3/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A2/M4/M1/_1_  (.A(\V3/V4/V2/s1 [3]),
    .B(net8),
    .Z(\V3/V4/V2/A2/M4/s1 ));
 AND2_X1 \V3/V4/V2/A2/M4/M2/_0_  (.A1(\V3/V4/V2/A2/M4/s1 ),
    .A2(\V3/V4/V2/A2/c3 ),
    .ZN(\V3/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A2/M4/M2/_1_  (.A(\V3/V4/V2/A2/M4/s1 ),
    .B(\V3/V4/V2/A2/c3 ),
    .Z(\V3/V4/V2/s2 [3]));
 OR2_X1 \V3/V4/V2/A2/M4/_0_  (.A1(\V3/V4/V2/A2/M4/c1 ),
    .A2(\V3/V4/V2/A2/M4/c2 ),
    .ZN(\V3/V4/V2/c2 ));
 AND2_X1 \V3/V4/V2/A3/M1/M1/_0_  (.A1(\V3/V4/V2/v4 [0]),
    .A2(\V3/V4/V2/s2 [2]),
    .ZN(\V3/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M1/M1/_1_  (.A(\V3/V4/V2/v4 [0]),
    .B(\V3/V4/V2/s2 [2]),
    .Z(\V3/V4/V2/A3/M1/s1 ));
 AND2_X1 \V3/V4/V2/A3/M1/M2/_0_  (.A1(\V3/V4/V2/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M1/M2/_1_  (.A(\V3/V4/V2/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/v2 [4]));
 OR2_X1 \V3/V4/V2/A3/M1/_0_  (.A1(\V3/V4/V2/A3/M1/c1 ),
    .A2(\V3/V4/V2/A3/M1/c2 ),
    .ZN(\V3/V4/V2/A3/c1 ));
 AND2_X1 \V3/V4/V2/A3/M2/M1/_0_  (.A1(\V3/V4/V2/v4 [1]),
    .A2(\V3/V4/V2/s2 [3]),
    .ZN(\V3/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M2/M1/_1_  (.A(\V3/V4/V2/v4 [1]),
    .B(\V3/V4/V2/s2 [3]),
    .Z(\V3/V4/V2/A3/M2/s1 ));
 AND2_X1 \V3/V4/V2/A3/M2/M2/_0_  (.A1(\V3/V4/V2/A3/M2/s1 ),
    .A2(\V3/V4/V2/A3/c1 ),
    .ZN(\V3/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M2/M2/_1_  (.A(\V3/V4/V2/A3/M2/s1 ),
    .B(\V3/V4/V2/A3/c1 ),
    .Z(\V3/V4/v2 [5]));
 OR2_X1 \V3/V4/V2/A3/M2/_0_  (.A1(\V3/V4/V2/A3/M2/c1 ),
    .A2(\V3/V4/V2/A3/M2/c2 ),
    .ZN(\V3/V4/V2/A3/c2 ));
 AND2_X1 \V3/V4/V2/A3/M3/M1/_0_  (.A1(\V3/V4/V2/v4 [2]),
    .A2(\V3/V4/V2/c3 ),
    .ZN(\V3/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M3/M1/_1_  (.A(\V3/V4/V2/v4 [2]),
    .B(\V3/V4/V2/c3 ),
    .Z(\V3/V4/V2/A3/M3/s1 ));
 AND2_X1 \V3/V4/V2/A3/M3/M2/_0_  (.A1(\V3/V4/V2/A3/M3/s1 ),
    .A2(\V3/V4/V2/A3/c2 ),
    .ZN(\V3/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M3/M2/_1_  (.A(\V3/V4/V2/A3/M3/s1 ),
    .B(\V3/V4/V2/A3/c2 ),
    .Z(\V3/V4/v2 [6]));
 OR2_X1 \V3/V4/V2/A3/M3/_0_  (.A1(\V3/V4/V2/A3/M3/c1 ),
    .A2(\V3/V4/V2/A3/M3/c2 ),
    .ZN(\V3/V4/V2/A3/c3 ));
 AND2_X1 \V3/V4/V2/A3/M4/M1/_0_  (.A1(\V3/V4/V2/v4 [3]),
    .A2(net8),
    .ZN(\V3/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V2/A3/M4/M1/_1_  (.A(\V3/V4/V2/v4 [3]),
    .B(net8),
    .Z(\V3/V4/V2/A3/M4/s1 ));
 AND2_X1 \V3/V4/V2/A3/M4/M2/_0_  (.A1(\V3/V4/V2/A3/M4/s1 ),
    .A2(\V3/V4/V2/A3/c3 ),
    .ZN(\V3/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V2/A3/M4/M2/_1_  (.A(\V3/V4/V2/A3/M4/s1 ),
    .B(\V3/V4/V2/A3/c3 ),
    .Z(\V3/V4/v2 [7]));
 OR2_X1 \V3/V4/V2/A3/M4/_0_  (.A1(\V3/V4/V2/A3/M4/c1 ),
    .A2(\V3/V4/V2/A3/M4/c2 ),
    .ZN(\V3/V4/V2/overflow ));
 AND2_X1 \V3/V4/V2/V1/HA1/_0_  (.A1(\V3/V4/V2/V1/w2 ),
    .A2(\V3/V4/V2/V1/w1 ),
    .ZN(\V3/V4/V2/V1/w4 ));
 XOR2_X2 \V3/V4/V2/V1/HA1/_1_  (.A(\V3/V4/V2/V1/w2 ),
    .B(\V3/V4/V2/V1/w1 ),
    .Z(\V3/V4/v2 [1]));
 AND2_X1 \V3/V4/V2/V1/HA2/_0_  (.A1(\V3/V4/V2/V1/w4 ),
    .A2(\V3/V4/V2/V1/w3 ),
    .ZN(\V3/V4/V2/v1 [3]));
 XOR2_X2 \V3/V4/V2/V1/HA2/_1_  (.A(\V3/V4/V2/V1/w4 ),
    .B(\V3/V4/V2/V1/w3 ),
    .Z(\V3/V4/V2/v1 [2]));
 AND2_X1 \V3/V4/V2/V1/_0_  (.A1(net45),
    .A2(net14),
    .ZN(\V3/V4/v2 [0]));
 AND2_X1 \V3/V4/V2/V1/_1_  (.A1(net45),
    .A2(B[25]),
    .ZN(\V3/V4/V2/V1/w1 ));
 AND2_X1 \V3/V4/V2/V1/_2_  (.A1(net14),
    .A2(net44),
    .ZN(\V3/V4/V2/V1/w2 ));
 AND2_X1 \V3/V4/V2/V1/_3_  (.A1(B[25]),
    .A2(net44),
    .ZN(\V3/V4/V2/V1/w3 ));
 AND2_X1 \V3/V4/V2/V2/HA1/_0_  (.A1(\V3/V4/V2/V2/w2 ),
    .A2(\V3/V4/V2/V2/w1 ),
    .ZN(\V3/V4/V2/V2/w4 ));
 XOR2_X2 \V3/V4/V2/V2/HA1/_1_  (.A(\V3/V4/V2/V2/w2 ),
    .B(\V3/V4/V2/V2/w1 ),
    .Z(\V3/V4/V2/v2 [1]));
 AND2_X1 \V3/V4/V2/V2/HA2/_0_  (.A1(\V3/V4/V2/V2/w4 ),
    .A2(\V3/V4/V2/V2/w3 ),
    .ZN(\V3/V4/V2/v2 [3]));
 XOR2_X2 \V3/V4/V2/V2/HA2/_1_  (.A(\V3/V4/V2/V2/w4 ),
    .B(\V3/V4/V2/V2/w3 ),
    .Z(\V3/V4/V2/v2 [2]));
 AND2_X1 \V3/V4/V2/V2/_0_  (.A1(net43),
    .A2(net14),
    .ZN(\V3/V4/V2/v2 [0]));
 AND2_X1 \V3/V4/V2/V2/_1_  (.A1(net43),
    .A2(B[25]),
    .ZN(\V3/V4/V2/V2/w1 ));
 AND2_X1 \V3/V4/V2/V2/_2_  (.A1(net14),
    .A2(net42),
    .ZN(\V3/V4/V2/V2/w2 ));
 AND2_X1 \V3/V4/V2/V2/_3_  (.A1(B[25]),
    .A2(net42),
    .ZN(\V3/V4/V2/V2/w3 ));
 AND2_X1 \V3/V4/V2/V3/HA1/_0_  (.A1(\V3/V4/V2/V3/w2 ),
    .A2(\V3/V4/V2/V3/w1 ),
    .ZN(\V3/V4/V2/V3/w4 ));
 XOR2_X2 \V3/V4/V2/V3/HA1/_1_  (.A(\V3/V4/V2/V3/w2 ),
    .B(\V3/V4/V2/V3/w1 ),
    .Z(\V3/V4/V2/v3 [1]));
 AND2_X1 \V3/V4/V2/V3/HA2/_0_  (.A1(\V3/V4/V2/V3/w4 ),
    .A2(\V3/V4/V2/V3/w3 ),
    .ZN(\V3/V4/V2/v3 [3]));
 XOR2_X2 \V3/V4/V2/V3/HA2/_1_  (.A(\V3/V4/V2/V3/w4 ),
    .B(\V3/V4/V2/V3/w3 ),
    .Z(\V3/V4/V2/v3 [2]));
 AND2_X1 \V3/V4/V2/V3/_0_  (.A1(net45),
    .A2(net13),
    .ZN(\V3/V4/V2/v3 [0]));
 AND2_X1 \V3/V4/V2/V3/_1_  (.A1(net45),
    .A2(B[27]),
    .ZN(\V3/V4/V2/V3/w1 ));
 AND2_X1 \V3/V4/V2/V3/_2_  (.A1(net13),
    .A2(net44),
    .ZN(\V3/V4/V2/V3/w2 ));
 AND2_X1 \V3/V4/V2/V3/_3_  (.A1(B[27]),
    .A2(net44),
    .ZN(\V3/V4/V2/V3/w3 ));
 AND2_X1 \V3/V4/V2/V4/HA1/_0_  (.A1(\V3/V4/V2/V4/w2 ),
    .A2(\V3/V4/V2/V4/w1 ),
    .ZN(\V3/V4/V2/V4/w4 ));
 XOR2_X2 \V3/V4/V2/V4/HA1/_1_  (.A(\V3/V4/V2/V4/w2 ),
    .B(\V3/V4/V2/V4/w1 ),
    .Z(\V3/V4/V2/v4 [1]));
 AND2_X1 \V3/V4/V2/V4/HA2/_0_  (.A1(\V3/V4/V2/V4/w4 ),
    .A2(\V3/V4/V2/V4/w3 ),
    .ZN(\V3/V4/V2/v4 [3]));
 XOR2_X2 \V3/V4/V2/V4/HA2/_1_  (.A(\V3/V4/V2/V4/w4 ),
    .B(\V3/V4/V2/V4/w3 ),
    .Z(\V3/V4/V2/v4 [2]));
 AND2_X1 \V3/V4/V2/V4/_0_  (.A1(net43),
    .A2(net13),
    .ZN(\V3/V4/V2/v4 [0]));
 AND2_X1 \V3/V4/V2/V4/_1_  (.A1(net43),
    .A2(B[27]),
    .ZN(\V3/V4/V2/V4/w1 ));
 AND2_X1 \V3/V4/V2/V4/_2_  (.A1(net13),
    .A2(net42),
    .ZN(\V3/V4/V2/V4/w2 ));
 AND2_X1 \V3/V4/V2/V4/_3_  (.A1(B[27]),
    .A2(net42),
    .ZN(\V3/V4/V2/V4/w3 ));
 OR2_X1 \V3/V4/V2/_0_  (.A1(\V3/V4/V2/c1 ),
    .A2(\V3/V4/V2/c2 ),
    .ZN(\V3/V4/V2/c3 ));
 AND2_X1 \V3/V4/V3/A1/M1/M1/_0_  (.A1(\V3/V4/V3/v2 [0]),
    .A2(\V3/V4/V3/v3 [0]),
    .ZN(\V3/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M1/M1/_1_  (.A(\V3/V4/V3/v2 [0]),
    .B(\V3/V4/V3/v3 [0]),
    .Z(\V3/V4/V3/A1/M1/s1 ));
 AND2_X1 \V3/V4/V3/A1/M1/M2/_0_  (.A1(\V3/V4/V3/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M1/M2/_1_  (.A(\V3/V4/V3/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/V3/s1 [0]));
 OR2_X1 \V3/V4/V3/A1/M1/_0_  (.A1(\V3/V4/V3/A1/M1/c1 ),
    .A2(\V3/V4/V3/A1/M1/c2 ),
    .ZN(\V3/V4/V3/A1/c1 ));
 AND2_X1 \V3/V4/V3/A1/M2/M1/_0_  (.A1(\V3/V4/V3/v2 [1]),
    .A2(\V3/V4/V3/v3 [1]),
    .ZN(\V3/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M2/M1/_1_  (.A(\V3/V4/V3/v2 [1]),
    .B(\V3/V4/V3/v3 [1]),
    .Z(\V3/V4/V3/A1/M2/s1 ));
 AND2_X1 \V3/V4/V3/A1/M2/M2/_0_  (.A1(\V3/V4/V3/A1/M2/s1 ),
    .A2(\V3/V4/V3/A1/c1 ),
    .ZN(\V3/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M2/M2/_1_  (.A(\V3/V4/V3/A1/M2/s1 ),
    .B(\V3/V4/V3/A1/c1 ),
    .Z(\V3/V4/V3/s1 [1]));
 OR2_X1 \V3/V4/V3/A1/M2/_0_  (.A1(\V3/V4/V3/A1/M2/c1 ),
    .A2(\V3/V4/V3/A1/M2/c2 ),
    .ZN(\V3/V4/V3/A1/c2 ));
 AND2_X1 \V3/V4/V3/A1/M3/M1/_0_  (.A1(\V3/V4/V3/v2 [2]),
    .A2(\V3/V4/V3/v3 [2]),
    .ZN(\V3/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M3/M1/_1_  (.A(\V3/V4/V3/v2 [2]),
    .B(\V3/V4/V3/v3 [2]),
    .Z(\V3/V4/V3/A1/M3/s1 ));
 AND2_X1 \V3/V4/V3/A1/M3/M2/_0_  (.A1(\V3/V4/V3/A1/M3/s1 ),
    .A2(\V3/V4/V3/A1/c2 ),
    .ZN(\V3/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M3/M2/_1_  (.A(\V3/V4/V3/A1/M3/s1 ),
    .B(\V3/V4/V3/A1/c2 ),
    .Z(\V3/V4/V3/s1 [2]));
 OR2_X1 \V3/V4/V3/A1/M3/_0_  (.A1(\V3/V4/V3/A1/M3/c1 ),
    .A2(\V3/V4/V3/A1/M3/c2 ),
    .ZN(\V3/V4/V3/A1/c3 ));
 AND2_X1 \V3/V4/V3/A1/M4/M1/_0_  (.A1(\V3/V4/V3/v2 [3]),
    .A2(\V3/V4/V3/v3 [3]),
    .ZN(\V3/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A1/M4/M1/_1_  (.A(\V3/V4/V3/v2 [3]),
    .B(\V3/V4/V3/v3 [3]),
    .Z(\V3/V4/V3/A1/M4/s1 ));
 AND2_X1 \V3/V4/V3/A1/M4/M2/_0_  (.A1(\V3/V4/V3/A1/M4/s1 ),
    .A2(\V3/V4/V3/A1/c3 ),
    .ZN(\V3/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A1/M4/M2/_1_  (.A(\V3/V4/V3/A1/M4/s1 ),
    .B(\V3/V4/V3/A1/c3 ),
    .Z(\V3/V4/V3/s1 [3]));
 OR2_X1 \V3/V4/V3/A1/M4/_0_  (.A1(\V3/V4/V3/A1/M4/c1 ),
    .A2(\V3/V4/V3/A1/M4/c2 ),
    .ZN(\V3/V4/V3/c1 ));
 AND2_X1 \V3/V4/V3/A2/M1/M1/_0_  (.A1(\V3/V4/V3/s1 [0]),
    .A2(\V3/V4/V3/v1 [2]),
    .ZN(\V3/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M1/M1/_1_  (.A(\V3/V4/V3/s1 [0]),
    .B(\V3/V4/V3/v1 [2]),
    .Z(\V3/V4/V3/A2/M1/s1 ));
 AND2_X1 \V3/V4/V3/A2/M1/M2/_0_  (.A1(\V3/V4/V3/A2/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M1/M2/_1_  (.A(\V3/V4/V3/A2/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/v3 [2]));
 OR2_X1 \V3/V4/V3/A2/M1/_0_  (.A1(\V3/V4/V3/A2/M1/c1 ),
    .A2(\V3/V4/V3/A2/M1/c2 ),
    .ZN(\V3/V4/V3/A2/c1 ));
 AND2_X1 \V3/V4/V3/A2/M2/M1/_0_  (.A1(\V3/V4/V3/s1 [1]),
    .A2(\V3/V4/V3/v1 [3]),
    .ZN(\V3/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M2/M1/_1_  (.A(\V3/V4/V3/s1 [1]),
    .B(\V3/V4/V3/v1 [3]),
    .Z(\V3/V4/V3/A2/M2/s1 ));
 AND2_X1 \V3/V4/V3/A2/M2/M2/_0_  (.A1(\V3/V4/V3/A2/M2/s1 ),
    .A2(\V3/V4/V3/A2/c1 ),
    .ZN(\V3/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M2/M2/_1_  (.A(\V3/V4/V3/A2/M2/s1 ),
    .B(\V3/V4/V3/A2/c1 ),
    .Z(\V3/V4/v3 [3]));
 OR2_X1 \V3/V4/V3/A2/M2/_0_  (.A1(\V3/V4/V3/A2/M2/c1 ),
    .A2(\V3/V4/V3/A2/M2/c2 ),
    .ZN(\V3/V4/V3/A2/c2 ));
 AND2_X1 \V3/V4/V3/A2/M3/M1/_0_  (.A1(\V3/V4/V3/s1 [2]),
    .A2(net8),
    .ZN(\V3/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M3/M1/_1_  (.A(\V3/V4/V3/s1 [2]),
    .B(net8),
    .Z(\V3/V4/V3/A2/M3/s1 ));
 AND2_X1 \V3/V4/V3/A2/M3/M2/_0_  (.A1(\V3/V4/V3/A2/M3/s1 ),
    .A2(\V3/V4/V3/A2/c2 ),
    .ZN(\V3/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M3/M2/_1_  (.A(\V3/V4/V3/A2/M3/s1 ),
    .B(\V3/V4/V3/A2/c2 ),
    .Z(\V3/V4/V3/s2 [2]));
 OR2_X1 \V3/V4/V3/A2/M3/_0_  (.A1(\V3/V4/V3/A2/M3/c1 ),
    .A2(\V3/V4/V3/A2/M3/c2 ),
    .ZN(\V3/V4/V3/A2/c3 ));
 AND2_X1 \V3/V4/V3/A2/M4/M1/_0_  (.A1(\V3/V4/V3/s1 [3]),
    .A2(net8),
    .ZN(\V3/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A2/M4/M1/_1_  (.A(\V3/V4/V3/s1 [3]),
    .B(net8),
    .Z(\V3/V4/V3/A2/M4/s1 ));
 AND2_X1 \V3/V4/V3/A2/M4/M2/_0_  (.A1(\V3/V4/V3/A2/M4/s1 ),
    .A2(\V3/V4/V3/A2/c3 ),
    .ZN(\V3/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A2/M4/M2/_1_  (.A(\V3/V4/V3/A2/M4/s1 ),
    .B(\V3/V4/V3/A2/c3 ),
    .Z(\V3/V4/V3/s2 [3]));
 OR2_X1 \V3/V4/V3/A2/M4/_0_  (.A1(\V3/V4/V3/A2/M4/c1 ),
    .A2(\V3/V4/V3/A2/M4/c2 ),
    .ZN(\V3/V4/V3/c2 ));
 AND2_X1 \V3/V4/V3/A3/M1/M1/_0_  (.A1(\V3/V4/V3/v4 [0]),
    .A2(\V3/V4/V3/s2 [2]),
    .ZN(\V3/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M1/M1/_1_  (.A(\V3/V4/V3/v4 [0]),
    .B(\V3/V4/V3/s2 [2]),
    .Z(\V3/V4/V3/A3/M1/s1 ));
 AND2_X1 \V3/V4/V3/A3/M1/M2/_0_  (.A1(\V3/V4/V3/A3/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M1/M2/_1_  (.A(\V3/V4/V3/A3/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/v3 [4]));
 OR2_X1 \V3/V4/V3/A3/M1/_0_  (.A1(\V3/V4/V3/A3/M1/c1 ),
    .A2(\V3/V4/V3/A3/M1/c2 ),
    .ZN(\V3/V4/V3/A3/c1 ));
 AND2_X1 \V3/V4/V3/A3/M2/M1/_0_  (.A1(\V3/V4/V3/v4 [1]),
    .A2(\V3/V4/V3/s2 [3]),
    .ZN(\V3/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M2/M1/_1_  (.A(\V3/V4/V3/v4 [1]),
    .B(\V3/V4/V3/s2 [3]),
    .Z(\V3/V4/V3/A3/M2/s1 ));
 AND2_X1 \V3/V4/V3/A3/M2/M2/_0_  (.A1(\V3/V4/V3/A3/M2/s1 ),
    .A2(\V3/V4/V3/A3/c1 ),
    .ZN(\V3/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M2/M2/_1_  (.A(\V3/V4/V3/A3/M2/s1 ),
    .B(\V3/V4/V3/A3/c1 ),
    .Z(\V3/V4/v3 [5]));
 OR2_X1 \V3/V4/V3/A3/M2/_0_  (.A1(\V3/V4/V3/A3/M2/c1 ),
    .A2(\V3/V4/V3/A3/M2/c2 ),
    .ZN(\V3/V4/V3/A3/c2 ));
 AND2_X1 \V3/V4/V3/A3/M3/M1/_0_  (.A1(\V3/V4/V3/v4 [2]),
    .A2(\V3/V4/V3/c3 ),
    .ZN(\V3/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M3/M1/_1_  (.A(\V3/V4/V3/v4 [2]),
    .B(\V3/V4/V3/c3 ),
    .Z(\V3/V4/V3/A3/M3/s1 ));
 AND2_X1 \V3/V4/V3/A3/M3/M2/_0_  (.A1(\V3/V4/V3/A3/M3/s1 ),
    .A2(\V3/V4/V3/A3/c2 ),
    .ZN(\V3/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M3/M2/_1_  (.A(\V3/V4/V3/A3/M3/s1 ),
    .B(\V3/V4/V3/A3/c2 ),
    .Z(\V3/V4/v3 [6]));
 OR2_X1 \V3/V4/V3/A3/M3/_0_  (.A1(\V3/V4/V3/A3/M3/c1 ),
    .A2(\V3/V4/V3/A3/M3/c2 ),
    .ZN(\V3/V4/V3/A3/c3 ));
 AND2_X1 \V3/V4/V3/A3/M4/M1/_0_  (.A1(\V3/V4/V3/v4 [3]),
    .A2(net8),
    .ZN(\V3/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V3/A3/M4/M1/_1_  (.A(\V3/V4/V3/v4 [3]),
    .B(net8),
    .Z(\V3/V4/V3/A3/M4/s1 ));
 AND2_X1 \V3/V4/V3/A3/M4/M2/_0_  (.A1(\V3/V4/V3/A3/M4/s1 ),
    .A2(\V3/V4/V3/A3/c3 ),
    .ZN(\V3/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V3/A3/M4/M2/_1_  (.A(\V3/V4/V3/A3/M4/s1 ),
    .B(\V3/V4/V3/A3/c3 ),
    .Z(\V3/V4/v3 [7]));
 OR2_X1 \V3/V4/V3/A3/M4/_0_  (.A1(\V3/V4/V3/A3/M4/c1 ),
    .A2(\V3/V4/V3/A3/M4/c2 ),
    .ZN(\V3/V4/V3/overflow ));
 AND2_X1 \V3/V4/V3/V1/HA1/_0_  (.A1(\V3/V4/V3/V1/w2 ),
    .A2(\V3/V4/V3/V1/w1 ),
    .ZN(\V3/V4/V3/V1/w4 ));
 XOR2_X2 \V3/V4/V3/V1/HA1/_1_  (.A(\V3/V4/V3/V1/w2 ),
    .B(\V3/V4/V3/V1/w1 ),
    .Z(\V3/V4/v3 [1]));
 AND2_X1 \V3/V4/V3/V1/HA2/_0_  (.A1(\V3/V4/V3/V1/w4 ),
    .A2(\V3/V4/V3/V1/w3 ),
    .ZN(\V3/V4/V3/v1 [3]));
 XOR2_X2 \V3/V4/V3/V1/HA2/_1_  (.A(\V3/V4/V3/V1/w4 ),
    .B(\V3/V4/V3/V1/w3 ),
    .Z(\V3/V4/V3/v1 [2]));
 AND2_X1 \V3/V4/V3/V1/_0_  (.A1(net25),
    .A2(B[28]),
    .ZN(\V3/V4/v3 [0]));
 AND2_X1 \V3/V4/V3/V1/_1_  (.A1(net25),
    .A2(B[29]),
    .ZN(\V3/V4/V3/V1/w1 ));
 AND2_X1 \V3/V4/V3/V1/_2_  (.A1(B[28]),
    .A2(net24),
    .ZN(\V3/V4/V3/V1/w2 ));
 AND2_X1 \V3/V4/V3/V1/_3_  (.A1(B[29]),
    .A2(net24),
    .ZN(\V3/V4/V3/V1/w3 ));
 AND2_X1 \V3/V4/V3/V2/HA1/_0_  (.A1(\V3/V4/V3/V2/w2 ),
    .A2(\V3/V4/V3/V2/w1 ),
    .ZN(\V3/V4/V3/V2/w4 ));
 XOR2_X2 \V3/V4/V3/V2/HA1/_1_  (.A(\V3/V4/V3/V2/w2 ),
    .B(\V3/V4/V3/V2/w1 ),
    .Z(\V3/V4/V3/v2 [1]));
 AND2_X1 \V3/V4/V3/V2/HA2/_0_  (.A1(\V3/V4/V3/V2/w4 ),
    .A2(\V3/V4/V3/V2/w3 ),
    .ZN(\V3/V4/V3/v2 [3]));
 XOR2_X2 \V3/V4/V3/V2/HA2/_1_  (.A(\V3/V4/V3/V2/w4 ),
    .B(\V3/V4/V3/V2/w3 ),
    .Z(\V3/V4/V3/v2 [2]));
 AND2_X1 \V3/V4/V3/V2/_0_  (.A1(net47),
    .A2(B[28]),
    .ZN(\V3/V4/V3/v2 [0]));
 AND2_X1 \V3/V4/V3/V2/_1_  (.A1(net47),
    .A2(B[29]),
    .ZN(\V3/V4/V3/V2/w1 ));
 AND2_X1 \V3/V4/V3/V2/_2_  (.A1(B[28]),
    .A2(net46),
    .ZN(\V3/V4/V3/V2/w2 ));
 AND2_X1 \V3/V4/V3/V2/_3_  (.A1(B[29]),
    .A2(net46),
    .ZN(\V3/V4/V3/V2/w3 ));
 AND2_X1 \V3/V4/V3/V3/HA1/_0_  (.A1(\V3/V4/V3/V3/w2 ),
    .A2(\V3/V4/V3/V3/w1 ),
    .ZN(\V3/V4/V3/V3/w4 ));
 XOR2_X2 \V3/V4/V3/V3/HA1/_1_  (.A(\V3/V4/V3/V3/w2 ),
    .B(\V3/V4/V3/V3/w1 ),
    .Z(\V3/V4/V3/v3 [1]));
 AND2_X1 \V3/V4/V3/V3/HA2/_0_  (.A1(\V3/V4/V3/V3/w4 ),
    .A2(\V3/V4/V3/V3/w3 ),
    .ZN(\V3/V4/V3/v3 [3]));
 XOR2_X2 \V3/V4/V3/V3/HA2/_1_  (.A(\V3/V4/V3/V3/w4 ),
    .B(\V3/V4/V3/V3/w3 ),
    .Z(\V3/V4/V3/v3 [2]));
 AND2_X1 \V3/V4/V3/V3/_0_  (.A1(net25),
    .A2(B[30]),
    .ZN(\V3/V4/V3/v3 [0]));
 AND2_X1 \V3/V4/V3/V3/_1_  (.A1(net25),
    .A2(B[31]),
    .ZN(\V3/V4/V3/V3/w1 ));
 AND2_X1 \V3/V4/V3/V3/_2_  (.A1(B[30]),
    .A2(net24),
    .ZN(\V3/V4/V3/V3/w2 ));
 AND2_X1 \V3/V4/V3/V3/_3_  (.A1(B[31]),
    .A2(net24),
    .ZN(\V3/V4/V3/V3/w3 ));
 AND2_X1 \V3/V4/V3/V4/HA1/_0_  (.A1(\V3/V4/V3/V4/w2 ),
    .A2(\V3/V4/V3/V4/w1 ),
    .ZN(\V3/V4/V3/V4/w4 ));
 XOR2_X2 \V3/V4/V3/V4/HA1/_1_  (.A(\V3/V4/V3/V4/w2 ),
    .B(\V3/V4/V3/V4/w1 ),
    .Z(\V3/V4/V3/v4 [1]));
 AND2_X1 \V3/V4/V3/V4/HA2/_0_  (.A1(\V3/V4/V3/V4/w4 ),
    .A2(\V3/V4/V3/V4/w3 ),
    .ZN(\V3/V4/V3/v4 [3]));
 XOR2_X2 \V3/V4/V3/V4/HA2/_1_  (.A(\V3/V4/V3/V4/w4 ),
    .B(\V3/V4/V3/V4/w3 ),
    .Z(\V3/V4/V3/v4 [2]));
 AND2_X1 \V3/V4/V3/V4/_0_  (.A1(net47),
    .A2(B[30]),
    .ZN(\V3/V4/V3/v4 [0]));
 AND2_X1 \V3/V4/V3/V4/_1_  (.A1(net47),
    .A2(B[31]),
    .ZN(\V3/V4/V3/V4/w1 ));
 AND2_X1 \V3/V4/V3/V4/_2_  (.A1(B[30]),
    .A2(net46),
    .ZN(\V3/V4/V3/V4/w2 ));
 AND2_X1 \V3/V4/V3/V4/_3_  (.A1(B[31]),
    .A2(net46),
    .ZN(\V3/V4/V3/V4/w3 ));
 OR2_X1 \V3/V4/V3/_0_  (.A1(\V3/V4/V3/c1 ),
    .A2(\V3/V4/V3/c2 ),
    .ZN(\V3/V4/V3/c3 ));
 AND2_X1 \V3/V4/V4/A1/M1/M1/_0_  (.A1(\V3/V4/V4/v2 [0]),
    .A2(\V3/V4/V4/v3 [0]),
    .ZN(\V3/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M1/M1/_1_  (.A(\V3/V4/V4/v2 [0]),
    .B(\V3/V4/V4/v3 [0]),
    .Z(\V3/V4/V4/A1/M1/s1 ));
 AND2_X1 \V3/V4/V4/A1/M1/M2/_0_  (.A1(\V3/V4/V4/A1/M1/s1 ),
    .A2(net8),
    .ZN(\V3/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M1/M2/_1_  (.A(\V3/V4/V4/A1/M1/s1 ),
    .B(net8),
    .Z(\V3/V4/V4/s1 [0]));
 OR2_X1 \V3/V4/V4/A1/M1/_0_  (.A1(\V3/V4/V4/A1/M1/c1 ),
    .A2(\V3/V4/V4/A1/M1/c2 ),
    .ZN(\V3/V4/V4/A1/c1 ));
 AND2_X1 \V3/V4/V4/A1/M2/M1/_0_  (.A1(\V3/V4/V4/v2 [1]),
    .A2(\V3/V4/V4/v3 [1]),
    .ZN(\V3/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M2/M1/_1_  (.A(\V3/V4/V4/v2 [1]),
    .B(\V3/V4/V4/v3 [1]),
    .Z(\V3/V4/V4/A1/M2/s1 ));
 AND2_X1 \V3/V4/V4/A1/M2/M2/_0_  (.A1(\V3/V4/V4/A1/M2/s1 ),
    .A2(\V3/V4/V4/A1/c1 ),
    .ZN(\V3/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M2/M2/_1_  (.A(\V3/V4/V4/A1/M2/s1 ),
    .B(\V3/V4/V4/A1/c1 ),
    .Z(\V3/V4/V4/s1 [1]));
 OR2_X1 \V3/V4/V4/A1/M2/_0_  (.A1(\V3/V4/V4/A1/M2/c1 ),
    .A2(\V3/V4/V4/A1/M2/c2 ),
    .ZN(\V3/V4/V4/A1/c2 ));
 AND2_X1 \V3/V4/V4/A1/M3/M1/_0_  (.A1(\V3/V4/V4/v2 [2]),
    .A2(\V3/V4/V4/v3 [2]),
    .ZN(\V3/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M3/M1/_1_  (.A(\V3/V4/V4/v2 [2]),
    .B(\V3/V4/V4/v3 [2]),
    .Z(\V3/V4/V4/A1/M3/s1 ));
 AND2_X1 \V3/V4/V4/A1/M3/M2/_0_  (.A1(\V3/V4/V4/A1/M3/s1 ),
    .A2(\V3/V4/V4/A1/c2 ),
    .ZN(\V3/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M3/M2/_1_  (.A(\V3/V4/V4/A1/M3/s1 ),
    .B(\V3/V4/V4/A1/c2 ),
    .Z(\V3/V4/V4/s1 [2]));
 OR2_X1 \V3/V4/V4/A1/M3/_0_  (.A1(\V3/V4/V4/A1/M3/c1 ),
    .A2(\V3/V4/V4/A1/M3/c2 ),
    .ZN(\V3/V4/V4/A1/c3 ));
 AND2_X1 \V3/V4/V4/A1/M4/M1/_0_  (.A1(\V3/V4/V4/v2 [3]),
    .A2(\V3/V4/V4/v3 [3]),
    .ZN(\V3/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A1/M4/M1/_1_  (.A(\V3/V4/V4/v2 [3]),
    .B(\V3/V4/V4/v3 [3]),
    .Z(\V3/V4/V4/A1/M4/s1 ));
 AND2_X1 \V3/V4/V4/A1/M4/M2/_0_  (.A1(\V3/V4/V4/A1/M4/s1 ),
    .A2(\V3/V4/V4/A1/c3 ),
    .ZN(\V3/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A1/M4/M2/_1_  (.A(\V3/V4/V4/A1/M4/s1 ),
    .B(\V3/V4/V4/A1/c3 ),
    .Z(\V3/V4/V4/s1 [3]));
 OR2_X1 \V3/V4/V4/A1/M4/_0_  (.A1(\V3/V4/V4/A1/M4/c1 ),
    .A2(\V3/V4/V4/A1/M4/c2 ),
    .ZN(\V3/V4/V4/c1 ));
 AND2_X1 \V3/V4/V4/A2/M1/M1/_0_  (.A1(\V3/V4/V4/s1 [0]),
    .A2(\V3/V4/V4/v1 [2]),
    .ZN(\V3/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M1/M1/_1_  (.A(\V3/V4/V4/s1 [0]),
    .B(\V3/V4/V4/v1 [2]),
    .Z(\V3/V4/V4/A2/M1/s1 ));
 AND2_X1 \V3/V4/V4/A2/M1/M2/_0_  (.A1(\V3/V4/V4/A2/M1/s1 ),
    .A2(net7),
    .ZN(\V3/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M1/M2/_1_  (.A(\V3/V4/V4/A2/M1/s1 ),
    .B(net7),
    .Z(\V3/V4/v4 [2]));
 OR2_X1 \V3/V4/V4/A2/M1/_0_  (.A1(\V3/V4/V4/A2/M1/c1 ),
    .A2(\V3/V4/V4/A2/M1/c2 ),
    .ZN(\V3/V4/V4/A2/c1 ));
 AND2_X1 \V3/V4/V4/A2/M2/M1/_0_  (.A1(\V3/V4/V4/s1 [1]),
    .A2(\V3/V4/V4/v1 [3]),
    .ZN(\V3/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M2/M1/_1_  (.A(\V3/V4/V4/s1 [1]),
    .B(\V3/V4/V4/v1 [3]),
    .Z(\V3/V4/V4/A2/M2/s1 ));
 AND2_X1 \V3/V4/V4/A2/M2/M2/_0_  (.A1(\V3/V4/V4/A2/M2/s1 ),
    .A2(\V3/V4/V4/A2/c1 ),
    .ZN(\V3/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M2/M2/_1_  (.A(\V3/V4/V4/A2/M2/s1 ),
    .B(\V3/V4/V4/A2/c1 ),
    .Z(\V3/V4/v4 [3]));
 OR2_X1 \V3/V4/V4/A2/M2/_0_  (.A1(\V3/V4/V4/A2/M2/c1 ),
    .A2(\V3/V4/V4/A2/M2/c2 ),
    .ZN(\V3/V4/V4/A2/c2 ));
 AND2_X1 \V3/V4/V4/A2/M3/M1/_0_  (.A1(\V3/V4/V4/s1 [2]),
    .A2(net8),
    .ZN(\V3/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M3/M1/_1_  (.A(\V3/V4/V4/s1 [2]),
    .B(net8),
    .Z(\V3/V4/V4/A2/M3/s1 ));
 AND2_X1 \V3/V4/V4/A2/M3/M2/_0_  (.A1(\V3/V4/V4/A2/M3/s1 ),
    .A2(\V3/V4/V4/A2/c2 ),
    .ZN(\V3/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M3/M2/_1_  (.A(\V3/V4/V4/A2/M3/s1 ),
    .B(\V3/V4/V4/A2/c2 ),
    .Z(\V3/V4/V4/s2 [2]));
 OR2_X1 \V3/V4/V4/A2/M3/_0_  (.A1(\V3/V4/V4/A2/M3/c1 ),
    .A2(\V3/V4/V4/A2/M3/c2 ),
    .ZN(\V3/V4/V4/A2/c3 ));
 AND2_X1 \V3/V4/V4/A2/M4/M1/_0_  (.A1(\V3/V4/V4/s1 [3]),
    .A2(net8),
    .ZN(\V3/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A2/M4/M1/_1_  (.A(\V3/V4/V4/s1 [3]),
    .B(net8),
    .Z(\V3/V4/V4/A2/M4/s1 ));
 AND2_X1 \V3/V4/V4/A2/M4/M2/_0_  (.A1(\V3/V4/V4/A2/M4/s1 ),
    .A2(\V3/V4/V4/A2/c3 ),
    .ZN(\V3/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A2/M4/M2/_1_  (.A(\V3/V4/V4/A2/M4/s1 ),
    .B(\V3/V4/V4/A2/c3 ),
    .Z(\V3/V4/V4/s2 [3]));
 OR2_X1 \V3/V4/V4/A2/M4/_0_  (.A1(\V3/V4/V4/A2/M4/c1 ),
    .A2(\V3/V4/V4/A2/M4/c2 ),
    .ZN(\V3/V4/V4/c2 ));
 AND2_X1 \V3/V4/V4/A3/M1/M1/_0_  (.A1(\V3/V4/V4/v4 [0]),
    .A2(\V3/V4/V4/s2 [2]),
    .ZN(\V3/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M1/M1/_1_  (.A(\V3/V4/V4/v4 [0]),
    .B(\V3/V4/V4/s2 [2]),
    .Z(\V3/V4/V4/A3/M1/s1 ));
 AND2_X1 \V3/V4/V4/A3/M1/M2/_0_  (.A1(\V3/V4/V4/A3/M1/s1 ),
    .A2(net7),
    .ZN(\V3/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M1/M2/_1_  (.A(\V3/V4/V4/A3/M1/s1 ),
    .B(net7),
    .Z(\V3/V4/v4 [4]));
 OR2_X1 \V3/V4/V4/A3/M1/_0_  (.A1(\V3/V4/V4/A3/M1/c1 ),
    .A2(\V3/V4/V4/A3/M1/c2 ),
    .ZN(\V3/V4/V4/A3/c1 ));
 AND2_X1 \V3/V4/V4/A3/M2/M1/_0_  (.A1(\V3/V4/V4/v4 [1]),
    .A2(\V3/V4/V4/s2 [3]),
    .ZN(\V3/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M2/M1/_1_  (.A(\V3/V4/V4/v4 [1]),
    .B(\V3/V4/V4/s2 [3]),
    .Z(\V3/V4/V4/A3/M2/s1 ));
 AND2_X1 \V3/V4/V4/A3/M2/M2/_0_  (.A1(\V3/V4/V4/A3/M2/s1 ),
    .A2(\V3/V4/V4/A3/c1 ),
    .ZN(\V3/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M2/M2/_1_  (.A(\V3/V4/V4/A3/M2/s1 ),
    .B(\V3/V4/V4/A3/c1 ),
    .Z(\V3/V4/v4 [5]));
 OR2_X1 \V3/V4/V4/A3/M2/_0_  (.A1(\V3/V4/V4/A3/M2/c1 ),
    .A2(\V3/V4/V4/A3/M2/c2 ),
    .ZN(\V3/V4/V4/A3/c2 ));
 AND2_X1 \V3/V4/V4/A3/M3/M1/_0_  (.A1(\V3/V4/V4/v4 [2]),
    .A2(\V3/V4/V4/c3 ),
    .ZN(\V3/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M3/M1/_1_  (.A(\V3/V4/V4/v4 [2]),
    .B(\V3/V4/V4/c3 ),
    .Z(\V3/V4/V4/A3/M3/s1 ));
 AND2_X1 \V3/V4/V4/A3/M3/M2/_0_  (.A1(\V3/V4/V4/A3/M3/s1 ),
    .A2(\V3/V4/V4/A3/c2 ),
    .ZN(\V3/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M3/M2/_1_  (.A(\V3/V4/V4/A3/M3/s1 ),
    .B(\V3/V4/V4/A3/c2 ),
    .Z(\V3/V4/v4 [6]));
 OR2_X1 \V3/V4/V4/A3/M3/_0_  (.A1(\V3/V4/V4/A3/M3/c1 ),
    .A2(\V3/V4/V4/A3/M3/c2 ),
    .ZN(\V3/V4/V4/A3/c3 ));
 AND2_X1 \V3/V4/V4/A3/M4/M1/_0_  (.A1(\V3/V4/V4/v4 [3]),
    .A2(net8),
    .ZN(\V3/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V3/V4/V4/A3/M4/M1/_1_  (.A(\V3/V4/V4/v4 [3]),
    .B(net8),
    .Z(\V3/V4/V4/A3/M4/s1 ));
 AND2_X1 \V3/V4/V4/A3/M4/M2/_0_  (.A1(\V3/V4/V4/A3/M4/s1 ),
    .A2(\V3/V4/V4/A3/c3 ),
    .ZN(\V3/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V3/V4/V4/A3/M4/M2/_1_  (.A(\V3/V4/V4/A3/M4/s1 ),
    .B(\V3/V4/V4/A3/c3 ),
    .Z(\V3/V4/v4 [7]));
 OR2_X1 \V3/V4/V4/A3/M4/_0_  (.A1(\V3/V4/V4/A3/M4/c1 ),
    .A2(\V3/V4/V4/A3/M4/c2 ),
    .ZN(\V3/V4/V4/overflow ));
 AND2_X1 \V3/V4/V4/V1/HA1/_0_  (.A1(\V3/V4/V4/V1/w2 ),
    .A2(\V3/V4/V4/V1/w1 ),
    .ZN(\V3/V4/V4/V1/w4 ));
 XOR2_X2 \V3/V4/V4/V1/HA1/_1_  (.A(\V3/V4/V4/V1/w2 ),
    .B(\V3/V4/V4/V1/w1 ),
    .Z(\V3/V4/v4 [1]));
 AND2_X1 \V3/V4/V4/V1/HA2/_0_  (.A1(\V3/V4/V4/V1/w4 ),
    .A2(\V3/V4/V4/V1/w3 ),
    .ZN(\V3/V4/V4/v1 [3]));
 XOR2_X2 \V3/V4/V4/V1/HA2/_1_  (.A(\V3/V4/V4/V1/w4 ),
    .B(\V3/V4/V4/V1/w3 ),
    .Z(\V3/V4/V4/v1 [2]));
 AND2_X1 \V3/V4/V4/V1/_0_  (.A1(net45),
    .A2(B[28]),
    .ZN(\V3/V4/v4 [0]));
 AND2_X1 \V3/V4/V4/V1/_1_  (.A1(net45),
    .A2(B[29]),
    .ZN(\V3/V4/V4/V1/w1 ));
 AND2_X1 \V3/V4/V4/V1/_2_  (.A1(B[28]),
    .A2(net44),
    .ZN(\V3/V4/V4/V1/w2 ));
 AND2_X1 \V3/V4/V4/V1/_3_  (.A1(B[29]),
    .A2(net44),
    .ZN(\V3/V4/V4/V1/w3 ));
 AND2_X1 \V3/V4/V4/V2/HA1/_0_  (.A1(\V3/V4/V4/V2/w2 ),
    .A2(\V3/V4/V4/V2/w1 ),
    .ZN(\V3/V4/V4/V2/w4 ));
 XOR2_X2 \V3/V4/V4/V2/HA1/_1_  (.A(\V3/V4/V4/V2/w2 ),
    .B(\V3/V4/V4/V2/w1 ),
    .Z(\V3/V4/V4/v2 [1]));
 AND2_X1 \V3/V4/V4/V2/HA2/_0_  (.A1(\V3/V4/V4/V2/w4 ),
    .A2(\V3/V4/V4/V2/w3 ),
    .ZN(\V3/V4/V4/v2 [3]));
 XOR2_X2 \V3/V4/V4/V2/HA2/_1_  (.A(\V3/V4/V4/V2/w4 ),
    .B(\V3/V4/V4/V2/w3 ),
    .Z(\V3/V4/V4/v2 [2]));
 AND2_X1 \V3/V4/V4/V2/_0_  (.A1(net43),
    .A2(B[28]),
    .ZN(\V3/V4/V4/v2 [0]));
 AND2_X1 \V3/V4/V4/V2/_1_  (.A1(net43),
    .A2(B[29]),
    .ZN(\V3/V4/V4/V2/w1 ));
 AND2_X1 \V3/V4/V4/V2/_2_  (.A1(B[28]),
    .A2(net42),
    .ZN(\V3/V4/V4/V2/w2 ));
 AND2_X1 \V3/V4/V4/V2/_3_  (.A1(B[29]),
    .A2(net42),
    .ZN(\V3/V4/V4/V2/w3 ));
 AND2_X1 \V3/V4/V4/V3/HA1/_0_  (.A1(\V3/V4/V4/V3/w2 ),
    .A2(\V3/V4/V4/V3/w1 ),
    .ZN(\V3/V4/V4/V3/w4 ));
 XOR2_X2 \V3/V4/V4/V3/HA1/_1_  (.A(\V3/V4/V4/V3/w2 ),
    .B(\V3/V4/V4/V3/w1 ),
    .Z(\V3/V4/V4/v3 [1]));
 AND2_X1 \V3/V4/V4/V3/HA2/_0_  (.A1(\V3/V4/V4/V3/w4 ),
    .A2(\V3/V4/V4/V3/w3 ),
    .ZN(\V3/V4/V4/v3 [3]));
 XOR2_X2 \V3/V4/V4/V3/HA2/_1_  (.A(\V3/V4/V4/V3/w4 ),
    .B(\V3/V4/V4/V3/w3 ),
    .Z(\V3/V4/V4/v3 [2]));
 AND2_X1 \V3/V4/V4/V3/_0_  (.A1(net45),
    .A2(B[30]),
    .ZN(\V3/V4/V4/v3 [0]));
 AND2_X1 \V3/V4/V4/V3/_1_  (.A1(net45),
    .A2(B[31]),
    .ZN(\V3/V4/V4/V3/w1 ));
 AND2_X1 \V3/V4/V4/V3/_2_  (.A1(B[30]),
    .A2(net44),
    .ZN(\V3/V4/V4/V3/w2 ));
 AND2_X1 \V3/V4/V4/V3/_3_  (.A1(B[31]),
    .A2(net44),
    .ZN(\V3/V4/V4/V3/w3 ));
 AND2_X1 \V3/V4/V4/V4/HA1/_0_  (.A1(\V3/V4/V4/V4/w2 ),
    .A2(\V3/V4/V4/V4/w1 ),
    .ZN(\V3/V4/V4/V4/w4 ));
 XOR2_X2 \V3/V4/V4/V4/HA1/_1_  (.A(\V3/V4/V4/V4/w2 ),
    .B(\V3/V4/V4/V4/w1 ),
    .Z(\V3/V4/V4/v4 [1]));
 AND2_X1 \V3/V4/V4/V4/HA2/_0_  (.A1(\V3/V4/V4/V4/w4 ),
    .A2(\V3/V4/V4/V4/w3 ),
    .ZN(\V3/V4/V4/v4 [3]));
 XOR2_X2 \V3/V4/V4/V4/HA2/_1_  (.A(\V3/V4/V4/V4/w4 ),
    .B(\V3/V4/V4/V4/w3 ),
    .Z(\V3/V4/V4/v4 [2]));
 AND2_X1 \V3/V4/V4/V4/_0_  (.A1(net43),
    .A2(B[30]),
    .ZN(\V3/V4/V4/v4 [0]));
 AND2_X1 \V3/V4/V4/V4/_1_  (.A1(net43),
    .A2(B[31]),
    .ZN(\V3/V4/V4/V4/w1 ));
 AND2_X1 \V3/V4/V4/V4/_2_  (.A1(B[30]),
    .A2(net42),
    .ZN(\V3/V4/V4/V4/w2 ));
 AND2_X1 \V3/V4/V4/V4/_3_  (.A1(B[31]),
    .A2(net42),
    .ZN(\V3/V4/V4/V4/w3 ));
 OR2_X1 \V3/V4/V4/_0_  (.A1(\V3/V4/V4/c1 ),
    .A2(\V3/V4/V4/c2 ),
    .ZN(\V3/V4/V4/c3 ));
 OR2_X1 \V3/V4/_0_  (.A1(\V3/V4/c1 ),
    .A2(\V3/V4/c2 ),
    .ZN(\V3/V4/c3 ));
 OR2_X1 \V3/_0_  (.A1(\V3/c1 ),
    .A2(\V3/c2 ),
    .ZN(\V3/c3 ));
 AND2_X1 \V4/A1/A1/A1/M1/M1/_0_  (.A1(\V4/v2 [0]),
    .A2(\V4/v3 [0]),
    .ZN(\V4/A1/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M1/M1/_1_  (.A(\V4/v2 [0]),
    .B(\V4/v3 [0]),
    .Z(\V4/A1/A1/A1/M1/s1 ));
 AND2_X1 \V4/A1/A1/A1/M1/M2/_0_  (.A1(\V4/A1/A1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/A1/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M1/M2/_1_  (.A(\V4/A1/A1/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/s1 [0]));
 OR2_X1 \V4/A1/A1/A1/M1/_0_  (.A1(\V4/A1/A1/A1/M1/c1 ),
    .A2(\V4/A1/A1/A1/M1/c2 ),
    .ZN(\V4/A1/A1/A1/c1 ));
 AND2_X1 \V4/A1/A1/A1/M2/M1/_0_  (.A1(\V4/v2 [1]),
    .A2(\V4/v3 [1]),
    .ZN(\V4/A1/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M2/M1/_1_  (.A(\V4/v2 [1]),
    .B(\V4/v3 [1]),
    .Z(\V4/A1/A1/A1/M2/s1 ));
 AND2_X1 \V4/A1/A1/A1/M2/M2/_0_  (.A1(\V4/A1/A1/A1/M2/s1 ),
    .A2(\V4/A1/A1/A1/c1 ),
    .ZN(\V4/A1/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M2/M2/_1_  (.A(\V4/A1/A1/A1/M2/s1 ),
    .B(\V4/A1/A1/A1/c1 ),
    .Z(\V4/s1 [1]));
 OR2_X1 \V4/A1/A1/A1/M2/_0_  (.A1(\V4/A1/A1/A1/M2/c1 ),
    .A2(\V4/A1/A1/A1/M2/c2 ),
    .ZN(\V4/A1/A1/A1/c2 ));
 AND2_X1 \V4/A1/A1/A1/M3/M1/_0_  (.A1(\V4/v2 [2]),
    .A2(\V4/v3 [2]),
    .ZN(\V4/A1/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M3/M1/_1_  (.A(\V4/v2 [2]),
    .B(\V4/v3 [2]),
    .Z(\V4/A1/A1/A1/M3/s1 ));
 AND2_X1 \V4/A1/A1/A1/M3/M2/_0_  (.A1(\V4/A1/A1/A1/M3/s1 ),
    .A2(\V4/A1/A1/A1/c2 ),
    .ZN(\V4/A1/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M3/M2/_1_  (.A(\V4/A1/A1/A1/M3/s1 ),
    .B(\V4/A1/A1/A1/c2 ),
    .Z(\V4/s1 [2]));
 OR2_X1 \V4/A1/A1/A1/M3/_0_  (.A1(\V4/A1/A1/A1/M3/c1 ),
    .A2(\V4/A1/A1/A1/M3/c2 ),
    .ZN(\V4/A1/A1/A1/c3 ));
 AND2_X1 \V4/A1/A1/A1/M4/M1/_0_  (.A1(\V4/v2 [3]),
    .A2(\V4/v3 [3]),
    .ZN(\V4/A1/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A1/A1/A1/M4/M1/_1_  (.A(\V4/v2 [3]),
    .B(\V4/v3 [3]),
    .Z(\V4/A1/A1/A1/M4/s1 ));
 AND2_X1 \V4/A1/A1/A1/M4/M2/_0_  (.A1(\V4/A1/A1/A1/M4/s1 ),
    .A2(\V4/A1/A1/A1/c3 ),
    .ZN(\V4/A1/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A1/A1/A1/M4/M2/_1_  (.A(\V4/A1/A1/A1/M4/s1 ),
    .B(\V4/A1/A1/A1/c3 ),
    .Z(\V4/s1 [3]));
 OR2_X1 \V4/A1/A1/A1/M4/_0_  (.A1(\V4/A1/A1/A1/M4/c1 ),
    .A2(\V4/A1/A1/A1/M4/c2 ),
    .ZN(\V4/A1/A1/c1 ));
 AND2_X1 \V4/A1/A1/A2/M1/M1/_0_  (.A1(\V4/v2 [4]),
    .A2(\V4/v3 [4]),
    .ZN(\V4/A1/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M1/M1/_1_  (.A(\V4/v2 [4]),
    .B(\V4/v3 [4]),
    .Z(\V4/A1/A1/A2/M1/s1 ));
 AND2_X1 \V4/A1/A1/A2/M1/M2/_0_  (.A1(\V4/A1/A1/A2/M1/s1 ),
    .A2(\V4/A1/A1/c1 ),
    .ZN(\V4/A1/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M1/M2/_1_  (.A(\V4/A1/A1/A2/M1/s1 ),
    .B(\V4/A1/A1/c1 ),
    .Z(\V4/s1 [4]));
 OR2_X1 \V4/A1/A1/A2/M1/_0_  (.A1(\V4/A1/A1/A2/M1/c1 ),
    .A2(\V4/A1/A1/A2/M1/c2 ),
    .ZN(\V4/A1/A1/A2/c1 ));
 AND2_X1 \V4/A1/A1/A2/M2/M1/_0_  (.A1(\V4/v2 [5]),
    .A2(\V4/v3 [5]),
    .ZN(\V4/A1/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M2/M1/_1_  (.A(\V4/v2 [5]),
    .B(\V4/v3 [5]),
    .Z(\V4/A1/A1/A2/M2/s1 ));
 AND2_X1 \V4/A1/A1/A2/M2/M2/_0_  (.A1(\V4/A1/A1/A2/M2/s1 ),
    .A2(\V4/A1/A1/A2/c1 ),
    .ZN(\V4/A1/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M2/M2/_1_  (.A(\V4/A1/A1/A2/M2/s1 ),
    .B(\V4/A1/A1/A2/c1 ),
    .Z(\V4/s1 [5]));
 OR2_X1 \V4/A1/A1/A2/M2/_0_  (.A1(\V4/A1/A1/A2/M2/c1 ),
    .A2(\V4/A1/A1/A2/M2/c2 ),
    .ZN(\V4/A1/A1/A2/c2 ));
 AND2_X1 \V4/A1/A1/A2/M3/M1/_0_  (.A1(\V4/v2 [6]),
    .A2(\V4/v3 [6]),
    .ZN(\V4/A1/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M3/M1/_1_  (.A(\V4/v2 [6]),
    .B(\V4/v3 [6]),
    .Z(\V4/A1/A1/A2/M3/s1 ));
 AND2_X1 \V4/A1/A1/A2/M3/M2/_0_  (.A1(\V4/A1/A1/A2/M3/s1 ),
    .A2(\V4/A1/A1/A2/c2 ),
    .ZN(\V4/A1/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M3/M2/_1_  (.A(\V4/A1/A1/A2/M3/s1 ),
    .B(\V4/A1/A1/A2/c2 ),
    .Z(\V4/s1 [6]));
 OR2_X1 \V4/A1/A1/A2/M3/_0_  (.A1(\V4/A1/A1/A2/M3/c1 ),
    .A2(\V4/A1/A1/A2/M3/c2 ),
    .ZN(\V4/A1/A1/A2/c3 ));
 AND2_X1 \V4/A1/A1/A2/M4/M1/_0_  (.A1(\V4/v2 [7]),
    .A2(\V4/v3 [7]),
    .ZN(\V4/A1/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A1/A1/A2/M4/M1/_1_  (.A(\V4/v2 [7]),
    .B(\V4/v3 [7]),
    .Z(\V4/A1/A1/A2/M4/s1 ));
 AND2_X1 \V4/A1/A1/A2/M4/M2/_0_  (.A1(\V4/A1/A1/A2/M4/s1 ),
    .A2(\V4/A1/A1/A2/c3 ),
    .ZN(\V4/A1/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A1/A1/A2/M4/M2/_1_  (.A(\V4/A1/A1/A2/M4/s1 ),
    .B(\V4/A1/A1/A2/c3 ),
    .Z(\V4/s1 [7]));
 OR2_X1 \V4/A1/A1/A2/M4/_0_  (.A1(\V4/A1/A1/A2/M4/c1 ),
    .A2(\V4/A1/A1/A2/M4/c2 ),
    .ZN(\V4/A1/c1 ));
 AND2_X1 \V4/A1/A2/A1/M1/M1/_0_  (.A1(\V4/v2 [8]),
    .A2(\V4/v3 [8]),
    .ZN(\V4/A1/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M1/M1/_1_  (.A(\V4/v2 [8]),
    .B(\V4/v3 [8]),
    .Z(\V4/A1/A2/A1/M1/s1 ));
 AND2_X1 \V4/A1/A2/A1/M1/M2/_0_  (.A1(\V4/A1/A2/A1/M1/s1 ),
    .A2(\V4/A1/c1 ),
    .ZN(\V4/A1/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M1/M2/_1_  (.A(\V4/A1/A2/A1/M1/s1 ),
    .B(\V4/A1/c1 ),
    .Z(\V4/s1 [8]));
 OR2_X1 \V4/A1/A2/A1/M1/_0_  (.A1(\V4/A1/A2/A1/M1/c1 ),
    .A2(\V4/A1/A2/A1/M1/c2 ),
    .ZN(\V4/A1/A2/A1/c1 ));
 AND2_X1 \V4/A1/A2/A1/M2/M1/_0_  (.A1(\V4/v2 [9]),
    .A2(\V4/v3 [9]),
    .ZN(\V4/A1/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M2/M1/_1_  (.A(\V4/v2 [9]),
    .B(\V4/v3 [9]),
    .Z(\V4/A1/A2/A1/M2/s1 ));
 AND2_X1 \V4/A1/A2/A1/M2/M2/_0_  (.A1(\V4/A1/A2/A1/M2/s1 ),
    .A2(\V4/A1/A2/A1/c1 ),
    .ZN(\V4/A1/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M2/M2/_1_  (.A(\V4/A1/A2/A1/M2/s1 ),
    .B(\V4/A1/A2/A1/c1 ),
    .Z(\V4/s1 [9]));
 OR2_X1 \V4/A1/A2/A1/M2/_0_  (.A1(\V4/A1/A2/A1/M2/c1 ),
    .A2(\V4/A1/A2/A1/M2/c2 ),
    .ZN(\V4/A1/A2/A1/c2 ));
 AND2_X1 \V4/A1/A2/A1/M3/M1/_0_  (.A1(\V4/v2 [10]),
    .A2(\V4/v3 [10]),
    .ZN(\V4/A1/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M3/M1/_1_  (.A(\V4/v2 [10]),
    .B(\V4/v3 [10]),
    .Z(\V4/A1/A2/A1/M3/s1 ));
 AND2_X1 \V4/A1/A2/A1/M3/M2/_0_  (.A1(\V4/A1/A2/A1/M3/s1 ),
    .A2(\V4/A1/A2/A1/c2 ),
    .ZN(\V4/A1/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M3/M2/_1_  (.A(\V4/A1/A2/A1/M3/s1 ),
    .B(\V4/A1/A2/A1/c2 ),
    .Z(\V4/s1 [10]));
 OR2_X1 \V4/A1/A2/A1/M3/_0_  (.A1(\V4/A1/A2/A1/M3/c1 ),
    .A2(\V4/A1/A2/A1/M3/c2 ),
    .ZN(\V4/A1/A2/A1/c3 ));
 AND2_X1 \V4/A1/A2/A1/M4/M1/_0_  (.A1(\V4/v2 [11]),
    .A2(\V4/v3 [11]),
    .ZN(\V4/A1/A2/A1/M4/c1 ));
 XOR2_X2 \V4/A1/A2/A1/M4/M1/_1_  (.A(\V4/v2 [11]),
    .B(\V4/v3 [11]),
    .Z(\V4/A1/A2/A1/M4/s1 ));
 AND2_X1 \V4/A1/A2/A1/M4/M2/_0_  (.A1(\V4/A1/A2/A1/M4/s1 ),
    .A2(\V4/A1/A2/A1/c3 ),
    .ZN(\V4/A1/A2/A1/M4/c2 ));
 XOR2_X2 \V4/A1/A2/A1/M4/M2/_1_  (.A(\V4/A1/A2/A1/M4/s1 ),
    .B(\V4/A1/A2/A1/c3 ),
    .Z(\V4/s1 [11]));
 OR2_X1 \V4/A1/A2/A1/M4/_0_  (.A1(\V4/A1/A2/A1/M4/c1 ),
    .A2(\V4/A1/A2/A1/M4/c2 ),
    .ZN(\V4/A1/A2/c1 ));
 AND2_X1 \V4/A1/A2/A2/M1/M1/_0_  (.A1(\V4/v2 [12]),
    .A2(\V4/v3 [12]),
    .ZN(\V4/A1/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M1/M1/_1_  (.A(\V4/v2 [12]),
    .B(\V4/v3 [12]),
    .Z(\V4/A1/A2/A2/M1/s1 ));
 AND2_X1 \V4/A1/A2/A2/M1/M2/_0_  (.A1(\V4/A1/A2/A2/M1/s1 ),
    .A2(\V4/A1/A2/c1 ),
    .ZN(\V4/A1/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M1/M2/_1_  (.A(\V4/A1/A2/A2/M1/s1 ),
    .B(\V4/A1/A2/c1 ),
    .Z(\V4/s1 [12]));
 OR2_X1 \V4/A1/A2/A2/M1/_0_  (.A1(\V4/A1/A2/A2/M1/c1 ),
    .A2(\V4/A1/A2/A2/M1/c2 ),
    .ZN(\V4/A1/A2/A2/c1 ));
 AND2_X1 \V4/A1/A2/A2/M2/M1/_0_  (.A1(\V4/v2 [13]),
    .A2(\V4/v3 [13]),
    .ZN(\V4/A1/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M2/M1/_1_  (.A(\V4/v2 [13]),
    .B(\V4/v3 [13]),
    .Z(\V4/A1/A2/A2/M2/s1 ));
 AND2_X1 \V4/A1/A2/A2/M2/M2/_0_  (.A1(\V4/A1/A2/A2/M2/s1 ),
    .A2(\V4/A1/A2/A2/c1 ),
    .ZN(\V4/A1/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M2/M2/_1_  (.A(\V4/A1/A2/A2/M2/s1 ),
    .B(\V4/A1/A2/A2/c1 ),
    .Z(\V4/s1 [13]));
 OR2_X1 \V4/A1/A2/A2/M2/_0_  (.A1(\V4/A1/A2/A2/M2/c1 ),
    .A2(\V4/A1/A2/A2/M2/c2 ),
    .ZN(\V4/A1/A2/A2/c2 ));
 AND2_X1 \V4/A1/A2/A2/M3/M1/_0_  (.A1(\V4/v2 [14]),
    .A2(\V4/v3 [14]),
    .ZN(\V4/A1/A2/A2/M3/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M3/M1/_1_  (.A(\V4/v2 [14]),
    .B(\V4/v3 [14]),
    .Z(\V4/A1/A2/A2/M3/s1 ));
 AND2_X1 \V4/A1/A2/A2/M3/M2/_0_  (.A1(\V4/A1/A2/A2/M3/s1 ),
    .A2(\V4/A1/A2/A2/c2 ),
    .ZN(\V4/A1/A2/A2/M3/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M3/M2/_1_  (.A(\V4/A1/A2/A2/M3/s1 ),
    .B(\V4/A1/A2/A2/c2 ),
    .Z(\V4/s1 [14]));
 OR2_X1 \V4/A1/A2/A2/M3/_0_  (.A1(\V4/A1/A2/A2/M3/c1 ),
    .A2(\V4/A1/A2/A2/M3/c2 ),
    .ZN(\V4/A1/A2/A2/c3 ));
 AND2_X1 \V4/A1/A2/A2/M4/M1/_0_  (.A1(\V4/v2 [15]),
    .A2(\V4/v3 [15]),
    .ZN(\V4/A1/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A1/A2/A2/M4/M1/_1_  (.A(\V4/v2 [15]),
    .B(\V4/v3 [15]),
    .Z(\V4/A1/A2/A2/M4/s1 ));
 AND2_X1 \V4/A1/A2/A2/M4/M2/_0_  (.A1(\V4/A1/A2/A2/M4/s1 ),
    .A2(\V4/A1/A2/A2/c3 ),
    .ZN(\V4/A1/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A1/A2/A2/M4/M2/_1_  (.A(\V4/A1/A2/A2/M4/s1 ),
    .B(\V4/A1/A2/A2/c3 ),
    .Z(\V4/s1 [15]));
 OR2_X1 \V4/A1/A2/A2/M4/_0_  (.A1(\V4/A1/A2/A2/M4/c1 ),
    .A2(\V4/A1/A2/A2/M4/c2 ),
    .ZN(\V4/c1 ));
 AND2_X1 \V4/A2/A1/A1/M1/M1/_0_  (.A1(\V4/s1 [0]),
    .A2(\V4/v1 [8]),
    .ZN(\V4/A2/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M1/M1/_1_  (.A(\V4/s1 [0]),
    .B(\V4/v1 [8]),
    .Z(\V4/A2/A1/A1/M1/s1 ));
 AND2_X1 \V4/A2/A1/A1/M1/M2/_0_  (.A1(\V4/A2/A1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/A2/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M1/M2/_1_  (.A(\V4/A2/A1/A1/M1/s1 ),
    .B(net9),
    .Z(v4[8]));
 OR2_X1 \V4/A2/A1/A1/M1/_0_  (.A1(\V4/A2/A1/A1/M1/c1 ),
    .A2(\V4/A2/A1/A1/M1/c2 ),
    .ZN(\V4/A2/A1/A1/c1 ));
 AND2_X1 \V4/A2/A1/A1/M2/M1/_0_  (.A1(\V4/s1 [1]),
    .A2(\V4/v1 [9]),
    .ZN(\V4/A2/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M2/M1/_1_  (.A(\V4/s1 [1]),
    .B(\V4/v1 [9]),
    .Z(\V4/A2/A1/A1/M2/s1 ));
 AND2_X1 \V4/A2/A1/A1/M2/M2/_0_  (.A1(\V4/A2/A1/A1/M2/s1 ),
    .A2(\V4/A2/A1/A1/c1 ),
    .ZN(\V4/A2/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M2/M2/_1_  (.A(\V4/A2/A1/A1/M2/s1 ),
    .B(\V4/A2/A1/A1/c1 ),
    .Z(v4[9]));
 OR2_X1 \V4/A2/A1/A1/M2/_0_  (.A1(\V4/A2/A1/A1/M2/c1 ),
    .A2(\V4/A2/A1/A1/M2/c2 ),
    .ZN(\V4/A2/A1/A1/c2 ));
 AND2_X1 \V4/A2/A1/A1/M3/M1/_0_  (.A1(\V4/s1 [2]),
    .A2(\V4/v1 [10]),
    .ZN(\V4/A2/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M3/M1/_1_  (.A(\V4/s1 [2]),
    .B(\V4/v1 [10]),
    .Z(\V4/A2/A1/A1/M3/s1 ));
 AND2_X1 \V4/A2/A1/A1/M3/M2/_0_  (.A1(\V4/A2/A1/A1/M3/s1 ),
    .A2(\V4/A2/A1/A1/c2 ),
    .ZN(\V4/A2/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M3/M2/_1_  (.A(\V4/A2/A1/A1/M3/s1 ),
    .B(\V4/A2/A1/A1/c2 ),
    .Z(v4[10]));
 OR2_X1 \V4/A2/A1/A1/M3/_0_  (.A1(\V4/A2/A1/A1/M3/c1 ),
    .A2(\V4/A2/A1/A1/M3/c2 ),
    .ZN(\V4/A2/A1/A1/c3 ));
 AND2_X1 \V4/A2/A1/A1/M4/M1/_0_  (.A1(\V4/s1 [3]),
    .A2(\V4/v1 [11]),
    .ZN(\V4/A2/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A2/A1/A1/M4/M1/_1_  (.A(\V4/s1 [3]),
    .B(\V4/v1 [11]),
    .Z(\V4/A2/A1/A1/M4/s1 ));
 AND2_X1 \V4/A2/A1/A1/M4/M2/_0_  (.A1(\V4/A2/A1/A1/M4/s1 ),
    .A2(\V4/A2/A1/A1/c3 ),
    .ZN(\V4/A2/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A2/A1/A1/M4/M2/_1_  (.A(\V4/A2/A1/A1/M4/s1 ),
    .B(\V4/A2/A1/A1/c3 ),
    .Z(v4[11]));
 OR2_X1 \V4/A2/A1/A1/M4/_0_  (.A1(\V4/A2/A1/A1/M4/c1 ),
    .A2(\V4/A2/A1/A1/M4/c2 ),
    .ZN(\V4/A2/A1/c1 ));
 AND2_X1 \V4/A2/A1/A2/M1/M1/_0_  (.A1(\V4/s1 [4]),
    .A2(\V4/v1 [12]),
    .ZN(\V4/A2/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M1/M1/_1_  (.A(\V4/s1 [4]),
    .B(\V4/v1 [12]),
    .Z(\V4/A2/A1/A2/M1/s1 ));
 AND2_X1 \V4/A2/A1/A2/M1/M2/_0_  (.A1(\V4/A2/A1/A2/M1/s1 ),
    .A2(\V4/A2/A1/c1 ),
    .ZN(\V4/A2/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M1/M2/_1_  (.A(\V4/A2/A1/A2/M1/s1 ),
    .B(\V4/A2/A1/c1 ),
    .Z(v4[12]));
 OR2_X1 \V4/A2/A1/A2/M1/_0_  (.A1(\V4/A2/A1/A2/M1/c1 ),
    .A2(\V4/A2/A1/A2/M1/c2 ),
    .ZN(\V4/A2/A1/A2/c1 ));
 AND2_X1 \V4/A2/A1/A2/M2/M1/_0_  (.A1(\V4/s1 [5]),
    .A2(\V4/v1 [13]),
    .ZN(\V4/A2/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M2/M1/_1_  (.A(\V4/s1 [5]),
    .B(\V4/v1 [13]),
    .Z(\V4/A2/A1/A2/M2/s1 ));
 AND2_X1 \V4/A2/A1/A2/M2/M2/_0_  (.A1(\V4/A2/A1/A2/M2/s1 ),
    .A2(\V4/A2/A1/A2/c1 ),
    .ZN(\V4/A2/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M2/M2/_1_  (.A(\V4/A2/A1/A2/M2/s1 ),
    .B(\V4/A2/A1/A2/c1 ),
    .Z(v4[13]));
 OR2_X1 \V4/A2/A1/A2/M2/_0_  (.A1(\V4/A2/A1/A2/M2/c1 ),
    .A2(\V4/A2/A1/A2/M2/c2 ),
    .ZN(\V4/A2/A1/A2/c2 ));
 AND2_X1 \V4/A2/A1/A2/M3/M1/_0_  (.A1(\V4/s1 [6]),
    .A2(\V4/v1 [14]),
    .ZN(\V4/A2/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M3/M1/_1_  (.A(\V4/s1 [6]),
    .B(\V4/v1 [14]),
    .Z(\V4/A2/A1/A2/M3/s1 ));
 AND2_X1 \V4/A2/A1/A2/M3/M2/_0_  (.A1(\V4/A2/A1/A2/M3/s1 ),
    .A2(\V4/A2/A1/A2/c2 ),
    .ZN(\V4/A2/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M3/M2/_1_  (.A(\V4/A2/A1/A2/M3/s1 ),
    .B(\V4/A2/A1/A2/c2 ),
    .Z(v4[14]));
 OR2_X1 \V4/A2/A1/A2/M3/_0_  (.A1(\V4/A2/A1/A2/M3/c1 ),
    .A2(\V4/A2/A1/A2/M3/c2 ),
    .ZN(\V4/A2/A1/A2/c3 ));
 AND2_X1 \V4/A2/A1/A2/M4/M1/_0_  (.A1(\V4/s1 [7]),
    .A2(\V4/v1 [15]),
    .ZN(\V4/A2/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A2/A1/A2/M4/M1/_1_  (.A(\V4/s1 [7]),
    .B(\V4/v1 [15]),
    .Z(\V4/A2/A1/A2/M4/s1 ));
 AND2_X1 \V4/A2/A1/A2/M4/M2/_0_  (.A1(\V4/A2/A1/A2/M4/s1 ),
    .A2(\V4/A2/A1/A2/c3 ),
    .ZN(\V4/A2/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A2/A1/A2/M4/M2/_1_  (.A(\V4/A2/A1/A2/M4/s1 ),
    .B(\V4/A2/A1/A2/c3 ),
    .Z(v4[15]));
 OR2_X1 \V4/A2/A1/A2/M4/_0_  (.A1(\V4/A2/A1/A2/M4/c1 ),
    .A2(\V4/A2/A1/A2/M4/c2 ),
    .ZN(\V4/A2/c1 ));
 AND2_X1 \V4/A2/A2/A1/M1/M1/_0_  (.A1(\V4/s1 [8]),
    .A2(net10),
    .ZN(\V4/A2/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M1/M1/_1_  (.A(\V4/s1 [8]),
    .B(net10),
    .Z(\V4/A2/A2/A1/M1/s1 ));
 AND2_X1 \V4/A2/A2/A1/M1/M2/_0_  (.A1(\V4/A2/A2/A1/M1/s1 ),
    .A2(\V4/A2/c1 ),
    .ZN(\V4/A2/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M1/M2/_1_  (.A(\V4/A2/A2/A1/M1/s1 ),
    .B(\V4/A2/c1 ),
    .Z(\V4/s2 [8]));
 OR2_X1 \V4/A2/A2/A1/M1/_0_  (.A1(\V4/A2/A2/A1/M1/c1 ),
    .A2(\V4/A2/A2/A1/M1/c2 ),
    .ZN(\V4/A2/A2/A1/c1 ));
 AND2_X1 \V4/A2/A2/A1/M2/M1/_0_  (.A1(\V4/s1 [9]),
    .A2(net1),
    .ZN(\V4/A2/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M2/M1/_1_  (.A(\V4/s1 [9]),
    .B(net1),
    .Z(\V4/A2/A2/A1/M2/s1 ));
 AND2_X1 \V4/A2/A2/A1/M2/M2/_0_  (.A1(\V4/A2/A2/A1/M2/s1 ),
    .A2(\V4/A2/A2/A1/c1 ),
    .ZN(\V4/A2/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M2/M2/_1_  (.A(\V4/A2/A2/A1/M2/s1 ),
    .B(\V4/A2/A2/A1/c1 ),
    .Z(\V4/s2 [9]));
 OR2_X1 \V4/A2/A2/A1/M2/_0_  (.A1(\V4/A2/A2/A1/M2/c1 ),
    .A2(\V4/A2/A2/A1/M2/c2 ),
    .ZN(\V4/A2/A2/A1/c2 ));
 AND2_X1 \V4/A2/A2/A1/M3/M1/_0_  (.A1(\V4/s1 [10]),
    .A2(net1),
    .ZN(\V4/A2/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M3/M1/_1_  (.A(\V4/s1 [10]),
    .B(net1),
    .Z(\V4/A2/A2/A1/M3/s1 ));
 AND2_X1 \V4/A2/A2/A1/M3/M2/_0_  (.A1(\V4/A2/A2/A1/M3/s1 ),
    .A2(\V4/A2/A2/A1/c2 ),
    .ZN(\V4/A2/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M3/M2/_1_  (.A(\V4/A2/A2/A1/M3/s1 ),
    .B(\V4/A2/A2/A1/c2 ),
    .Z(\V4/s2 [10]));
 OR2_X1 \V4/A2/A2/A1/M3/_0_  (.A1(\V4/A2/A2/A1/M3/c1 ),
    .A2(\V4/A2/A2/A1/M3/c2 ),
    .ZN(\V4/A2/A2/A1/c3 ));
 AND2_X1 \V4/A2/A2/A1/M4/M1/_0_  (.A1(\V4/s1 [11]),
    .A2(net1),
    .ZN(\V4/A2/A2/A1/M4/c1 ));
 XOR2_X2 \V4/A2/A2/A1/M4/M1/_1_  (.A(\V4/s1 [11]),
    .B(net1),
    .Z(\V4/A2/A2/A1/M4/s1 ));
 AND2_X1 \V4/A2/A2/A1/M4/M2/_0_  (.A1(\V4/A2/A2/A1/M4/s1 ),
    .A2(\V4/A2/A2/A1/c3 ),
    .ZN(\V4/A2/A2/A1/M4/c2 ));
 XOR2_X2 \V4/A2/A2/A1/M4/M2/_1_  (.A(\V4/A2/A2/A1/M4/s1 ),
    .B(\V4/A2/A2/A1/c3 ),
    .Z(\V4/s2 [11]));
 OR2_X1 \V4/A2/A2/A1/M4/_0_  (.A1(\V4/A2/A2/A1/M4/c1 ),
    .A2(\V4/A2/A2/A1/M4/c2 ),
    .ZN(\V4/A2/A2/c1 ));
 AND2_X1 \V4/A2/A2/A2/M1/M1/_0_  (.A1(\V4/s1 [12]),
    .A2(net1),
    .ZN(\V4/A2/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M1/M1/_1_  (.A(\V4/s1 [12]),
    .B(net1),
    .Z(\V4/A2/A2/A2/M1/s1 ));
 AND2_X1 \V4/A2/A2/A2/M1/M2/_0_  (.A1(\V4/A2/A2/A2/M1/s1 ),
    .A2(\V4/A2/A2/c1 ),
    .ZN(\V4/A2/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M1/M2/_1_  (.A(\V4/A2/A2/A2/M1/s1 ),
    .B(\V4/A2/A2/c1 ),
    .Z(\V4/s2 [12]));
 OR2_X1 \V4/A2/A2/A2/M1/_0_  (.A1(\V4/A2/A2/A2/M1/c1 ),
    .A2(\V4/A2/A2/A2/M1/c2 ),
    .ZN(\V4/A2/A2/A2/c1 ));
 AND2_X1 \V4/A2/A2/A2/M2/M1/_0_  (.A1(\V4/s1 [13]),
    .A2(net1),
    .ZN(\V4/A2/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M2/M1/_1_  (.A(\V4/s1 [13]),
    .B(net1),
    .Z(\V4/A2/A2/A2/M2/s1 ));
 AND2_X1 \V4/A2/A2/A2/M2/M2/_0_  (.A1(\V4/A2/A2/A2/M2/s1 ),
    .A2(\V4/A2/A2/A2/c1 ),
    .ZN(\V4/A2/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M2/M2/_1_  (.A(\V4/A2/A2/A2/M2/s1 ),
    .B(\V4/A2/A2/A2/c1 ),
    .Z(\V4/s2 [13]));
 OR2_X1 \V4/A2/A2/A2/M2/_0_  (.A1(\V4/A2/A2/A2/M2/c1 ),
    .A2(\V4/A2/A2/A2/M2/c2 ),
    .ZN(\V4/A2/A2/A2/c2 ));
 AND2_X1 \V4/A2/A2/A2/M3/M1/_0_  (.A1(\V4/s1 [14]),
    .A2(net1),
    .ZN(\V4/A2/A2/A2/M3/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M3/M1/_1_  (.A(\V4/s1 [14]),
    .B(net1),
    .Z(\V4/A2/A2/A2/M3/s1 ));
 AND2_X1 \V4/A2/A2/A2/M3/M2/_0_  (.A1(\V4/A2/A2/A2/M3/s1 ),
    .A2(\V4/A2/A2/A2/c2 ),
    .ZN(\V4/A2/A2/A2/M3/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M3/M2/_1_  (.A(\V4/A2/A2/A2/M3/s1 ),
    .B(\V4/A2/A2/A2/c2 ),
    .Z(\V4/s2 [14]));
 OR2_X1 \V4/A2/A2/A2/M3/_0_  (.A1(\V4/A2/A2/A2/M3/c1 ),
    .A2(\V4/A2/A2/A2/M3/c2 ),
    .ZN(\V4/A2/A2/A2/c3 ));
 AND2_X1 \V4/A2/A2/A2/M4/M1/_0_  (.A1(\V4/s1 [15]),
    .A2(net1),
    .ZN(\V4/A2/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A2/A2/A2/M4/M1/_1_  (.A(\V4/s1 [15]),
    .B(net1),
    .Z(\V4/A2/A2/A2/M4/s1 ));
 AND2_X1 \V4/A2/A2/A2/M4/M2/_0_  (.A1(\V4/A2/A2/A2/M4/s1 ),
    .A2(\V4/A2/A2/A2/c3 ),
    .ZN(\V4/A2/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A2/A2/A2/M4/M2/_1_  (.A(\V4/A2/A2/A2/M4/s1 ),
    .B(\V4/A2/A2/A2/c3 ),
    .Z(\V4/s2 [15]));
 OR2_X1 \V4/A2/A2/A2/M4/_0_  (.A1(\V4/A2/A2/A2/M4/c1 ),
    .A2(\V4/A2/A2/A2/M4/c2 ),
    .ZN(\V4/c2 ));
 AND2_X1 \V4/A3/A1/A1/M1/M1/_0_  (.A1(\V4/v4 [0]),
    .A2(\V4/s2 [8]),
    .ZN(\V4/A3/A1/A1/M1/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M1/M1/_1_  (.A(\V4/v4 [0]),
    .B(\V4/s2 [8]),
    .Z(\V4/A3/A1/A1/M1/s1 ));
 AND2_X1 \V4/A3/A1/A1/M1/M2/_0_  (.A1(\V4/A3/A1/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/A3/A1/A1/M1/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M1/M2/_1_  (.A(\V4/A3/A1/A1/M1/s1 ),
    .B(net1),
    .Z(v4[16]));
 OR2_X1 \V4/A3/A1/A1/M1/_0_  (.A1(\V4/A3/A1/A1/M1/c1 ),
    .A2(\V4/A3/A1/A1/M1/c2 ),
    .ZN(\V4/A3/A1/A1/c1 ));
 AND2_X1 \V4/A3/A1/A1/M2/M1/_0_  (.A1(\V4/v4 [1]),
    .A2(\V4/s2 [9]),
    .ZN(\V4/A3/A1/A1/M2/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M2/M1/_1_  (.A(\V4/v4 [1]),
    .B(\V4/s2 [9]),
    .Z(\V4/A3/A1/A1/M2/s1 ));
 AND2_X1 \V4/A3/A1/A1/M2/M2/_0_  (.A1(\V4/A3/A1/A1/M2/s1 ),
    .A2(\V4/A3/A1/A1/c1 ),
    .ZN(\V4/A3/A1/A1/M2/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M2/M2/_1_  (.A(\V4/A3/A1/A1/M2/s1 ),
    .B(\V4/A3/A1/A1/c1 ),
    .Z(v4[17]));
 OR2_X1 \V4/A3/A1/A1/M2/_0_  (.A1(\V4/A3/A1/A1/M2/c1 ),
    .A2(\V4/A3/A1/A1/M2/c2 ),
    .ZN(\V4/A3/A1/A1/c2 ));
 AND2_X1 \V4/A3/A1/A1/M3/M1/_0_  (.A1(\V4/v4 [2]),
    .A2(\V4/s2 [10]),
    .ZN(\V4/A3/A1/A1/M3/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M3/M1/_1_  (.A(\V4/v4 [2]),
    .B(\V4/s2 [10]),
    .Z(\V4/A3/A1/A1/M3/s1 ));
 AND2_X1 \V4/A3/A1/A1/M3/M2/_0_  (.A1(\V4/A3/A1/A1/M3/s1 ),
    .A2(\V4/A3/A1/A1/c2 ),
    .ZN(\V4/A3/A1/A1/M3/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M3/M2/_1_  (.A(\V4/A3/A1/A1/M3/s1 ),
    .B(\V4/A3/A1/A1/c2 ),
    .Z(v4[18]));
 OR2_X1 \V4/A3/A1/A1/M3/_0_  (.A1(\V4/A3/A1/A1/M3/c1 ),
    .A2(\V4/A3/A1/A1/M3/c2 ),
    .ZN(\V4/A3/A1/A1/c3 ));
 AND2_X1 \V4/A3/A1/A1/M4/M1/_0_  (.A1(\V4/v4 [3]),
    .A2(\V4/s2 [11]),
    .ZN(\V4/A3/A1/A1/M4/c1 ));
 XOR2_X2 \V4/A3/A1/A1/M4/M1/_1_  (.A(\V4/v4 [3]),
    .B(\V4/s2 [11]),
    .Z(\V4/A3/A1/A1/M4/s1 ));
 AND2_X1 \V4/A3/A1/A1/M4/M2/_0_  (.A1(\V4/A3/A1/A1/M4/s1 ),
    .A2(\V4/A3/A1/A1/c3 ),
    .ZN(\V4/A3/A1/A1/M4/c2 ));
 XOR2_X2 \V4/A3/A1/A1/M4/M2/_1_  (.A(\V4/A3/A1/A1/M4/s1 ),
    .B(\V4/A3/A1/A1/c3 ),
    .Z(v4[19]));
 OR2_X1 \V4/A3/A1/A1/M4/_0_  (.A1(\V4/A3/A1/A1/M4/c1 ),
    .A2(\V4/A3/A1/A1/M4/c2 ),
    .ZN(\V4/A3/A1/c1 ));
 AND2_X1 \V4/A3/A1/A2/M1/M1/_0_  (.A1(\V4/v4 [4]),
    .A2(\V4/s2 [12]),
    .ZN(\V4/A3/A1/A2/M1/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M1/M1/_1_  (.A(\V4/v4 [4]),
    .B(\V4/s2 [12]),
    .Z(\V4/A3/A1/A2/M1/s1 ));
 AND2_X1 \V4/A3/A1/A2/M1/M2/_0_  (.A1(\V4/A3/A1/A2/M1/s1 ),
    .A2(\V4/A3/A1/c1 ),
    .ZN(\V4/A3/A1/A2/M1/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M1/M2/_1_  (.A(\V4/A3/A1/A2/M1/s1 ),
    .B(\V4/A3/A1/c1 ),
    .Z(v4[20]));
 OR2_X1 \V4/A3/A1/A2/M1/_0_  (.A1(\V4/A3/A1/A2/M1/c1 ),
    .A2(\V4/A3/A1/A2/M1/c2 ),
    .ZN(\V4/A3/A1/A2/c1 ));
 AND2_X1 \V4/A3/A1/A2/M2/M1/_0_  (.A1(\V4/v4 [5]),
    .A2(\V4/s2 [13]),
    .ZN(\V4/A3/A1/A2/M2/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M2/M1/_1_  (.A(\V4/v4 [5]),
    .B(\V4/s2 [13]),
    .Z(\V4/A3/A1/A2/M2/s1 ));
 AND2_X1 \V4/A3/A1/A2/M2/M2/_0_  (.A1(\V4/A3/A1/A2/M2/s1 ),
    .A2(\V4/A3/A1/A2/c1 ),
    .ZN(\V4/A3/A1/A2/M2/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M2/M2/_1_  (.A(\V4/A3/A1/A2/M2/s1 ),
    .B(\V4/A3/A1/A2/c1 ),
    .Z(v4[21]));
 OR2_X1 \V4/A3/A1/A2/M2/_0_  (.A1(\V4/A3/A1/A2/M2/c1 ),
    .A2(\V4/A3/A1/A2/M2/c2 ),
    .ZN(\V4/A3/A1/A2/c2 ));
 AND2_X1 \V4/A3/A1/A2/M3/M1/_0_  (.A1(\V4/v4 [6]),
    .A2(\V4/s2 [14]),
    .ZN(\V4/A3/A1/A2/M3/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M3/M1/_1_  (.A(\V4/v4 [6]),
    .B(\V4/s2 [14]),
    .Z(\V4/A3/A1/A2/M3/s1 ));
 AND2_X1 \V4/A3/A1/A2/M3/M2/_0_  (.A1(\V4/A3/A1/A2/M3/s1 ),
    .A2(\V4/A3/A1/A2/c2 ),
    .ZN(\V4/A3/A1/A2/M3/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M3/M2/_1_  (.A(\V4/A3/A1/A2/M3/s1 ),
    .B(\V4/A3/A1/A2/c2 ),
    .Z(v4[22]));
 OR2_X1 \V4/A3/A1/A2/M3/_0_  (.A1(\V4/A3/A1/A2/M3/c1 ),
    .A2(\V4/A3/A1/A2/M3/c2 ),
    .ZN(\V4/A3/A1/A2/c3 ));
 AND2_X1 \V4/A3/A1/A2/M4/M1/_0_  (.A1(\V4/v4 [7]),
    .A2(\V4/s2 [15]),
    .ZN(\V4/A3/A1/A2/M4/c1 ));
 XOR2_X2 \V4/A3/A1/A2/M4/M1/_1_  (.A(\V4/v4 [7]),
    .B(\V4/s2 [15]),
    .Z(\V4/A3/A1/A2/M4/s1 ));
 AND2_X1 \V4/A3/A1/A2/M4/M2/_0_  (.A1(\V4/A3/A1/A2/M4/s1 ),
    .A2(\V4/A3/A1/A2/c3 ),
    .ZN(\V4/A3/A1/A2/M4/c2 ));
 XOR2_X2 \V4/A3/A1/A2/M4/M2/_1_  (.A(\V4/A3/A1/A2/M4/s1 ),
    .B(\V4/A3/A1/A2/c3 ),
    .Z(v4[23]));
 OR2_X1 \V4/A3/A1/A2/M4/_0_  (.A1(\V4/A3/A1/A2/M4/c1 ),
    .A2(\V4/A3/A1/A2/M4/c2 ),
    .ZN(\V4/A3/c1 ));
 AND2_X1 \V4/A3/A2/A1/M1/M1/_0_  (.A1(\V4/v4 [8]),
    .A2(\V4/c3 ),
    .ZN(\V4/A3/A2/A1/M1/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M1/M1/_1_  (.A(\V4/v4 [8]),
    .B(\V4/c3 ),
    .Z(\V4/A3/A2/A1/M1/s1 ));
 AND2_X1 \V4/A3/A2/A1/M1/M2/_0_  (.A1(\V4/A3/A2/A1/M1/s1 ),
    .A2(\V4/A3/c1 ),
    .ZN(\V4/A3/A2/A1/M1/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M1/M2/_1_  (.A(\V4/A3/A2/A1/M1/s1 ),
    .B(\V4/A3/c1 ),
    .Z(v4[24]));
 OR2_X1 \V4/A3/A2/A1/M1/_0_  (.A1(\V4/A3/A2/A1/M1/c1 ),
    .A2(\V4/A3/A2/A1/M1/c2 ),
    .ZN(\V4/A3/A2/A1/c1 ));
 AND2_X1 \V4/A3/A2/A1/M2/M1/_0_  (.A1(\V4/v4 [9]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M2/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M2/M1/_1_  (.A(\V4/v4 [9]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M2/s1 ));
 AND2_X1 \V4/A3/A2/A1/M2/M2/_0_  (.A1(\V4/A3/A2/A1/M2/s1 ),
    .A2(\V4/A3/A2/A1/c1 ),
    .ZN(\V4/A3/A2/A1/M2/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M2/M2/_1_  (.A(\V4/A3/A2/A1/M2/s1 ),
    .B(\V4/A3/A2/A1/c1 ),
    .Z(v4[25]));
 OR2_X1 \V4/A3/A2/A1/M2/_0_  (.A1(\V4/A3/A2/A1/M2/c1 ),
    .A2(\V4/A3/A2/A1/M2/c2 ),
    .ZN(\V4/A3/A2/A1/c2 ));
 AND2_X1 \V4/A3/A2/A1/M3/M1/_0_  (.A1(\V4/v4 [10]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M3/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M3/M1/_1_  (.A(\V4/v4 [10]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M3/s1 ));
 AND2_X1 \V4/A3/A2/A1/M3/M2/_0_  (.A1(\V4/A3/A2/A1/M3/s1 ),
    .A2(\V4/A3/A2/A1/c2 ),
    .ZN(\V4/A3/A2/A1/M3/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M3/M2/_1_  (.A(\V4/A3/A2/A1/M3/s1 ),
    .B(\V4/A3/A2/A1/c2 ),
    .Z(v4[26]));
 OR2_X1 \V4/A3/A2/A1/M3/_0_  (.A1(\V4/A3/A2/A1/M3/c1 ),
    .A2(\V4/A3/A2/A1/M3/c2 ),
    .ZN(\V4/A3/A2/A1/c3 ));
 AND2_X1 \V4/A3/A2/A1/M4/M1/_0_  (.A1(\V4/v4 [11]),
    .A2(ground),
    .ZN(\V4/A3/A2/A1/M4/c1 ));
 XOR2_X2 \V4/A3/A2/A1/M4/M1/_1_  (.A(\V4/v4 [11]),
    .B(ground),
    .Z(\V4/A3/A2/A1/M4/s1 ));
 AND2_X1 \V4/A3/A2/A1/M4/M2/_0_  (.A1(\V4/A3/A2/A1/M4/s1 ),
    .A2(\V4/A3/A2/A1/c3 ),
    .ZN(\V4/A3/A2/A1/M4/c2 ));
 XOR2_X2 \V4/A3/A2/A1/M4/M2/_1_  (.A(\V4/A3/A2/A1/M4/s1 ),
    .B(\V4/A3/A2/A1/c3 ),
    .Z(v4[27]));
 OR2_X1 \V4/A3/A2/A1/M4/_0_  (.A1(\V4/A3/A2/A1/M4/c1 ),
    .A2(\V4/A3/A2/A1/M4/c2 ),
    .ZN(\V4/A3/A2/c1 ));
 AND2_X1 \V4/A3/A2/A2/M1/M1/_0_  (.A1(\V4/v4 [12]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M1/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M1/M1/_1_  (.A(\V4/v4 [12]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M1/s1 ));
 AND2_X1 \V4/A3/A2/A2/M1/M2/_0_  (.A1(\V4/A3/A2/A2/M1/s1 ),
    .A2(\V4/A3/A2/c1 ),
    .ZN(\V4/A3/A2/A2/M1/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M1/M2/_1_  (.A(\V4/A3/A2/A2/M1/s1 ),
    .B(\V4/A3/A2/c1 ),
    .Z(v4[28]));
 OR2_X1 \V4/A3/A2/A2/M1/_0_  (.A1(\V4/A3/A2/A2/M1/c1 ),
    .A2(\V4/A3/A2/A2/M1/c2 ),
    .ZN(\V4/A3/A2/A2/c1 ));
 AND2_X1 \V4/A3/A2/A2/M2/M1/_0_  (.A1(\V4/v4 [13]),
    .A2(net10),
    .ZN(\V4/A3/A2/A2/M2/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M2/M1/_1_  (.A(\V4/v4 [13]),
    .B(net10),
    .Z(\V4/A3/A2/A2/M2/s1 ));
 AND2_X1 \V4/A3/A2/A2/M2/M2/_0_  (.A1(\V4/A3/A2/A2/M2/s1 ),
    .A2(\V4/A3/A2/A2/c1 ),
    .ZN(\V4/A3/A2/A2/M2/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M2/M2/_1_  (.A(\V4/A3/A2/A2/M2/s1 ),
    .B(\V4/A3/A2/A2/c1 ),
    .Z(v4[29]));
 OR2_X1 \V4/A3/A2/A2/M2/_0_  (.A1(\V4/A3/A2/A2/M2/c1 ),
    .A2(\V4/A3/A2/A2/M2/c2 ),
    .ZN(\V4/A3/A2/A2/c2 ));
 AND2_X1 \V4/A3/A2/A2/M3/M1/_0_  (.A1(\V4/v4 [14]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M3/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M3/M1/_1_  (.A(\V4/v4 [14]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M3/s1 ));
 AND2_X1 \V4/A3/A2/A2/M3/M2/_0_  (.A1(\V4/A3/A2/A2/M3/s1 ),
    .A2(\V4/A3/A2/A2/c2 ),
    .ZN(\V4/A3/A2/A2/M3/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M3/M2/_1_  (.A(\V4/A3/A2/A2/M3/s1 ),
    .B(\V4/A3/A2/A2/c2 ),
    .Z(v4[30]));
 OR2_X1 \V4/A3/A2/A2/M3/_0_  (.A1(\V4/A3/A2/A2/M3/c1 ),
    .A2(\V4/A3/A2/A2/M3/c2 ),
    .ZN(\V4/A3/A2/A2/c3 ));
 AND2_X1 \V4/A3/A2/A2/M4/M1/_0_  (.A1(\V4/v4 [15]),
    .A2(ground),
    .ZN(\V4/A3/A2/A2/M4/c1 ));
 XOR2_X2 \V4/A3/A2/A2/M4/M1/_1_  (.A(\V4/v4 [15]),
    .B(ground),
    .Z(\V4/A3/A2/A2/M4/s1 ));
 AND2_X1 \V4/A3/A2/A2/M4/M2/_0_  (.A1(\V4/A3/A2/A2/M4/s1 ),
    .A2(\V4/A3/A2/A2/c3 ),
    .ZN(\V4/A3/A2/A2/M4/c2 ));
 XOR2_X2 \V4/A3/A2/A2/M4/M2/_1_  (.A(\V4/A3/A2/A2/M4/s1 ),
    .B(\V4/A3/A2/A2/c3 ),
    .Z(v4[31]));
 OR2_X1 \V4/A3/A2/A2/M4/_0_  (.A1(\V4/A3/A2/A2/M4/c1 ),
    .A2(\V4/A3/A2/A2/M4/c2 ),
    .ZN(\V4/overflow ));
 AND2_X1 \V4/V1/A1/A1/M1/M1/_0_  (.A1(\V4/V1/v2 [0]),
    .A2(\V4/V1/v3 [0]),
    .ZN(\V4/V1/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M1/M1/_1_  (.A(\V4/V1/v2 [0]),
    .B(\V4/V1/v3 [0]),
    .Z(\V4/V1/A1/A1/M1/s1 ));
 AND2_X1 \V4/V1/A1/A1/M1/M2/_0_  (.A1(\V4/V1/A1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M1/M2/_1_  (.A(\V4/V1/A1/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/V1/s1 [0]));
 OR2_X1 \V4/V1/A1/A1/M1/_0_  (.A1(\V4/V1/A1/A1/M1/c1 ),
    .A2(\V4/V1/A1/A1/M1/c2 ),
    .ZN(\V4/V1/A1/A1/c1 ));
 AND2_X1 \V4/V1/A1/A1/M2/M1/_0_  (.A1(\V4/V1/v2 [1]),
    .A2(\V4/V1/v3 [1]),
    .ZN(\V4/V1/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M2/M1/_1_  (.A(\V4/V1/v2 [1]),
    .B(\V4/V1/v3 [1]),
    .Z(\V4/V1/A1/A1/M2/s1 ));
 AND2_X1 \V4/V1/A1/A1/M2/M2/_0_  (.A1(\V4/V1/A1/A1/M2/s1 ),
    .A2(\V4/V1/A1/A1/c1 ),
    .ZN(\V4/V1/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M2/M2/_1_  (.A(\V4/V1/A1/A1/M2/s1 ),
    .B(\V4/V1/A1/A1/c1 ),
    .Z(\V4/V1/s1 [1]));
 OR2_X1 \V4/V1/A1/A1/M2/_0_  (.A1(\V4/V1/A1/A1/M2/c1 ),
    .A2(\V4/V1/A1/A1/M2/c2 ),
    .ZN(\V4/V1/A1/A1/c2 ));
 AND2_X1 \V4/V1/A1/A1/M3/M1/_0_  (.A1(\V4/V1/v2 [2]),
    .A2(\V4/V1/v3 [2]),
    .ZN(\V4/V1/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M3/M1/_1_  (.A(\V4/V1/v2 [2]),
    .B(\V4/V1/v3 [2]),
    .Z(\V4/V1/A1/A1/M3/s1 ));
 AND2_X1 \V4/V1/A1/A1/M3/M2/_0_  (.A1(\V4/V1/A1/A1/M3/s1 ),
    .A2(\V4/V1/A1/A1/c2 ),
    .ZN(\V4/V1/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M3/M2/_1_  (.A(\V4/V1/A1/A1/M3/s1 ),
    .B(\V4/V1/A1/A1/c2 ),
    .Z(\V4/V1/s1 [2]));
 OR2_X1 \V4/V1/A1/A1/M3/_0_  (.A1(\V4/V1/A1/A1/M3/c1 ),
    .A2(\V4/V1/A1/A1/M3/c2 ),
    .ZN(\V4/V1/A1/A1/c3 ));
 AND2_X1 \V4/V1/A1/A1/M4/M1/_0_  (.A1(\V4/V1/v2 [3]),
    .A2(\V4/V1/v3 [3]),
    .ZN(\V4/V1/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A1/A1/M4/M1/_1_  (.A(\V4/V1/v2 [3]),
    .B(\V4/V1/v3 [3]),
    .Z(\V4/V1/A1/A1/M4/s1 ));
 AND2_X1 \V4/V1/A1/A1/M4/M2/_0_  (.A1(\V4/V1/A1/A1/M4/s1 ),
    .A2(\V4/V1/A1/A1/c3 ),
    .ZN(\V4/V1/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A1/A1/M4/M2/_1_  (.A(\V4/V1/A1/A1/M4/s1 ),
    .B(\V4/V1/A1/A1/c3 ),
    .Z(\V4/V1/s1 [3]));
 OR2_X1 \V4/V1/A1/A1/M4/_0_  (.A1(\V4/V1/A1/A1/M4/c1 ),
    .A2(\V4/V1/A1/A1/M4/c2 ),
    .ZN(\V4/V1/A1/c1 ));
 AND2_X1 \V4/V1/A1/A2/M1/M1/_0_  (.A1(\V4/V1/v2 [4]),
    .A2(\V4/V1/v3 [4]),
    .ZN(\V4/V1/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M1/M1/_1_  (.A(\V4/V1/v2 [4]),
    .B(\V4/V1/v3 [4]),
    .Z(\V4/V1/A1/A2/M1/s1 ));
 AND2_X1 \V4/V1/A1/A2/M1/M2/_0_  (.A1(\V4/V1/A1/A2/M1/s1 ),
    .A2(\V4/V1/A1/c1 ),
    .ZN(\V4/V1/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M1/M2/_1_  (.A(\V4/V1/A1/A2/M1/s1 ),
    .B(\V4/V1/A1/c1 ),
    .Z(\V4/V1/s1 [4]));
 OR2_X1 \V4/V1/A1/A2/M1/_0_  (.A1(\V4/V1/A1/A2/M1/c1 ),
    .A2(\V4/V1/A1/A2/M1/c2 ),
    .ZN(\V4/V1/A1/A2/c1 ));
 AND2_X1 \V4/V1/A1/A2/M2/M1/_0_  (.A1(\V4/V1/v2 [5]),
    .A2(\V4/V1/v3 [5]),
    .ZN(\V4/V1/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M2/M1/_1_  (.A(\V4/V1/v2 [5]),
    .B(\V4/V1/v3 [5]),
    .Z(\V4/V1/A1/A2/M2/s1 ));
 AND2_X1 \V4/V1/A1/A2/M2/M2/_0_  (.A1(\V4/V1/A1/A2/M2/s1 ),
    .A2(\V4/V1/A1/A2/c1 ),
    .ZN(\V4/V1/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M2/M2/_1_  (.A(\V4/V1/A1/A2/M2/s1 ),
    .B(\V4/V1/A1/A2/c1 ),
    .Z(\V4/V1/s1 [5]));
 OR2_X1 \V4/V1/A1/A2/M2/_0_  (.A1(\V4/V1/A1/A2/M2/c1 ),
    .A2(\V4/V1/A1/A2/M2/c2 ),
    .ZN(\V4/V1/A1/A2/c2 ));
 AND2_X1 \V4/V1/A1/A2/M3/M1/_0_  (.A1(\V4/V1/v2 [6]),
    .A2(\V4/V1/v3 [6]),
    .ZN(\V4/V1/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M3/M1/_1_  (.A(\V4/V1/v2 [6]),
    .B(\V4/V1/v3 [6]),
    .Z(\V4/V1/A1/A2/M3/s1 ));
 AND2_X1 \V4/V1/A1/A2/M3/M2/_0_  (.A1(\V4/V1/A1/A2/M3/s1 ),
    .A2(\V4/V1/A1/A2/c2 ),
    .ZN(\V4/V1/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M3/M2/_1_  (.A(\V4/V1/A1/A2/M3/s1 ),
    .B(\V4/V1/A1/A2/c2 ),
    .Z(\V4/V1/s1 [6]));
 OR2_X1 \V4/V1/A1/A2/M3/_0_  (.A1(\V4/V1/A1/A2/M3/c1 ),
    .A2(\V4/V1/A1/A2/M3/c2 ),
    .ZN(\V4/V1/A1/A2/c3 ));
 AND2_X1 \V4/V1/A1/A2/M4/M1/_0_  (.A1(\V4/V1/v2 [7]),
    .A2(\V4/V1/v3 [7]),
    .ZN(\V4/V1/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A1/A2/M4/M1/_1_  (.A(\V4/V1/v2 [7]),
    .B(\V4/V1/v3 [7]),
    .Z(\V4/V1/A1/A2/M4/s1 ));
 AND2_X1 \V4/V1/A1/A2/M4/M2/_0_  (.A1(\V4/V1/A1/A2/M4/s1 ),
    .A2(\V4/V1/A1/A2/c3 ),
    .ZN(\V4/V1/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A1/A2/M4/M2/_1_  (.A(\V4/V1/A1/A2/M4/s1 ),
    .B(\V4/V1/A1/A2/c3 ),
    .Z(\V4/V1/s1 [7]));
 OR2_X1 \V4/V1/A1/A2/M4/_0_  (.A1(\V4/V1/A1/A2/M4/c1 ),
    .A2(\V4/V1/A1/A2/M4/c2 ),
    .ZN(\V4/V1/c1 ));
 AND2_X1 \V4/V1/A2/A1/M1/M1/_0_  (.A1(\V4/V1/s1 [0]),
    .A2(\V4/V1/v1 [4]),
    .ZN(\V4/V1/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M1/M1/_1_  (.A(\V4/V1/s1 [0]),
    .B(\V4/V1/v1 [4]),
    .Z(\V4/V1/A2/A1/M1/s1 ));
 AND2_X1 \V4/V1/A2/A1/M1/M2/_0_  (.A1(\V4/V1/A2/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M1/M2/_1_  (.A(\V4/V1/A2/A1/M1/s1 ),
    .B(net9),
    .Z(v4[4]));
 OR2_X1 \V4/V1/A2/A1/M1/_0_  (.A1(\V4/V1/A2/A1/M1/c1 ),
    .A2(\V4/V1/A2/A1/M1/c2 ),
    .ZN(\V4/V1/A2/A1/c1 ));
 AND2_X1 \V4/V1/A2/A1/M2/M1/_0_  (.A1(\V4/V1/s1 [1]),
    .A2(\V4/V1/v1 [5]),
    .ZN(\V4/V1/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M2/M1/_1_  (.A(\V4/V1/s1 [1]),
    .B(\V4/V1/v1 [5]),
    .Z(\V4/V1/A2/A1/M2/s1 ));
 AND2_X1 \V4/V1/A2/A1/M2/M2/_0_  (.A1(\V4/V1/A2/A1/M2/s1 ),
    .A2(\V4/V1/A2/A1/c1 ),
    .ZN(\V4/V1/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M2/M2/_1_  (.A(\V4/V1/A2/A1/M2/s1 ),
    .B(\V4/V1/A2/A1/c1 ),
    .Z(v4[5]));
 OR2_X1 \V4/V1/A2/A1/M2/_0_  (.A1(\V4/V1/A2/A1/M2/c1 ),
    .A2(\V4/V1/A2/A1/M2/c2 ),
    .ZN(\V4/V1/A2/A1/c2 ));
 AND2_X1 \V4/V1/A2/A1/M3/M1/_0_  (.A1(\V4/V1/s1 [2]),
    .A2(\V4/V1/v1 [6]),
    .ZN(\V4/V1/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M3/M1/_1_  (.A(\V4/V1/s1 [2]),
    .B(\V4/V1/v1 [6]),
    .Z(\V4/V1/A2/A1/M3/s1 ));
 AND2_X1 \V4/V1/A2/A1/M3/M2/_0_  (.A1(\V4/V1/A2/A1/M3/s1 ),
    .A2(\V4/V1/A2/A1/c2 ),
    .ZN(\V4/V1/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M3/M2/_1_  (.A(\V4/V1/A2/A1/M3/s1 ),
    .B(\V4/V1/A2/A1/c2 ),
    .Z(v4[6]));
 OR2_X1 \V4/V1/A2/A1/M3/_0_  (.A1(\V4/V1/A2/A1/M3/c1 ),
    .A2(\V4/V1/A2/A1/M3/c2 ),
    .ZN(\V4/V1/A2/A1/c3 ));
 AND2_X1 \V4/V1/A2/A1/M4/M1/_0_  (.A1(\V4/V1/s1 [3]),
    .A2(\V4/V1/v1 [7]),
    .ZN(\V4/V1/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A2/A1/M4/M1/_1_  (.A(\V4/V1/s1 [3]),
    .B(\V4/V1/v1 [7]),
    .Z(\V4/V1/A2/A1/M4/s1 ));
 AND2_X1 \V4/V1/A2/A1/M4/M2/_0_  (.A1(\V4/V1/A2/A1/M4/s1 ),
    .A2(\V4/V1/A2/A1/c3 ),
    .ZN(\V4/V1/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A2/A1/M4/M2/_1_  (.A(\V4/V1/A2/A1/M4/s1 ),
    .B(\V4/V1/A2/A1/c3 ),
    .Z(v4[7]));
 OR2_X1 \V4/V1/A2/A1/M4/_0_  (.A1(\V4/V1/A2/A1/M4/c1 ),
    .A2(\V4/V1/A2/A1/M4/c2 ),
    .ZN(\V4/V1/A2/c1 ));
 AND2_X1 \V4/V1/A2/A2/M1/M1/_0_  (.A1(\V4/V1/s1 [4]),
    .A2(net10),
    .ZN(\V4/V1/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M1/M1/_1_  (.A(\V4/V1/s1 [4]),
    .B(net10),
    .Z(\V4/V1/A2/A2/M1/s1 ));
 AND2_X1 \V4/V1/A2/A2/M1/M2/_0_  (.A1(\V4/V1/A2/A2/M1/s1 ),
    .A2(\V4/V1/A2/c1 ),
    .ZN(\V4/V1/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M1/M2/_1_  (.A(\V4/V1/A2/A2/M1/s1 ),
    .B(\V4/V1/A2/c1 ),
    .Z(\V4/V1/s2 [4]));
 OR2_X1 \V4/V1/A2/A2/M1/_0_  (.A1(\V4/V1/A2/A2/M1/c1 ),
    .A2(\V4/V1/A2/A2/M1/c2 ),
    .ZN(\V4/V1/A2/A2/c1 ));
 AND2_X1 \V4/V1/A2/A2/M2/M1/_0_  (.A1(\V4/V1/s1 [5]),
    .A2(net10),
    .ZN(\V4/V1/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M2/M1/_1_  (.A(\V4/V1/s1 [5]),
    .B(net10),
    .Z(\V4/V1/A2/A2/M2/s1 ));
 AND2_X1 \V4/V1/A2/A2/M2/M2/_0_  (.A1(\V4/V1/A2/A2/M2/s1 ),
    .A2(\V4/V1/A2/A2/c1 ),
    .ZN(\V4/V1/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M2/M2/_1_  (.A(\V4/V1/A2/A2/M2/s1 ),
    .B(\V4/V1/A2/A2/c1 ),
    .Z(\V4/V1/s2 [5]));
 OR2_X1 \V4/V1/A2/A2/M2/_0_  (.A1(\V4/V1/A2/A2/M2/c1 ),
    .A2(\V4/V1/A2/A2/M2/c2 ),
    .ZN(\V4/V1/A2/A2/c2 ));
 AND2_X1 \V4/V1/A2/A2/M3/M1/_0_  (.A1(\V4/V1/s1 [6]),
    .A2(net10),
    .ZN(\V4/V1/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M3/M1/_1_  (.A(\V4/V1/s1 [6]),
    .B(net10),
    .Z(\V4/V1/A2/A2/M3/s1 ));
 AND2_X1 \V4/V1/A2/A2/M3/M2/_0_  (.A1(\V4/V1/A2/A2/M3/s1 ),
    .A2(\V4/V1/A2/A2/c2 ),
    .ZN(\V4/V1/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M3/M2/_1_  (.A(\V4/V1/A2/A2/M3/s1 ),
    .B(\V4/V1/A2/A2/c2 ),
    .Z(\V4/V1/s2 [6]));
 OR2_X1 \V4/V1/A2/A2/M3/_0_  (.A1(\V4/V1/A2/A2/M3/c1 ),
    .A2(\V4/V1/A2/A2/M3/c2 ),
    .ZN(\V4/V1/A2/A2/c3 ));
 AND2_X1 \V4/V1/A2/A2/M4/M1/_0_  (.A1(\V4/V1/s1 [7]),
    .A2(net1),
    .ZN(\V4/V1/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A2/A2/M4/M1/_1_  (.A(\V4/V1/s1 [7]),
    .B(net1),
    .Z(\V4/V1/A2/A2/M4/s1 ));
 AND2_X1 \V4/V1/A2/A2/M4/M2/_0_  (.A1(\V4/V1/A2/A2/M4/s1 ),
    .A2(\V4/V1/A2/A2/c3 ),
    .ZN(\V4/V1/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A2/A2/M4/M2/_1_  (.A(\V4/V1/A2/A2/M4/s1 ),
    .B(\V4/V1/A2/A2/c3 ),
    .Z(\V4/V1/s2 [7]));
 OR2_X1 \V4/V1/A2/A2/M4/_0_  (.A1(\V4/V1/A2/A2/M4/c1 ),
    .A2(\V4/V1/A2/A2/M4/c2 ),
    .ZN(\V4/V1/c2 ));
 AND2_X1 \V4/V1/A3/A1/M1/M1/_0_  (.A1(\V4/V1/v4 [0]),
    .A2(\V4/V1/s2 [4]),
    .ZN(\V4/V1/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M1/M1/_1_  (.A(\V4/V1/v4 [0]),
    .B(\V4/V1/s2 [4]),
    .Z(\V4/V1/A3/A1/M1/s1 ));
 AND2_X1 \V4/V1/A3/A1/M1/M2/_0_  (.A1(\V4/V1/A3/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M1/M2/_1_  (.A(\V4/V1/A3/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/v1 [8]));
 OR2_X1 \V4/V1/A3/A1/M1/_0_  (.A1(\V4/V1/A3/A1/M1/c1 ),
    .A2(\V4/V1/A3/A1/M1/c2 ),
    .ZN(\V4/V1/A3/A1/c1 ));
 AND2_X1 \V4/V1/A3/A1/M2/M1/_0_  (.A1(\V4/V1/v4 [1]),
    .A2(\V4/V1/s2 [5]),
    .ZN(\V4/V1/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M2/M1/_1_  (.A(\V4/V1/v4 [1]),
    .B(\V4/V1/s2 [5]),
    .Z(\V4/V1/A3/A1/M2/s1 ));
 AND2_X1 \V4/V1/A3/A1/M2/M2/_0_  (.A1(\V4/V1/A3/A1/M2/s1 ),
    .A2(\V4/V1/A3/A1/c1 ),
    .ZN(\V4/V1/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M2/M2/_1_  (.A(\V4/V1/A3/A1/M2/s1 ),
    .B(\V4/V1/A3/A1/c1 ),
    .Z(\V4/v1 [9]));
 OR2_X1 \V4/V1/A3/A1/M2/_0_  (.A1(\V4/V1/A3/A1/M2/c1 ),
    .A2(\V4/V1/A3/A1/M2/c2 ),
    .ZN(\V4/V1/A3/A1/c2 ));
 AND2_X1 \V4/V1/A3/A1/M3/M1/_0_  (.A1(\V4/V1/v4 [2]),
    .A2(\V4/V1/s2 [6]),
    .ZN(\V4/V1/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M3/M1/_1_  (.A(\V4/V1/v4 [2]),
    .B(\V4/V1/s2 [6]),
    .Z(\V4/V1/A3/A1/M3/s1 ));
 AND2_X1 \V4/V1/A3/A1/M3/M2/_0_  (.A1(\V4/V1/A3/A1/M3/s1 ),
    .A2(\V4/V1/A3/A1/c2 ),
    .ZN(\V4/V1/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M3/M2/_1_  (.A(\V4/V1/A3/A1/M3/s1 ),
    .B(\V4/V1/A3/A1/c2 ),
    .Z(\V4/v1 [10]));
 OR2_X1 \V4/V1/A3/A1/M3/_0_  (.A1(\V4/V1/A3/A1/M3/c1 ),
    .A2(\V4/V1/A3/A1/M3/c2 ),
    .ZN(\V4/V1/A3/A1/c3 ));
 AND2_X1 \V4/V1/A3/A1/M4/M1/_0_  (.A1(\V4/V1/v4 [3]),
    .A2(\V4/V1/s2 [7]),
    .ZN(\V4/V1/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V1/A3/A1/M4/M1/_1_  (.A(\V4/V1/v4 [3]),
    .B(\V4/V1/s2 [7]),
    .Z(\V4/V1/A3/A1/M4/s1 ));
 AND2_X1 \V4/V1/A3/A1/M4/M2/_0_  (.A1(\V4/V1/A3/A1/M4/s1 ),
    .A2(\V4/V1/A3/A1/c3 ),
    .ZN(\V4/V1/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V1/A3/A1/M4/M2/_1_  (.A(\V4/V1/A3/A1/M4/s1 ),
    .B(\V4/V1/A3/A1/c3 ),
    .Z(\V4/v1 [11]));
 OR2_X1 \V4/V1/A3/A1/M4/_0_  (.A1(\V4/V1/A3/A1/M4/c1 ),
    .A2(\V4/V1/A3/A1/M4/c2 ),
    .ZN(\V4/V1/A3/c1 ));
 AND2_X1 \V4/V1/A3/A2/M1/M1/_0_  (.A1(\V4/V1/v4 [4]),
    .A2(\V4/V1/c3 ),
    .ZN(\V4/V1/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M1/M1/_1_  (.A(\V4/V1/v4 [4]),
    .B(\V4/V1/c3 ),
    .Z(\V4/V1/A3/A2/M1/s1 ));
 AND2_X1 \V4/V1/A3/A2/M1/M2/_0_  (.A1(\V4/V1/A3/A2/M1/s1 ),
    .A2(\V4/V1/A3/c1 ),
    .ZN(\V4/V1/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M1/M2/_1_  (.A(\V4/V1/A3/A2/M1/s1 ),
    .B(\V4/V1/A3/c1 ),
    .Z(\V4/v1 [12]));
 OR2_X1 \V4/V1/A3/A2/M1/_0_  (.A1(\V4/V1/A3/A2/M1/c1 ),
    .A2(\V4/V1/A3/A2/M1/c2 ),
    .ZN(\V4/V1/A3/A2/c1 ));
 AND2_X1 \V4/V1/A3/A2/M2/M1/_0_  (.A1(\V4/V1/v4 [5]),
    .A2(net1),
    .ZN(\V4/V1/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M2/M1/_1_  (.A(\V4/V1/v4 [5]),
    .B(net1),
    .Z(\V4/V1/A3/A2/M2/s1 ));
 AND2_X1 \V4/V1/A3/A2/M2/M2/_0_  (.A1(\V4/V1/A3/A2/M2/s1 ),
    .A2(\V4/V1/A3/A2/c1 ),
    .ZN(\V4/V1/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M2/M2/_1_  (.A(\V4/V1/A3/A2/M2/s1 ),
    .B(\V4/V1/A3/A2/c1 ),
    .Z(\V4/v1 [13]));
 OR2_X1 \V4/V1/A3/A2/M2/_0_  (.A1(\V4/V1/A3/A2/M2/c1 ),
    .A2(\V4/V1/A3/A2/M2/c2 ),
    .ZN(\V4/V1/A3/A2/c2 ));
 AND2_X1 \V4/V1/A3/A2/M3/M1/_0_  (.A1(\V4/V1/v4 [6]),
    .A2(net1),
    .ZN(\V4/V1/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M3/M1/_1_  (.A(\V4/V1/v4 [6]),
    .B(net1),
    .Z(\V4/V1/A3/A2/M3/s1 ));
 AND2_X1 \V4/V1/A3/A2/M3/M2/_0_  (.A1(\V4/V1/A3/A2/M3/s1 ),
    .A2(\V4/V1/A3/A2/c2 ),
    .ZN(\V4/V1/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M3/M2/_1_  (.A(\V4/V1/A3/A2/M3/s1 ),
    .B(\V4/V1/A3/A2/c2 ),
    .Z(\V4/v1 [14]));
 OR2_X1 \V4/V1/A3/A2/M3/_0_  (.A1(\V4/V1/A3/A2/M3/c1 ),
    .A2(\V4/V1/A3/A2/M3/c2 ),
    .ZN(\V4/V1/A3/A2/c3 ));
 AND2_X1 \V4/V1/A3/A2/M4/M1/_0_  (.A1(\V4/V1/v4 [7]),
    .A2(net1),
    .ZN(\V4/V1/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V1/A3/A2/M4/M1/_1_  (.A(\V4/V1/v4 [7]),
    .B(net1),
    .Z(\V4/V1/A3/A2/M4/s1 ));
 AND2_X1 \V4/V1/A3/A2/M4/M2/_0_  (.A1(\V4/V1/A3/A2/M4/s1 ),
    .A2(\V4/V1/A3/A2/c3 ),
    .ZN(\V4/V1/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V1/A3/A2/M4/M2/_1_  (.A(\V4/V1/A3/A2/M4/s1 ),
    .B(\V4/V1/A3/A2/c3 ),
    .Z(\V4/v1 [15]));
 OR2_X1 \V4/V1/A3/A2/M4/_0_  (.A1(\V4/V1/A3/A2/M4/c1 ),
    .A2(\V4/V1/A3/A2/M4/c2 ),
    .ZN(\V4/V1/overflow ));
 AND2_X1 \V4/V1/V1/A1/M1/M1/_0_  (.A1(\V4/V1/V1/v2 [0]),
    .A2(\V4/V1/V1/v3 [0]),
    .ZN(\V4/V1/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M1/M1/_1_  (.A(\V4/V1/V1/v2 [0]),
    .B(\V4/V1/V1/v3 [0]),
    .Z(\V4/V1/V1/A1/M1/s1 ));
 AND2_X1 \V4/V1/V1/A1/M1/M2/_0_  (.A1(\V4/V1/V1/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M1/M2/_1_  (.A(\V4/V1/V1/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/V1/V1/s1 [0]));
 OR2_X1 \V4/V1/V1/A1/M1/_0_  (.A1(\V4/V1/V1/A1/M1/c1 ),
    .A2(\V4/V1/V1/A1/M1/c2 ),
    .ZN(\V4/V1/V1/A1/c1 ));
 AND2_X1 \V4/V1/V1/A1/M2/M1/_0_  (.A1(\V4/V1/V1/v2 [1]),
    .A2(\V4/V1/V1/v3 [1]),
    .ZN(\V4/V1/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M2/M1/_1_  (.A(\V4/V1/V1/v2 [1]),
    .B(\V4/V1/V1/v3 [1]),
    .Z(\V4/V1/V1/A1/M2/s1 ));
 AND2_X1 \V4/V1/V1/A1/M2/M2/_0_  (.A1(\V4/V1/V1/A1/M2/s1 ),
    .A2(\V4/V1/V1/A1/c1 ),
    .ZN(\V4/V1/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M2/M2/_1_  (.A(\V4/V1/V1/A1/M2/s1 ),
    .B(\V4/V1/V1/A1/c1 ),
    .Z(\V4/V1/V1/s1 [1]));
 OR2_X1 \V4/V1/V1/A1/M2/_0_  (.A1(\V4/V1/V1/A1/M2/c1 ),
    .A2(\V4/V1/V1/A1/M2/c2 ),
    .ZN(\V4/V1/V1/A1/c2 ));
 AND2_X1 \V4/V1/V1/A1/M3/M1/_0_  (.A1(\V4/V1/V1/v2 [2]),
    .A2(\V4/V1/V1/v3 [2]),
    .ZN(\V4/V1/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M3/M1/_1_  (.A(\V4/V1/V1/v2 [2]),
    .B(\V4/V1/V1/v3 [2]),
    .Z(\V4/V1/V1/A1/M3/s1 ));
 AND2_X1 \V4/V1/V1/A1/M3/M2/_0_  (.A1(\V4/V1/V1/A1/M3/s1 ),
    .A2(\V4/V1/V1/A1/c2 ),
    .ZN(\V4/V1/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M3/M2/_1_  (.A(\V4/V1/V1/A1/M3/s1 ),
    .B(\V4/V1/V1/A1/c2 ),
    .Z(\V4/V1/V1/s1 [2]));
 OR2_X1 \V4/V1/V1/A1/M3/_0_  (.A1(\V4/V1/V1/A1/M3/c1 ),
    .A2(\V4/V1/V1/A1/M3/c2 ),
    .ZN(\V4/V1/V1/A1/c3 ));
 AND2_X1 \V4/V1/V1/A1/M4/M1/_0_  (.A1(\V4/V1/V1/v2 [3]),
    .A2(\V4/V1/V1/v3 [3]),
    .ZN(\V4/V1/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A1/M4/M1/_1_  (.A(\V4/V1/V1/v2 [3]),
    .B(\V4/V1/V1/v3 [3]),
    .Z(\V4/V1/V1/A1/M4/s1 ));
 AND2_X1 \V4/V1/V1/A1/M4/M2/_0_  (.A1(\V4/V1/V1/A1/M4/s1 ),
    .A2(\V4/V1/V1/A1/c3 ),
    .ZN(\V4/V1/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A1/M4/M2/_1_  (.A(\V4/V1/V1/A1/M4/s1 ),
    .B(\V4/V1/V1/A1/c3 ),
    .Z(\V4/V1/V1/s1 [3]));
 OR2_X1 \V4/V1/V1/A1/M4/_0_  (.A1(\V4/V1/V1/A1/M4/c1 ),
    .A2(\V4/V1/V1/A1/M4/c2 ),
    .ZN(\V4/V1/V1/c1 ));
 AND2_X1 \V4/V1/V1/A2/M1/M1/_0_  (.A1(\V4/V1/V1/s1 [0]),
    .A2(\V4/V1/V1/v1 [2]),
    .ZN(\V4/V1/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M1/M1/_1_  (.A(\V4/V1/V1/s1 [0]),
    .B(\V4/V1/V1/v1 [2]),
    .Z(\V4/V1/V1/A2/M1/s1 ));
 AND2_X1 \V4/V1/V1/A2/M1/M2/_0_  (.A1(\V4/V1/V1/A2/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M1/M2/_1_  (.A(\V4/V1/V1/A2/M1/s1 ),
    .B(net9),
    .Z(v4[2]));
 OR2_X1 \V4/V1/V1/A2/M1/_0_  (.A1(\V4/V1/V1/A2/M1/c1 ),
    .A2(\V4/V1/V1/A2/M1/c2 ),
    .ZN(\V4/V1/V1/A2/c1 ));
 AND2_X1 \V4/V1/V1/A2/M2/M1/_0_  (.A1(\V4/V1/V1/s1 [1]),
    .A2(\V4/V1/V1/v1 [3]),
    .ZN(\V4/V1/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M2/M1/_1_  (.A(\V4/V1/V1/s1 [1]),
    .B(\V4/V1/V1/v1 [3]),
    .Z(\V4/V1/V1/A2/M2/s1 ));
 AND2_X1 \V4/V1/V1/A2/M2/M2/_0_  (.A1(\V4/V1/V1/A2/M2/s1 ),
    .A2(\V4/V1/V1/A2/c1 ),
    .ZN(\V4/V1/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M2/M2/_1_  (.A(\V4/V1/V1/A2/M2/s1 ),
    .B(\V4/V1/V1/A2/c1 ),
    .Z(v4[3]));
 OR2_X1 \V4/V1/V1/A2/M2/_0_  (.A1(\V4/V1/V1/A2/M2/c1 ),
    .A2(\V4/V1/V1/A2/M2/c2 ),
    .ZN(\V4/V1/V1/A2/c2 ));
 AND2_X1 \V4/V1/V1/A2/M3/M1/_0_  (.A1(\V4/V1/V1/s1 [2]),
    .A2(net9),
    .ZN(\V4/V1/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M3/M1/_1_  (.A(\V4/V1/V1/s1 [2]),
    .B(net9),
    .Z(\V4/V1/V1/A2/M3/s1 ));
 AND2_X1 \V4/V1/V1/A2/M3/M2/_0_  (.A1(\V4/V1/V1/A2/M3/s1 ),
    .A2(\V4/V1/V1/A2/c2 ),
    .ZN(\V4/V1/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M3/M2/_1_  (.A(\V4/V1/V1/A2/M3/s1 ),
    .B(\V4/V1/V1/A2/c2 ),
    .Z(\V4/V1/V1/s2 [2]));
 OR2_X1 \V4/V1/V1/A2/M3/_0_  (.A1(\V4/V1/V1/A2/M3/c1 ),
    .A2(\V4/V1/V1/A2/M3/c2 ),
    .ZN(\V4/V1/V1/A2/c3 ));
 AND2_X1 \V4/V1/V1/A2/M4/M1/_0_  (.A1(\V4/V1/V1/s1 [3]),
    .A2(net9),
    .ZN(\V4/V1/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A2/M4/M1/_1_  (.A(\V4/V1/V1/s1 [3]),
    .B(net9),
    .Z(\V4/V1/V1/A2/M4/s1 ));
 AND2_X1 \V4/V1/V1/A2/M4/M2/_0_  (.A1(\V4/V1/V1/A2/M4/s1 ),
    .A2(\V4/V1/V1/A2/c3 ),
    .ZN(\V4/V1/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A2/M4/M2/_1_  (.A(\V4/V1/V1/A2/M4/s1 ),
    .B(\V4/V1/V1/A2/c3 ),
    .Z(\V4/V1/V1/s2 [3]));
 OR2_X1 \V4/V1/V1/A2/M4/_0_  (.A1(\V4/V1/V1/A2/M4/c1 ),
    .A2(\V4/V1/V1/A2/M4/c2 ),
    .ZN(\V4/V1/V1/c2 ));
 AND2_X1 \V4/V1/V1/A3/M1/M1/_0_  (.A1(\V4/V1/V1/v4 [0]),
    .A2(\V4/V1/V1/s2 [2]),
    .ZN(\V4/V1/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M1/M1/_1_  (.A(\V4/V1/V1/v4 [0]),
    .B(\V4/V1/V1/s2 [2]),
    .Z(\V4/V1/V1/A3/M1/s1 ));
 AND2_X1 \V4/V1/V1/A3/M1/M2/_0_  (.A1(\V4/V1/V1/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V1/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M1/M2/_1_  (.A(\V4/V1/V1/A3/M1/s1 ),
    .B(net9),
    .Z(\V4/V1/v1 [4]));
 OR2_X1 \V4/V1/V1/A3/M1/_0_  (.A1(\V4/V1/V1/A3/M1/c1 ),
    .A2(\V4/V1/V1/A3/M1/c2 ),
    .ZN(\V4/V1/V1/A3/c1 ));
 AND2_X1 \V4/V1/V1/A3/M2/M1/_0_  (.A1(\V4/V1/V1/v4 [1]),
    .A2(\V4/V1/V1/s2 [3]),
    .ZN(\V4/V1/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M2/M1/_1_  (.A(\V4/V1/V1/v4 [1]),
    .B(\V4/V1/V1/s2 [3]),
    .Z(\V4/V1/V1/A3/M2/s1 ));
 AND2_X1 \V4/V1/V1/A3/M2/M2/_0_  (.A1(\V4/V1/V1/A3/M2/s1 ),
    .A2(\V4/V1/V1/A3/c1 ),
    .ZN(\V4/V1/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M2/M2/_1_  (.A(\V4/V1/V1/A3/M2/s1 ),
    .B(\V4/V1/V1/A3/c1 ),
    .Z(\V4/V1/v1 [5]));
 OR2_X1 \V4/V1/V1/A3/M2/_0_  (.A1(\V4/V1/V1/A3/M2/c1 ),
    .A2(\V4/V1/V1/A3/M2/c2 ),
    .ZN(\V4/V1/V1/A3/c2 ));
 AND2_X1 \V4/V1/V1/A3/M3/M1/_0_  (.A1(\V4/V1/V1/v4 [2]),
    .A2(\V4/V1/V1/c3 ),
    .ZN(\V4/V1/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M3/M1/_1_  (.A(\V4/V1/V1/v4 [2]),
    .B(\V4/V1/V1/c3 ),
    .Z(\V4/V1/V1/A3/M3/s1 ));
 AND2_X1 \V4/V1/V1/A3/M3/M2/_0_  (.A1(\V4/V1/V1/A3/M3/s1 ),
    .A2(\V4/V1/V1/A3/c2 ),
    .ZN(\V4/V1/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M3/M2/_1_  (.A(\V4/V1/V1/A3/M3/s1 ),
    .B(\V4/V1/V1/A3/c2 ),
    .Z(\V4/V1/v1 [6]));
 OR2_X1 \V4/V1/V1/A3/M3/_0_  (.A1(\V4/V1/V1/A3/M3/c1 ),
    .A2(\V4/V1/V1/A3/M3/c2 ),
    .ZN(\V4/V1/V1/A3/c3 ));
 AND2_X1 \V4/V1/V1/A3/M4/M1/_0_  (.A1(\V4/V1/V1/v4 [3]),
    .A2(net10),
    .ZN(\V4/V1/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V1/A3/M4/M1/_1_  (.A(\V4/V1/V1/v4 [3]),
    .B(net10),
    .Z(\V4/V1/V1/A3/M4/s1 ));
 AND2_X1 \V4/V1/V1/A3/M4/M2/_0_  (.A1(\V4/V1/V1/A3/M4/s1 ),
    .A2(\V4/V1/V1/A3/c3 ),
    .ZN(\V4/V1/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V1/A3/M4/M2/_1_  (.A(\V4/V1/V1/A3/M4/s1 ),
    .B(\V4/V1/V1/A3/c3 ),
    .Z(\V4/V1/v1 [7]));
 OR2_X1 \V4/V1/V1/A3/M4/_0_  (.A1(\V4/V1/V1/A3/M4/c1 ),
    .A2(\V4/V1/V1/A3/M4/c2 ),
    .ZN(\V4/V1/V1/overflow ));
 AND2_X1 \V4/V1/V1/V1/HA1/_0_  (.A1(\V4/V1/V1/V1/w2 ),
    .A2(\V4/V1/V1/V1/w1 ),
    .ZN(\V4/V1/V1/V1/w4 ));
 XOR2_X2 \V4/V1/V1/V1/HA1/_1_  (.A(\V4/V1/V1/V1/w2 ),
    .B(\V4/V1/V1/V1/w1 ),
    .Z(v4[1]));
 AND2_X1 \V4/V1/V1/V1/HA2/_0_  (.A1(\V4/V1/V1/V1/w4 ),
    .A2(\V4/V1/V1/V1/w3 ),
    .ZN(\V4/V1/V1/v1 [3]));
 XOR2_X2 \V4/V1/V1/V1/HA2/_1_  (.A(\V4/V1/V1/V1/w4 ),
    .B(\V4/V1/V1/V1/w3 ),
    .Z(\V4/V1/V1/v1 [2]));
 AND2_X1 \V4/V1/V1/V1/_0_  (.A1(net41),
    .A2(net22),
    .ZN(v4[0]));
 AND2_X1 \V4/V1/V1/V1/_1_  (.A1(net41),
    .A2(net21),
    .ZN(\V4/V1/V1/V1/w1 ));
 AND2_X1 \V4/V1/V1/V1/_2_  (.A1(net22),
    .A2(net40),
    .ZN(\V4/V1/V1/V1/w2 ));
 AND2_X1 \V4/V1/V1/V1/_3_  (.A1(net21),
    .A2(net40),
    .ZN(\V4/V1/V1/V1/w3 ));
 AND2_X1 \V4/V1/V1/V2/HA1/_0_  (.A1(\V4/V1/V1/V2/w2 ),
    .A2(\V4/V1/V1/V2/w1 ),
    .ZN(\V4/V1/V1/V2/w4 ));
 XOR2_X2 \V4/V1/V1/V2/HA1/_1_  (.A(\V4/V1/V1/V2/w2 ),
    .B(\V4/V1/V1/V2/w1 ),
    .Z(\V4/V1/V1/v2 [1]));
 AND2_X1 \V4/V1/V1/V2/HA2/_0_  (.A1(\V4/V1/V1/V2/w4 ),
    .A2(\V4/V1/V1/V2/w3 ),
    .ZN(\V4/V1/V1/v2 [3]));
 XOR2_X2 \V4/V1/V1/V2/HA2/_1_  (.A(\V4/V1/V1/V2/w4 ),
    .B(\V4/V1/V1/V2/w3 ),
    .Z(\V4/V1/V1/v2 [2]));
 AND2_X1 \V4/V1/V1/V2/_0_  (.A1(net39),
    .A2(net22),
    .ZN(\V4/V1/V1/v2 [0]));
 AND2_X1 \V4/V1/V1/V2/_1_  (.A1(net39),
    .A2(net21),
    .ZN(\V4/V1/V1/V2/w1 ));
 AND2_X1 \V4/V1/V1/V2/_2_  (.A1(net22),
    .A2(net38),
    .ZN(\V4/V1/V1/V2/w2 ));
 AND2_X1 \V4/V1/V1/V2/_3_  (.A1(net21),
    .A2(net38),
    .ZN(\V4/V1/V1/V2/w3 ));
 AND2_X1 \V4/V1/V1/V3/HA1/_0_  (.A1(\V4/V1/V1/V3/w2 ),
    .A2(\V4/V1/V1/V3/w1 ),
    .ZN(\V4/V1/V1/V3/w4 ));
 XOR2_X2 \V4/V1/V1/V3/HA1/_1_  (.A(\V4/V1/V1/V3/w2 ),
    .B(\V4/V1/V1/V3/w1 ),
    .Z(\V4/V1/V1/v3 [1]));
 AND2_X1 \V4/V1/V1/V3/HA2/_0_  (.A1(\V4/V1/V1/V3/w4 ),
    .A2(\V4/V1/V1/V3/w3 ),
    .ZN(\V4/V1/V1/v3 [3]));
 XOR2_X2 \V4/V1/V1/V3/HA2/_1_  (.A(\V4/V1/V1/V3/w4 ),
    .B(\V4/V1/V1/V3/w3 ),
    .Z(\V4/V1/V1/v3 [2]));
 AND2_X1 \V4/V1/V1/V3/_0_  (.A1(net41),
    .A2(net20),
    .ZN(\V4/V1/V1/v3 [0]));
 AND2_X1 \V4/V1/V1/V3/_1_  (.A1(net41),
    .A2(net19),
    .ZN(\V4/V1/V1/V3/w1 ));
 AND2_X1 \V4/V1/V1/V3/_2_  (.A1(net20),
    .A2(net40),
    .ZN(\V4/V1/V1/V3/w2 ));
 AND2_X1 \V4/V1/V1/V3/_3_  (.A1(net19),
    .A2(net40),
    .ZN(\V4/V1/V1/V3/w3 ));
 AND2_X1 \V4/V1/V1/V4/HA1/_0_  (.A1(\V4/V1/V1/V4/w2 ),
    .A2(\V4/V1/V1/V4/w1 ),
    .ZN(\V4/V1/V1/V4/w4 ));
 XOR2_X2 \V4/V1/V1/V4/HA1/_1_  (.A(\V4/V1/V1/V4/w2 ),
    .B(\V4/V1/V1/V4/w1 ),
    .Z(\V4/V1/V1/v4 [1]));
 AND2_X1 \V4/V1/V1/V4/HA2/_0_  (.A1(\V4/V1/V1/V4/w4 ),
    .A2(\V4/V1/V1/V4/w3 ),
    .ZN(\V4/V1/V1/v4 [3]));
 XOR2_X2 \V4/V1/V1/V4/HA2/_1_  (.A(\V4/V1/V1/V4/w4 ),
    .B(\V4/V1/V1/V4/w3 ),
    .Z(\V4/V1/V1/v4 [2]));
 AND2_X1 \V4/V1/V1/V4/_0_  (.A1(net39),
    .A2(net20),
    .ZN(\V4/V1/V1/v4 [0]));
 AND2_X1 \V4/V1/V1/V4/_1_  (.A1(net39),
    .A2(net19),
    .ZN(\V4/V1/V1/V4/w1 ));
 AND2_X1 \V4/V1/V1/V4/_2_  (.A1(net20),
    .A2(net38),
    .ZN(\V4/V1/V1/V4/w2 ));
 AND2_X1 \V4/V1/V1/V4/_3_  (.A1(net19),
    .A2(net38),
    .ZN(\V4/V1/V1/V4/w3 ));
 OR2_X1 \V4/V1/V1/_0_  (.A1(\V4/V1/V1/c1 ),
    .A2(\V4/V1/V1/c2 ),
    .ZN(\V4/V1/V1/c3 ));
 AND2_X1 \V4/V1/V2/A1/M1/M1/_0_  (.A1(\V4/V1/V2/v2 [0]),
    .A2(\V4/V1/V2/v3 [0]),
    .ZN(\V4/V1/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M1/M1/_1_  (.A(\V4/V1/V2/v2 [0]),
    .B(\V4/V1/V2/v3 [0]),
    .Z(\V4/V1/V2/A1/M1/s1 ));
 AND2_X1 \V4/V1/V2/A1/M1/M2/_0_  (.A1(\V4/V1/V2/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V1/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M1/M2/_1_  (.A(\V4/V1/V2/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V1/V2/s1 [0]));
 OR2_X1 \V4/V1/V2/A1/M1/_0_  (.A1(\V4/V1/V2/A1/M1/c1 ),
    .A2(\V4/V1/V2/A1/M1/c2 ),
    .ZN(\V4/V1/V2/A1/c1 ));
 AND2_X1 \V4/V1/V2/A1/M2/M1/_0_  (.A1(\V4/V1/V2/v2 [1]),
    .A2(\V4/V1/V2/v3 [1]),
    .ZN(\V4/V1/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M2/M1/_1_  (.A(\V4/V1/V2/v2 [1]),
    .B(\V4/V1/V2/v3 [1]),
    .Z(\V4/V1/V2/A1/M2/s1 ));
 AND2_X1 \V4/V1/V2/A1/M2/M2/_0_  (.A1(\V4/V1/V2/A1/M2/s1 ),
    .A2(\V4/V1/V2/A1/c1 ),
    .ZN(\V4/V1/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M2/M2/_1_  (.A(\V4/V1/V2/A1/M2/s1 ),
    .B(\V4/V1/V2/A1/c1 ),
    .Z(\V4/V1/V2/s1 [1]));
 OR2_X1 \V4/V1/V2/A1/M2/_0_  (.A1(\V4/V1/V2/A1/M2/c1 ),
    .A2(\V4/V1/V2/A1/M2/c2 ),
    .ZN(\V4/V1/V2/A1/c2 ));
 AND2_X1 \V4/V1/V2/A1/M3/M1/_0_  (.A1(\V4/V1/V2/v2 [2]),
    .A2(\V4/V1/V2/v3 [2]),
    .ZN(\V4/V1/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M3/M1/_1_  (.A(\V4/V1/V2/v2 [2]),
    .B(\V4/V1/V2/v3 [2]),
    .Z(\V4/V1/V2/A1/M3/s1 ));
 AND2_X1 \V4/V1/V2/A1/M3/M2/_0_  (.A1(\V4/V1/V2/A1/M3/s1 ),
    .A2(\V4/V1/V2/A1/c2 ),
    .ZN(\V4/V1/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M3/M2/_1_  (.A(\V4/V1/V2/A1/M3/s1 ),
    .B(\V4/V1/V2/A1/c2 ),
    .Z(\V4/V1/V2/s1 [2]));
 OR2_X1 \V4/V1/V2/A1/M3/_0_  (.A1(\V4/V1/V2/A1/M3/c1 ),
    .A2(\V4/V1/V2/A1/M3/c2 ),
    .ZN(\V4/V1/V2/A1/c3 ));
 AND2_X1 \V4/V1/V2/A1/M4/M1/_0_  (.A1(\V4/V1/V2/v2 [3]),
    .A2(\V4/V1/V2/v3 [3]),
    .ZN(\V4/V1/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A1/M4/M1/_1_  (.A(\V4/V1/V2/v2 [3]),
    .B(\V4/V1/V2/v3 [3]),
    .Z(\V4/V1/V2/A1/M4/s1 ));
 AND2_X1 \V4/V1/V2/A1/M4/M2/_0_  (.A1(\V4/V1/V2/A1/M4/s1 ),
    .A2(\V4/V1/V2/A1/c3 ),
    .ZN(\V4/V1/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A1/M4/M2/_1_  (.A(\V4/V1/V2/A1/M4/s1 ),
    .B(\V4/V1/V2/A1/c3 ),
    .Z(\V4/V1/V2/s1 [3]));
 OR2_X1 \V4/V1/V2/A1/M4/_0_  (.A1(\V4/V1/V2/A1/M4/c1 ),
    .A2(\V4/V1/V2/A1/M4/c2 ),
    .ZN(\V4/V1/V2/c1 ));
 AND2_X1 \V4/V1/V2/A2/M1/M1/_0_  (.A1(\V4/V1/V2/s1 [0]),
    .A2(\V4/V1/V2/v1 [2]),
    .ZN(\V4/V1/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M1/M1/_1_  (.A(\V4/V1/V2/s1 [0]),
    .B(\V4/V1/V2/v1 [2]),
    .Z(\V4/V1/V2/A2/M1/s1 ));
 AND2_X1 \V4/V1/V2/A2/M1/M2/_0_  (.A1(\V4/V1/V2/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V1/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M1/M2/_1_  (.A(\V4/V1/V2/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/v2 [2]));
 OR2_X1 \V4/V1/V2/A2/M1/_0_  (.A1(\V4/V1/V2/A2/M1/c1 ),
    .A2(\V4/V1/V2/A2/M1/c2 ),
    .ZN(\V4/V1/V2/A2/c1 ));
 AND2_X1 \V4/V1/V2/A2/M2/M1/_0_  (.A1(\V4/V1/V2/s1 [1]),
    .A2(\V4/V1/V2/v1 [3]),
    .ZN(\V4/V1/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M2/M1/_1_  (.A(\V4/V1/V2/s1 [1]),
    .B(\V4/V1/V2/v1 [3]),
    .Z(\V4/V1/V2/A2/M2/s1 ));
 AND2_X1 \V4/V1/V2/A2/M2/M2/_0_  (.A1(\V4/V1/V2/A2/M2/s1 ),
    .A2(\V4/V1/V2/A2/c1 ),
    .ZN(\V4/V1/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M2/M2/_1_  (.A(\V4/V1/V2/A2/M2/s1 ),
    .B(\V4/V1/V2/A2/c1 ),
    .Z(\V4/V1/v2 [3]));
 OR2_X1 \V4/V1/V2/A2/M2/_0_  (.A1(\V4/V1/V2/A2/M2/c1 ),
    .A2(\V4/V1/V2/A2/M2/c2 ),
    .ZN(\V4/V1/V2/A2/c2 ));
 AND2_X1 \V4/V1/V2/A2/M3/M1/_0_  (.A1(\V4/V1/V2/s1 [2]),
    .A2(net1),
    .ZN(\V4/V1/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M3/M1/_1_  (.A(\V4/V1/V2/s1 [2]),
    .B(net1),
    .Z(\V4/V1/V2/A2/M3/s1 ));
 AND2_X1 \V4/V1/V2/A2/M3/M2/_0_  (.A1(\V4/V1/V2/A2/M3/s1 ),
    .A2(\V4/V1/V2/A2/c2 ),
    .ZN(\V4/V1/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M3/M2/_1_  (.A(\V4/V1/V2/A2/M3/s1 ),
    .B(\V4/V1/V2/A2/c2 ),
    .Z(\V4/V1/V2/s2 [2]));
 OR2_X1 \V4/V1/V2/A2/M3/_0_  (.A1(\V4/V1/V2/A2/M3/c1 ),
    .A2(\V4/V1/V2/A2/M3/c2 ),
    .ZN(\V4/V1/V2/A2/c3 ));
 AND2_X1 \V4/V1/V2/A2/M4/M1/_0_  (.A1(\V4/V1/V2/s1 [3]),
    .A2(net1),
    .ZN(\V4/V1/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A2/M4/M1/_1_  (.A(\V4/V1/V2/s1 [3]),
    .B(net1),
    .Z(\V4/V1/V2/A2/M4/s1 ));
 AND2_X1 \V4/V1/V2/A2/M4/M2/_0_  (.A1(\V4/V1/V2/A2/M4/s1 ),
    .A2(\V4/V1/V2/A2/c3 ),
    .ZN(\V4/V1/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A2/M4/M2/_1_  (.A(\V4/V1/V2/A2/M4/s1 ),
    .B(\V4/V1/V2/A2/c3 ),
    .Z(\V4/V1/V2/s2 [3]));
 OR2_X1 \V4/V1/V2/A2/M4/_0_  (.A1(\V4/V1/V2/A2/M4/c1 ),
    .A2(\V4/V1/V2/A2/M4/c2 ),
    .ZN(\V4/V1/V2/c2 ));
 AND2_X1 \V4/V1/V2/A3/M1/M1/_0_  (.A1(\V4/V1/V2/v4 [0]),
    .A2(\V4/V1/V2/s2 [2]),
    .ZN(\V4/V1/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M1/M1/_1_  (.A(\V4/V1/V2/v4 [0]),
    .B(\V4/V1/V2/s2 [2]),
    .Z(\V4/V1/V2/A3/M1/s1 ));
 AND2_X1 \V4/V1/V2/A3/M1/M2/_0_  (.A1(\V4/V1/V2/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V1/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M1/M2/_1_  (.A(\V4/V1/V2/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/v2 [4]));
 OR2_X1 \V4/V1/V2/A3/M1/_0_  (.A1(\V4/V1/V2/A3/M1/c1 ),
    .A2(\V4/V1/V2/A3/M1/c2 ),
    .ZN(\V4/V1/V2/A3/c1 ));
 AND2_X1 \V4/V1/V2/A3/M2/M1/_0_  (.A1(\V4/V1/V2/v4 [1]),
    .A2(\V4/V1/V2/s2 [3]),
    .ZN(\V4/V1/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M2/M1/_1_  (.A(\V4/V1/V2/v4 [1]),
    .B(\V4/V1/V2/s2 [3]),
    .Z(\V4/V1/V2/A3/M2/s1 ));
 AND2_X1 \V4/V1/V2/A3/M2/M2/_0_  (.A1(\V4/V1/V2/A3/M2/s1 ),
    .A2(\V4/V1/V2/A3/c1 ),
    .ZN(\V4/V1/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M2/M2/_1_  (.A(\V4/V1/V2/A3/M2/s1 ),
    .B(\V4/V1/V2/A3/c1 ),
    .Z(\V4/V1/v2 [5]));
 OR2_X1 \V4/V1/V2/A3/M2/_0_  (.A1(\V4/V1/V2/A3/M2/c1 ),
    .A2(\V4/V1/V2/A3/M2/c2 ),
    .ZN(\V4/V1/V2/A3/c2 ));
 AND2_X1 \V4/V1/V2/A3/M3/M1/_0_  (.A1(\V4/V1/V2/v4 [2]),
    .A2(\V4/V1/V2/c3 ),
    .ZN(\V4/V1/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M3/M1/_1_  (.A(\V4/V1/V2/v4 [2]),
    .B(\V4/V1/V2/c3 ),
    .Z(\V4/V1/V2/A3/M3/s1 ));
 AND2_X1 \V4/V1/V2/A3/M3/M2/_0_  (.A1(\V4/V1/V2/A3/M3/s1 ),
    .A2(\V4/V1/V2/A3/c2 ),
    .ZN(\V4/V1/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M3/M2/_1_  (.A(\V4/V1/V2/A3/M3/s1 ),
    .B(\V4/V1/V2/A3/c2 ),
    .Z(\V4/V1/v2 [6]));
 OR2_X1 \V4/V1/V2/A3/M3/_0_  (.A1(\V4/V1/V2/A3/M3/c1 ),
    .A2(\V4/V1/V2/A3/M3/c2 ),
    .ZN(\V4/V1/V2/A3/c3 ));
 AND2_X1 \V4/V1/V2/A3/M4/M1/_0_  (.A1(\V4/V1/V2/v4 [3]),
    .A2(net1),
    .ZN(\V4/V1/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V2/A3/M4/M1/_1_  (.A(\V4/V1/V2/v4 [3]),
    .B(net1),
    .Z(\V4/V1/V2/A3/M4/s1 ));
 AND2_X1 \V4/V1/V2/A3/M4/M2/_0_  (.A1(\V4/V1/V2/A3/M4/s1 ),
    .A2(\V4/V1/V2/A3/c3 ),
    .ZN(\V4/V1/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V2/A3/M4/M2/_1_  (.A(\V4/V1/V2/A3/M4/s1 ),
    .B(\V4/V1/V2/A3/c3 ),
    .Z(\V4/V1/v2 [7]));
 OR2_X1 \V4/V1/V2/A3/M4/_0_  (.A1(\V4/V1/V2/A3/M4/c1 ),
    .A2(\V4/V1/V2/A3/M4/c2 ),
    .ZN(\V4/V1/V2/overflow ));
 AND2_X1 \V4/V1/V2/V1/HA1/_0_  (.A1(\V4/V1/V2/V1/w2 ),
    .A2(\V4/V1/V2/V1/w1 ),
    .ZN(\V4/V1/V2/V1/w4 ));
 XOR2_X2 \V4/V1/V2/V1/HA1/_1_  (.A(\V4/V1/V2/V1/w2 ),
    .B(\V4/V1/V2/V1/w1 ),
    .Z(\V4/V1/v2 [1]));
 AND2_X1 \V4/V1/V2/V1/HA2/_0_  (.A1(\V4/V1/V2/V1/w4 ),
    .A2(\V4/V1/V2/V1/w3 ),
    .ZN(\V4/V1/V2/v1 [3]));
 XOR2_X2 \V4/V1/V2/V1/HA2/_1_  (.A(\V4/V1/V2/V1/w4 ),
    .B(\V4/V1/V2/V1/w3 ),
    .Z(\V4/V1/V2/v1 [2]));
 AND2_X1 \V4/V1/V2/V1/_0_  (.A1(net37),
    .A2(net22),
    .ZN(\V4/V1/v2 [0]));
 AND2_X1 \V4/V1/V2/V1/_1_  (.A1(net37),
    .A2(net21),
    .ZN(\V4/V1/V2/V1/w1 ));
 AND2_X1 \V4/V1/V2/V1/_2_  (.A1(net22),
    .A2(net36),
    .ZN(\V4/V1/V2/V1/w2 ));
 AND2_X1 \V4/V1/V2/V1/_3_  (.A1(net21),
    .A2(net36),
    .ZN(\V4/V1/V2/V1/w3 ));
 AND2_X1 \V4/V1/V2/V2/HA1/_0_  (.A1(\V4/V1/V2/V2/w2 ),
    .A2(\V4/V1/V2/V2/w1 ),
    .ZN(\V4/V1/V2/V2/w4 ));
 XOR2_X2 \V4/V1/V2/V2/HA1/_1_  (.A(\V4/V1/V2/V2/w2 ),
    .B(\V4/V1/V2/V2/w1 ),
    .Z(\V4/V1/V2/v2 [1]));
 AND2_X1 \V4/V1/V2/V2/HA2/_0_  (.A1(\V4/V1/V2/V2/w4 ),
    .A2(\V4/V1/V2/V2/w3 ),
    .ZN(\V4/V1/V2/v2 [3]));
 XOR2_X2 \V4/V1/V2/V2/HA2/_1_  (.A(\V4/V1/V2/V2/w4 ),
    .B(\V4/V1/V2/V2/w3 ),
    .Z(\V4/V1/V2/v2 [2]));
 AND2_X1 \V4/V1/V2/V2/_0_  (.A1(net35),
    .A2(net22),
    .ZN(\V4/V1/V2/v2 [0]));
 AND2_X1 \V4/V1/V2/V2/_1_  (.A1(net35),
    .A2(net21),
    .ZN(\V4/V1/V2/V2/w1 ));
 AND2_X1 \V4/V1/V2/V2/_2_  (.A1(net22),
    .A2(net34),
    .ZN(\V4/V1/V2/V2/w2 ));
 AND2_X1 \V4/V1/V2/V2/_3_  (.A1(net21),
    .A2(net34),
    .ZN(\V4/V1/V2/V2/w3 ));
 AND2_X1 \V4/V1/V2/V3/HA1/_0_  (.A1(\V4/V1/V2/V3/w2 ),
    .A2(\V4/V1/V2/V3/w1 ),
    .ZN(\V4/V1/V2/V3/w4 ));
 XOR2_X2 \V4/V1/V2/V3/HA1/_1_  (.A(\V4/V1/V2/V3/w2 ),
    .B(\V4/V1/V2/V3/w1 ),
    .Z(\V4/V1/V2/v3 [1]));
 AND2_X1 \V4/V1/V2/V3/HA2/_0_  (.A1(\V4/V1/V2/V3/w4 ),
    .A2(\V4/V1/V2/V3/w3 ),
    .ZN(\V4/V1/V2/v3 [3]));
 XOR2_X2 \V4/V1/V2/V3/HA2/_1_  (.A(\V4/V1/V2/V3/w4 ),
    .B(\V4/V1/V2/V3/w3 ),
    .Z(\V4/V1/V2/v3 [2]));
 AND2_X1 \V4/V1/V2/V3/_0_  (.A1(net37),
    .A2(net20),
    .ZN(\V4/V1/V2/v3 [0]));
 AND2_X1 \V4/V1/V2/V3/_1_  (.A1(net37),
    .A2(net19),
    .ZN(\V4/V1/V2/V3/w1 ));
 AND2_X1 \V4/V1/V2/V3/_2_  (.A1(net20),
    .A2(net36),
    .ZN(\V4/V1/V2/V3/w2 ));
 AND2_X1 \V4/V1/V2/V3/_3_  (.A1(B[19]),
    .A2(net36),
    .ZN(\V4/V1/V2/V3/w3 ));
 AND2_X1 \V4/V1/V2/V4/HA1/_0_  (.A1(\V4/V1/V2/V4/w2 ),
    .A2(\V4/V1/V2/V4/w1 ),
    .ZN(\V4/V1/V2/V4/w4 ));
 XOR2_X2 \V4/V1/V2/V4/HA1/_1_  (.A(\V4/V1/V2/V4/w2 ),
    .B(\V4/V1/V2/V4/w1 ),
    .Z(\V4/V1/V2/v4 [1]));
 AND2_X1 \V4/V1/V2/V4/HA2/_0_  (.A1(\V4/V1/V2/V4/w4 ),
    .A2(\V4/V1/V2/V4/w3 ),
    .ZN(\V4/V1/V2/v4 [3]));
 XOR2_X2 \V4/V1/V2/V4/HA2/_1_  (.A(\V4/V1/V2/V4/w4 ),
    .B(\V4/V1/V2/V4/w3 ),
    .Z(\V4/V1/V2/v4 [2]));
 AND2_X1 \V4/V1/V2/V4/_0_  (.A1(net35),
    .A2(net20),
    .ZN(\V4/V1/V2/v4 [0]));
 AND2_X1 \V4/V1/V2/V4/_1_  (.A1(net35),
    .A2(B[19]),
    .ZN(\V4/V1/V2/V4/w1 ));
 AND2_X1 \V4/V1/V2/V4/_2_  (.A1(B[18]),
    .A2(net34),
    .ZN(\V4/V1/V2/V4/w2 ));
 AND2_X1 \V4/V1/V2/V4/_3_  (.A1(B[19]),
    .A2(net34),
    .ZN(\V4/V1/V2/V4/w3 ));
 OR2_X1 \V4/V1/V2/_0_  (.A1(\V4/V1/V2/c1 ),
    .A2(\V4/V1/V2/c2 ),
    .ZN(\V4/V1/V2/c3 ));
 AND2_X1 \V4/V1/V3/A1/M1/M1/_0_  (.A1(\V4/V1/V3/v2 [0]),
    .A2(\V4/V1/V3/v3 [0]),
    .ZN(\V4/V1/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M1/M1/_1_  (.A(\V4/V1/V3/v2 [0]),
    .B(\V4/V1/V3/v3 [0]),
    .Z(\V4/V1/V3/A1/M1/s1 ));
 AND2_X1 \V4/V1/V3/A1/M1/M2/_0_  (.A1(\V4/V1/V3/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V1/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M1/M2/_1_  (.A(\V4/V1/V3/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/V3/s1 [0]));
 OR2_X1 \V4/V1/V3/A1/M1/_0_  (.A1(\V4/V1/V3/A1/M1/c1 ),
    .A2(\V4/V1/V3/A1/M1/c2 ),
    .ZN(\V4/V1/V3/A1/c1 ));
 AND2_X1 \V4/V1/V3/A1/M2/M1/_0_  (.A1(\V4/V1/V3/v2 [1]),
    .A2(\V4/V1/V3/v3 [1]),
    .ZN(\V4/V1/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M2/M1/_1_  (.A(\V4/V1/V3/v2 [1]),
    .B(\V4/V1/V3/v3 [1]),
    .Z(\V4/V1/V3/A1/M2/s1 ));
 AND2_X1 \V4/V1/V3/A1/M2/M2/_0_  (.A1(\V4/V1/V3/A1/M2/s1 ),
    .A2(\V4/V1/V3/A1/c1 ),
    .ZN(\V4/V1/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M2/M2/_1_  (.A(\V4/V1/V3/A1/M2/s1 ),
    .B(\V4/V1/V3/A1/c1 ),
    .Z(\V4/V1/V3/s1 [1]));
 OR2_X1 \V4/V1/V3/A1/M2/_0_  (.A1(\V4/V1/V3/A1/M2/c1 ),
    .A2(\V4/V1/V3/A1/M2/c2 ),
    .ZN(\V4/V1/V3/A1/c2 ));
 AND2_X1 \V4/V1/V3/A1/M3/M1/_0_  (.A1(\V4/V1/V3/v2 [2]),
    .A2(\V4/V1/V3/v3 [2]),
    .ZN(\V4/V1/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M3/M1/_1_  (.A(\V4/V1/V3/v2 [2]),
    .B(\V4/V1/V3/v3 [2]),
    .Z(\V4/V1/V3/A1/M3/s1 ));
 AND2_X1 \V4/V1/V3/A1/M3/M2/_0_  (.A1(\V4/V1/V3/A1/M3/s1 ),
    .A2(\V4/V1/V3/A1/c2 ),
    .ZN(\V4/V1/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M3/M2/_1_  (.A(\V4/V1/V3/A1/M3/s1 ),
    .B(\V4/V1/V3/A1/c2 ),
    .Z(\V4/V1/V3/s1 [2]));
 OR2_X1 \V4/V1/V3/A1/M3/_0_  (.A1(\V4/V1/V3/A1/M3/c1 ),
    .A2(\V4/V1/V3/A1/M3/c2 ),
    .ZN(\V4/V1/V3/A1/c3 ));
 AND2_X1 \V4/V1/V3/A1/M4/M1/_0_  (.A1(\V4/V1/V3/v2 [3]),
    .A2(\V4/V1/V3/v3 [3]),
    .ZN(\V4/V1/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A1/M4/M1/_1_  (.A(\V4/V1/V3/v2 [3]),
    .B(\V4/V1/V3/v3 [3]),
    .Z(\V4/V1/V3/A1/M4/s1 ));
 AND2_X1 \V4/V1/V3/A1/M4/M2/_0_  (.A1(\V4/V1/V3/A1/M4/s1 ),
    .A2(\V4/V1/V3/A1/c3 ),
    .ZN(\V4/V1/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A1/M4/M2/_1_  (.A(\V4/V1/V3/A1/M4/s1 ),
    .B(\V4/V1/V3/A1/c3 ),
    .Z(\V4/V1/V3/s1 [3]));
 OR2_X1 \V4/V1/V3/A1/M4/_0_  (.A1(\V4/V1/V3/A1/M4/c1 ),
    .A2(\V4/V1/V3/A1/M4/c2 ),
    .ZN(\V4/V1/V3/c1 ));
 AND2_X1 \V4/V1/V3/A2/M1/M1/_0_  (.A1(\V4/V1/V3/s1 [0]),
    .A2(\V4/V1/V3/v1 [2]),
    .ZN(\V4/V1/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M1/M1/_1_  (.A(\V4/V1/V3/s1 [0]),
    .B(\V4/V1/V3/v1 [2]),
    .Z(\V4/V1/V3/A2/M1/s1 ));
 AND2_X1 \V4/V1/V3/A2/M1/M2/_0_  (.A1(\V4/V1/V3/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V1/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M1/M2/_1_  (.A(\V4/V1/V3/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/v3 [2]));
 OR2_X1 \V4/V1/V3/A2/M1/_0_  (.A1(\V4/V1/V3/A2/M1/c1 ),
    .A2(\V4/V1/V3/A2/M1/c2 ),
    .ZN(\V4/V1/V3/A2/c1 ));
 AND2_X1 \V4/V1/V3/A2/M2/M1/_0_  (.A1(\V4/V1/V3/s1 [1]),
    .A2(\V4/V1/V3/v1 [3]),
    .ZN(\V4/V1/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M2/M1/_1_  (.A(\V4/V1/V3/s1 [1]),
    .B(\V4/V1/V3/v1 [3]),
    .Z(\V4/V1/V3/A2/M2/s1 ));
 AND2_X1 \V4/V1/V3/A2/M2/M2/_0_  (.A1(\V4/V1/V3/A2/M2/s1 ),
    .A2(\V4/V1/V3/A2/c1 ),
    .ZN(\V4/V1/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M2/M2/_1_  (.A(\V4/V1/V3/A2/M2/s1 ),
    .B(\V4/V1/V3/A2/c1 ),
    .Z(\V4/V1/v3 [3]));
 OR2_X1 \V4/V1/V3/A2/M2/_0_  (.A1(\V4/V1/V3/A2/M2/c1 ),
    .A2(\V4/V1/V3/A2/M2/c2 ),
    .ZN(\V4/V1/V3/A2/c2 ));
 AND2_X1 \V4/V1/V3/A2/M3/M1/_0_  (.A1(\V4/V1/V3/s1 [2]),
    .A2(net10),
    .ZN(\V4/V1/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M3/M1/_1_  (.A(\V4/V1/V3/s1 [2]),
    .B(net10),
    .Z(\V4/V1/V3/A2/M3/s1 ));
 AND2_X1 \V4/V1/V3/A2/M3/M2/_0_  (.A1(\V4/V1/V3/A2/M3/s1 ),
    .A2(\V4/V1/V3/A2/c2 ),
    .ZN(\V4/V1/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M3/M2/_1_  (.A(\V4/V1/V3/A2/M3/s1 ),
    .B(\V4/V1/V3/A2/c2 ),
    .Z(\V4/V1/V3/s2 [2]));
 OR2_X1 \V4/V1/V3/A2/M3/_0_  (.A1(\V4/V1/V3/A2/M3/c1 ),
    .A2(\V4/V1/V3/A2/M3/c2 ),
    .ZN(\V4/V1/V3/A2/c3 ));
 AND2_X1 \V4/V1/V3/A2/M4/M1/_0_  (.A1(\V4/V1/V3/s1 [3]),
    .A2(net1),
    .ZN(\V4/V1/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A2/M4/M1/_1_  (.A(\V4/V1/V3/s1 [3]),
    .B(net1),
    .Z(\V4/V1/V3/A2/M4/s1 ));
 AND2_X1 \V4/V1/V3/A2/M4/M2/_0_  (.A1(\V4/V1/V3/A2/M4/s1 ),
    .A2(\V4/V1/V3/A2/c3 ),
    .ZN(\V4/V1/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A2/M4/M2/_1_  (.A(\V4/V1/V3/A2/M4/s1 ),
    .B(\V4/V1/V3/A2/c3 ),
    .Z(\V4/V1/V3/s2 [3]));
 OR2_X1 \V4/V1/V3/A2/M4/_0_  (.A1(\V4/V1/V3/A2/M4/c1 ),
    .A2(\V4/V1/V3/A2/M4/c2 ),
    .ZN(\V4/V1/V3/c2 ));
 AND2_X1 \V4/V1/V3/A3/M1/M1/_0_  (.A1(\V4/V1/V3/v4 [0]),
    .A2(\V4/V1/V3/s2 [2]),
    .ZN(\V4/V1/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M1/M1/_1_  (.A(\V4/V1/V3/v4 [0]),
    .B(\V4/V1/V3/s2 [2]),
    .Z(\V4/V1/V3/A3/M1/s1 ));
 AND2_X1 \V4/V1/V3/A3/M1/M2/_0_  (.A1(\V4/V1/V3/A3/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V1/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M1/M2/_1_  (.A(\V4/V1/V3/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/v3 [4]));
 OR2_X1 \V4/V1/V3/A3/M1/_0_  (.A1(\V4/V1/V3/A3/M1/c1 ),
    .A2(\V4/V1/V3/A3/M1/c2 ),
    .ZN(\V4/V1/V3/A3/c1 ));
 AND2_X1 \V4/V1/V3/A3/M2/M1/_0_  (.A1(\V4/V1/V3/v4 [1]),
    .A2(\V4/V1/V3/s2 [3]),
    .ZN(\V4/V1/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M2/M1/_1_  (.A(\V4/V1/V3/v4 [1]),
    .B(\V4/V1/V3/s2 [3]),
    .Z(\V4/V1/V3/A3/M2/s1 ));
 AND2_X1 \V4/V1/V3/A3/M2/M2/_0_  (.A1(\V4/V1/V3/A3/M2/s1 ),
    .A2(\V4/V1/V3/A3/c1 ),
    .ZN(\V4/V1/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M2/M2/_1_  (.A(\V4/V1/V3/A3/M2/s1 ),
    .B(\V4/V1/V3/A3/c1 ),
    .Z(\V4/V1/v3 [5]));
 OR2_X1 \V4/V1/V3/A3/M2/_0_  (.A1(\V4/V1/V3/A3/M2/c1 ),
    .A2(\V4/V1/V3/A3/M2/c2 ),
    .ZN(\V4/V1/V3/A3/c2 ));
 AND2_X1 \V4/V1/V3/A3/M3/M1/_0_  (.A1(\V4/V1/V3/v4 [2]),
    .A2(\V4/V1/V3/c3 ),
    .ZN(\V4/V1/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M3/M1/_1_  (.A(\V4/V1/V3/v4 [2]),
    .B(\V4/V1/V3/c3 ),
    .Z(\V4/V1/V3/A3/M3/s1 ));
 AND2_X1 \V4/V1/V3/A3/M3/M2/_0_  (.A1(\V4/V1/V3/A3/M3/s1 ),
    .A2(\V4/V1/V3/A3/c2 ),
    .ZN(\V4/V1/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M3/M2/_1_  (.A(\V4/V1/V3/A3/M3/s1 ),
    .B(\V4/V1/V3/A3/c2 ),
    .Z(\V4/V1/v3 [6]));
 OR2_X1 \V4/V1/V3/A3/M3/_0_  (.A1(\V4/V1/V3/A3/M3/c1 ),
    .A2(\V4/V1/V3/A3/M3/c2 ),
    .ZN(\V4/V1/V3/A3/c3 ));
 AND2_X1 \V4/V1/V3/A3/M4/M1/_0_  (.A1(\V4/V1/V3/v4 [3]),
    .A2(net1),
    .ZN(\V4/V1/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V3/A3/M4/M1/_1_  (.A(\V4/V1/V3/v4 [3]),
    .B(net1),
    .Z(\V4/V1/V3/A3/M4/s1 ));
 AND2_X1 \V4/V1/V3/A3/M4/M2/_0_  (.A1(\V4/V1/V3/A3/M4/s1 ),
    .A2(\V4/V1/V3/A3/c3 ),
    .ZN(\V4/V1/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V3/A3/M4/M2/_1_  (.A(\V4/V1/V3/A3/M4/s1 ),
    .B(\V4/V1/V3/A3/c3 ),
    .Z(\V4/V1/v3 [7]));
 OR2_X1 \V4/V1/V3/A3/M4/_0_  (.A1(\V4/V1/V3/A3/M4/c1 ),
    .A2(\V4/V1/V3/A3/M4/c2 ),
    .ZN(\V4/V1/V3/overflow ));
 AND2_X1 \V4/V1/V3/V1/HA1/_0_  (.A1(\V4/V1/V3/V1/w2 ),
    .A2(\V4/V1/V3/V1/w1 ),
    .ZN(\V4/V1/V3/V1/w4 ));
 XOR2_X2 \V4/V1/V3/V1/HA1/_1_  (.A(\V4/V1/V3/V1/w2 ),
    .B(\V4/V1/V3/V1/w1 ),
    .Z(\V4/V1/v3 [1]));
 AND2_X1 \V4/V1/V3/V1/HA2/_0_  (.A1(\V4/V1/V3/V1/w4 ),
    .A2(\V4/V1/V3/V1/w3 ),
    .ZN(\V4/V1/V3/v1 [3]));
 XOR2_X2 \V4/V1/V3/V1/HA2/_1_  (.A(\V4/V1/V3/V1/w4 ),
    .B(\V4/V1/V3/V1/w3 ),
    .Z(\V4/V1/V3/v1 [2]));
 AND2_X1 \V4/V1/V3/V1/_0_  (.A1(net41),
    .A2(B[20]),
    .ZN(\V4/V1/v3 [0]));
 AND2_X1 \V4/V1/V3/V1/_1_  (.A1(net41),
    .A2(B[21]),
    .ZN(\V4/V1/V3/V1/w1 ));
 AND2_X1 \V4/V1/V3/V1/_2_  (.A1(B[20]),
    .A2(net40),
    .ZN(\V4/V1/V3/V1/w2 ));
 AND2_X1 \V4/V1/V3/V1/_3_  (.A1(B[21]),
    .A2(net40),
    .ZN(\V4/V1/V3/V1/w3 ));
 AND2_X1 \V4/V1/V3/V2/HA1/_0_  (.A1(\V4/V1/V3/V2/w2 ),
    .A2(\V4/V1/V3/V2/w1 ),
    .ZN(\V4/V1/V3/V2/w4 ));
 XOR2_X2 \V4/V1/V3/V2/HA1/_1_  (.A(\V4/V1/V3/V2/w2 ),
    .B(\V4/V1/V3/V2/w1 ),
    .Z(\V4/V1/V3/v2 [1]));
 AND2_X1 \V4/V1/V3/V2/HA2/_0_  (.A1(\V4/V1/V3/V2/w4 ),
    .A2(\V4/V1/V3/V2/w3 ),
    .ZN(\V4/V1/V3/v2 [3]));
 XOR2_X2 \V4/V1/V3/V2/HA2/_1_  (.A(\V4/V1/V3/V2/w4 ),
    .B(\V4/V1/V3/V2/w3 ),
    .Z(\V4/V1/V3/v2 [2]));
 AND2_X1 \V4/V1/V3/V2/_0_  (.A1(net39),
    .A2(B[20]),
    .ZN(\V4/V1/V3/v2 [0]));
 AND2_X1 \V4/V1/V3/V2/_1_  (.A1(net39),
    .A2(B[21]),
    .ZN(\V4/V1/V3/V2/w1 ));
 AND2_X1 \V4/V1/V3/V2/_2_  (.A1(B[20]),
    .A2(net38),
    .ZN(\V4/V1/V3/V2/w2 ));
 AND2_X1 \V4/V1/V3/V2/_3_  (.A1(B[21]),
    .A2(net38),
    .ZN(\V4/V1/V3/V2/w3 ));
 AND2_X1 \V4/V1/V3/V3/HA1/_0_  (.A1(\V4/V1/V3/V3/w2 ),
    .A2(\V4/V1/V3/V3/w1 ),
    .ZN(\V4/V1/V3/V3/w4 ));
 XOR2_X2 \V4/V1/V3/V3/HA1/_1_  (.A(\V4/V1/V3/V3/w2 ),
    .B(\V4/V1/V3/V3/w1 ),
    .Z(\V4/V1/V3/v3 [1]));
 AND2_X1 \V4/V1/V3/V3/HA2/_0_  (.A1(\V4/V1/V3/V3/w4 ),
    .A2(\V4/V1/V3/V3/w3 ),
    .ZN(\V4/V1/V3/v3 [3]));
 XOR2_X2 \V4/V1/V3/V3/HA2/_1_  (.A(\V4/V1/V3/V3/w4 ),
    .B(\V4/V1/V3/V3/w3 ),
    .Z(\V4/V1/V3/v3 [2]));
 AND2_X1 \V4/V1/V3/V3/_0_  (.A1(net41),
    .A2(net16),
    .ZN(\V4/V1/V3/v3 [0]));
 AND2_X1 \V4/V1/V3/V3/_1_  (.A1(net41),
    .A2(net15),
    .ZN(\V4/V1/V3/V3/w1 ));
 AND2_X1 \V4/V1/V3/V3/_2_  (.A1(net16),
    .A2(net40),
    .ZN(\V4/V1/V3/V3/w2 ));
 AND2_X1 \V4/V1/V3/V3/_3_  (.A1(net15),
    .A2(net40),
    .ZN(\V4/V1/V3/V3/w3 ));
 AND2_X1 \V4/V1/V3/V4/HA1/_0_  (.A1(\V4/V1/V3/V4/w2 ),
    .A2(\V4/V1/V3/V4/w1 ),
    .ZN(\V4/V1/V3/V4/w4 ));
 XOR2_X2 \V4/V1/V3/V4/HA1/_1_  (.A(\V4/V1/V3/V4/w2 ),
    .B(\V4/V1/V3/V4/w1 ),
    .Z(\V4/V1/V3/v4 [1]));
 AND2_X1 \V4/V1/V3/V4/HA2/_0_  (.A1(\V4/V1/V3/V4/w4 ),
    .A2(\V4/V1/V3/V4/w3 ),
    .ZN(\V4/V1/V3/v4 [3]));
 XOR2_X2 \V4/V1/V3/V4/HA2/_1_  (.A(\V4/V1/V3/V4/w4 ),
    .B(\V4/V1/V3/V4/w3 ),
    .Z(\V4/V1/V3/v4 [2]));
 AND2_X1 \V4/V1/V3/V4/_0_  (.A1(net39),
    .A2(net16),
    .ZN(\V4/V1/V3/v4 [0]));
 AND2_X1 \V4/V1/V3/V4/_1_  (.A1(net39),
    .A2(net15),
    .ZN(\V4/V1/V3/V4/w1 ));
 AND2_X1 \V4/V1/V3/V4/_2_  (.A1(net16),
    .A2(net38),
    .ZN(\V4/V1/V3/V4/w2 ));
 AND2_X1 \V4/V1/V3/V4/_3_  (.A1(net15),
    .A2(net38),
    .ZN(\V4/V1/V3/V4/w3 ));
 OR2_X1 \V4/V1/V3/_0_  (.A1(\V4/V1/V3/c1 ),
    .A2(\V4/V1/V3/c2 ),
    .ZN(\V4/V1/V3/c3 ));
 AND2_X1 \V4/V1/V4/A1/M1/M1/_0_  (.A1(\V4/V1/V4/v2 [0]),
    .A2(\V4/V1/V4/v3 [0]),
    .ZN(\V4/V1/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M1/M1/_1_  (.A(\V4/V1/V4/v2 [0]),
    .B(\V4/V1/V4/v3 [0]),
    .Z(\V4/V1/V4/A1/M1/s1 ));
 AND2_X1 \V4/V1/V4/A1/M1/M2/_0_  (.A1(\V4/V1/V4/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V1/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M1/M2/_1_  (.A(\V4/V1/V4/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V1/V4/s1 [0]));
 OR2_X1 \V4/V1/V4/A1/M1/_0_  (.A1(\V4/V1/V4/A1/M1/c1 ),
    .A2(\V4/V1/V4/A1/M1/c2 ),
    .ZN(\V4/V1/V4/A1/c1 ));
 AND2_X1 \V4/V1/V4/A1/M2/M1/_0_  (.A1(\V4/V1/V4/v2 [1]),
    .A2(\V4/V1/V4/v3 [1]),
    .ZN(\V4/V1/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M2/M1/_1_  (.A(\V4/V1/V4/v2 [1]),
    .B(\V4/V1/V4/v3 [1]),
    .Z(\V4/V1/V4/A1/M2/s1 ));
 AND2_X1 \V4/V1/V4/A1/M2/M2/_0_  (.A1(\V4/V1/V4/A1/M2/s1 ),
    .A2(\V4/V1/V4/A1/c1 ),
    .ZN(\V4/V1/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M2/M2/_1_  (.A(\V4/V1/V4/A1/M2/s1 ),
    .B(\V4/V1/V4/A1/c1 ),
    .Z(\V4/V1/V4/s1 [1]));
 OR2_X1 \V4/V1/V4/A1/M2/_0_  (.A1(\V4/V1/V4/A1/M2/c1 ),
    .A2(\V4/V1/V4/A1/M2/c2 ),
    .ZN(\V4/V1/V4/A1/c2 ));
 AND2_X1 \V4/V1/V4/A1/M3/M1/_0_  (.A1(\V4/V1/V4/v2 [2]),
    .A2(\V4/V1/V4/v3 [2]),
    .ZN(\V4/V1/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M3/M1/_1_  (.A(\V4/V1/V4/v2 [2]),
    .B(\V4/V1/V4/v3 [2]),
    .Z(\V4/V1/V4/A1/M3/s1 ));
 AND2_X1 \V4/V1/V4/A1/M3/M2/_0_  (.A1(\V4/V1/V4/A1/M3/s1 ),
    .A2(\V4/V1/V4/A1/c2 ),
    .ZN(\V4/V1/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M3/M2/_1_  (.A(\V4/V1/V4/A1/M3/s1 ),
    .B(\V4/V1/V4/A1/c2 ),
    .Z(\V4/V1/V4/s1 [2]));
 OR2_X1 \V4/V1/V4/A1/M3/_0_  (.A1(\V4/V1/V4/A1/M3/c1 ),
    .A2(\V4/V1/V4/A1/M3/c2 ),
    .ZN(\V4/V1/V4/A1/c3 ));
 AND2_X1 \V4/V1/V4/A1/M4/M1/_0_  (.A1(\V4/V1/V4/v2 [3]),
    .A2(\V4/V1/V4/v3 [3]),
    .ZN(\V4/V1/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A1/M4/M1/_1_  (.A(\V4/V1/V4/v2 [3]),
    .B(\V4/V1/V4/v3 [3]),
    .Z(\V4/V1/V4/A1/M4/s1 ));
 AND2_X1 \V4/V1/V4/A1/M4/M2/_0_  (.A1(\V4/V1/V4/A1/M4/s1 ),
    .A2(\V4/V1/V4/A1/c3 ),
    .ZN(\V4/V1/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A1/M4/M2/_1_  (.A(\V4/V1/V4/A1/M4/s1 ),
    .B(\V4/V1/V4/A1/c3 ),
    .Z(\V4/V1/V4/s1 [3]));
 OR2_X1 \V4/V1/V4/A1/M4/_0_  (.A1(\V4/V1/V4/A1/M4/c1 ),
    .A2(\V4/V1/V4/A1/M4/c2 ),
    .ZN(\V4/V1/V4/c1 ));
 AND2_X1 \V4/V1/V4/A2/M1/M1/_0_  (.A1(\V4/V1/V4/s1 [0]),
    .A2(\V4/V1/V4/v1 [2]),
    .ZN(\V4/V1/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M1/M1/_1_  (.A(\V4/V1/V4/s1 [0]),
    .B(\V4/V1/V4/v1 [2]),
    .Z(\V4/V1/V4/A2/M1/s1 ));
 AND2_X1 \V4/V1/V4/A2/M1/M2/_0_  (.A1(\V4/V1/V4/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V1/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M1/M2/_1_  (.A(\V4/V1/V4/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V1/v4 [2]));
 OR2_X1 \V4/V1/V4/A2/M1/_0_  (.A1(\V4/V1/V4/A2/M1/c1 ),
    .A2(\V4/V1/V4/A2/M1/c2 ),
    .ZN(\V4/V1/V4/A2/c1 ));
 AND2_X1 \V4/V1/V4/A2/M2/M1/_0_  (.A1(\V4/V1/V4/s1 [1]),
    .A2(\V4/V1/V4/v1 [3]),
    .ZN(\V4/V1/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M2/M1/_1_  (.A(\V4/V1/V4/s1 [1]),
    .B(\V4/V1/V4/v1 [3]),
    .Z(\V4/V1/V4/A2/M2/s1 ));
 AND2_X1 \V4/V1/V4/A2/M2/M2/_0_  (.A1(\V4/V1/V4/A2/M2/s1 ),
    .A2(\V4/V1/V4/A2/c1 ),
    .ZN(\V4/V1/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M2/M2/_1_  (.A(\V4/V1/V4/A2/M2/s1 ),
    .B(\V4/V1/V4/A2/c1 ),
    .Z(\V4/V1/v4 [3]));
 OR2_X1 \V4/V1/V4/A2/M2/_0_  (.A1(\V4/V1/V4/A2/M2/c1 ),
    .A2(\V4/V1/V4/A2/M2/c2 ),
    .ZN(\V4/V1/V4/A2/c2 ));
 AND2_X1 \V4/V1/V4/A2/M3/M1/_0_  (.A1(\V4/V1/V4/s1 [2]),
    .A2(net1),
    .ZN(\V4/V1/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M3/M1/_1_  (.A(\V4/V1/V4/s1 [2]),
    .B(net1),
    .Z(\V4/V1/V4/A2/M3/s1 ));
 AND2_X1 \V4/V1/V4/A2/M3/M2/_0_  (.A1(\V4/V1/V4/A2/M3/s1 ),
    .A2(\V4/V1/V4/A2/c2 ),
    .ZN(\V4/V1/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M3/M2/_1_  (.A(\V4/V1/V4/A2/M3/s1 ),
    .B(\V4/V1/V4/A2/c2 ),
    .Z(\V4/V1/V4/s2 [2]));
 OR2_X1 \V4/V1/V4/A2/M3/_0_  (.A1(\V4/V1/V4/A2/M3/c1 ),
    .A2(\V4/V1/V4/A2/M3/c2 ),
    .ZN(\V4/V1/V4/A2/c3 ));
 AND2_X1 \V4/V1/V4/A2/M4/M1/_0_  (.A1(\V4/V1/V4/s1 [3]),
    .A2(net1),
    .ZN(\V4/V1/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A2/M4/M1/_1_  (.A(\V4/V1/V4/s1 [3]),
    .B(net1),
    .Z(\V4/V1/V4/A2/M4/s1 ));
 AND2_X1 \V4/V1/V4/A2/M4/M2/_0_  (.A1(\V4/V1/V4/A2/M4/s1 ),
    .A2(\V4/V1/V4/A2/c3 ),
    .ZN(\V4/V1/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A2/M4/M2/_1_  (.A(\V4/V1/V4/A2/M4/s1 ),
    .B(\V4/V1/V4/A2/c3 ),
    .Z(\V4/V1/V4/s2 [3]));
 OR2_X1 \V4/V1/V4/A2/M4/_0_  (.A1(\V4/V1/V4/A2/M4/c1 ),
    .A2(\V4/V1/V4/A2/M4/c2 ),
    .ZN(\V4/V1/V4/c2 ));
 AND2_X1 \V4/V1/V4/A3/M1/M1/_0_  (.A1(\V4/V1/V4/v4 [0]),
    .A2(\V4/V1/V4/s2 [2]),
    .ZN(\V4/V1/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M1/M1/_1_  (.A(\V4/V1/V4/v4 [0]),
    .B(\V4/V1/V4/s2 [2]),
    .Z(\V4/V1/V4/A3/M1/s1 ));
 AND2_X1 \V4/V1/V4/A3/M1/M2/_0_  (.A1(\V4/V1/V4/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V1/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M1/M2/_1_  (.A(\V4/V1/V4/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V1/v4 [4]));
 OR2_X1 \V4/V1/V4/A3/M1/_0_  (.A1(\V4/V1/V4/A3/M1/c1 ),
    .A2(\V4/V1/V4/A3/M1/c2 ),
    .ZN(\V4/V1/V4/A3/c1 ));
 AND2_X1 \V4/V1/V4/A3/M2/M1/_0_  (.A1(\V4/V1/V4/v4 [1]),
    .A2(\V4/V1/V4/s2 [3]),
    .ZN(\V4/V1/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M2/M1/_1_  (.A(\V4/V1/V4/v4 [1]),
    .B(\V4/V1/V4/s2 [3]),
    .Z(\V4/V1/V4/A3/M2/s1 ));
 AND2_X1 \V4/V1/V4/A3/M2/M2/_0_  (.A1(\V4/V1/V4/A3/M2/s1 ),
    .A2(\V4/V1/V4/A3/c1 ),
    .ZN(\V4/V1/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M2/M2/_1_  (.A(\V4/V1/V4/A3/M2/s1 ),
    .B(\V4/V1/V4/A3/c1 ),
    .Z(\V4/V1/v4 [5]));
 OR2_X1 \V4/V1/V4/A3/M2/_0_  (.A1(\V4/V1/V4/A3/M2/c1 ),
    .A2(\V4/V1/V4/A3/M2/c2 ),
    .ZN(\V4/V1/V4/A3/c2 ));
 AND2_X1 \V4/V1/V4/A3/M3/M1/_0_  (.A1(\V4/V1/V4/v4 [2]),
    .A2(\V4/V1/V4/c3 ),
    .ZN(\V4/V1/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M3/M1/_1_  (.A(\V4/V1/V4/v4 [2]),
    .B(\V4/V1/V4/c3 ),
    .Z(\V4/V1/V4/A3/M3/s1 ));
 AND2_X1 \V4/V1/V4/A3/M3/M2/_0_  (.A1(\V4/V1/V4/A3/M3/s1 ),
    .A2(\V4/V1/V4/A3/c2 ),
    .ZN(\V4/V1/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M3/M2/_1_  (.A(\V4/V1/V4/A3/M3/s1 ),
    .B(\V4/V1/V4/A3/c2 ),
    .Z(\V4/V1/v4 [6]));
 OR2_X1 \V4/V1/V4/A3/M3/_0_  (.A1(\V4/V1/V4/A3/M3/c1 ),
    .A2(\V4/V1/V4/A3/M3/c2 ),
    .ZN(\V4/V1/V4/A3/c3 ));
 AND2_X1 \V4/V1/V4/A3/M4/M1/_0_  (.A1(\V4/V1/V4/v4 [3]),
    .A2(net1),
    .ZN(\V4/V1/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V1/V4/A3/M4/M1/_1_  (.A(\V4/V1/V4/v4 [3]),
    .B(net1),
    .Z(\V4/V1/V4/A3/M4/s1 ));
 AND2_X1 \V4/V1/V4/A3/M4/M2/_0_  (.A1(\V4/V1/V4/A3/M4/s1 ),
    .A2(\V4/V1/V4/A3/c3 ),
    .ZN(\V4/V1/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V1/V4/A3/M4/M2/_1_  (.A(\V4/V1/V4/A3/M4/s1 ),
    .B(\V4/V1/V4/A3/c3 ),
    .Z(\V4/V1/v4 [7]));
 OR2_X1 \V4/V1/V4/A3/M4/_0_  (.A1(\V4/V1/V4/A3/M4/c1 ),
    .A2(\V4/V1/V4/A3/M4/c2 ),
    .ZN(\V4/V1/V4/overflow ));
 AND2_X1 \V4/V1/V4/V1/HA1/_0_  (.A1(\V4/V1/V4/V1/w2 ),
    .A2(\V4/V1/V4/V1/w1 ),
    .ZN(\V4/V1/V4/V1/w4 ));
 XOR2_X2 \V4/V1/V4/V1/HA1/_1_  (.A(\V4/V1/V4/V1/w2 ),
    .B(\V4/V1/V4/V1/w1 ),
    .Z(\V4/V1/v4 [1]));
 AND2_X1 \V4/V1/V4/V1/HA2/_0_  (.A1(\V4/V1/V4/V1/w4 ),
    .A2(\V4/V1/V4/V1/w3 ),
    .ZN(\V4/V1/V4/v1 [3]));
 XOR2_X2 \V4/V1/V4/V1/HA2/_1_  (.A(\V4/V1/V4/V1/w4 ),
    .B(\V4/V1/V4/V1/w3 ),
    .Z(\V4/V1/V4/v1 [2]));
 AND2_X1 \V4/V1/V4/V1/_0_  (.A1(net37),
    .A2(net18),
    .ZN(\V4/V1/v4 [0]));
 AND2_X1 \V4/V1/V4/V1/_1_  (.A1(net37),
    .A2(net17),
    .ZN(\V4/V1/V4/V1/w1 ));
 AND2_X1 \V4/V1/V4/V1/_2_  (.A1(net18),
    .A2(net36),
    .ZN(\V4/V1/V4/V1/w2 ));
 AND2_X1 \V4/V1/V4/V1/_3_  (.A1(net17),
    .A2(net36),
    .ZN(\V4/V1/V4/V1/w3 ));
 AND2_X1 \V4/V1/V4/V2/HA1/_0_  (.A1(\V4/V1/V4/V2/w2 ),
    .A2(\V4/V1/V4/V2/w1 ),
    .ZN(\V4/V1/V4/V2/w4 ));
 XOR2_X2 \V4/V1/V4/V2/HA1/_1_  (.A(\V4/V1/V4/V2/w2 ),
    .B(\V4/V1/V4/V2/w1 ),
    .Z(\V4/V1/V4/v2 [1]));
 AND2_X1 \V4/V1/V4/V2/HA2/_0_  (.A1(\V4/V1/V4/V2/w4 ),
    .A2(\V4/V1/V4/V2/w3 ),
    .ZN(\V4/V1/V4/v2 [3]));
 XOR2_X2 \V4/V1/V4/V2/HA2/_1_  (.A(\V4/V1/V4/V2/w4 ),
    .B(\V4/V1/V4/V2/w3 ),
    .Z(\V4/V1/V4/v2 [2]));
 AND2_X1 \V4/V1/V4/V2/_0_  (.A1(net35),
    .A2(net18),
    .ZN(\V4/V1/V4/v2 [0]));
 AND2_X1 \V4/V1/V4/V2/_1_  (.A1(net35),
    .A2(net17),
    .ZN(\V4/V1/V4/V2/w1 ));
 AND2_X1 \V4/V1/V4/V2/_2_  (.A1(net18),
    .A2(net34),
    .ZN(\V4/V1/V4/V2/w2 ));
 AND2_X1 \V4/V1/V4/V2/_3_  (.A1(net17),
    .A2(net34),
    .ZN(\V4/V1/V4/V2/w3 ));
 AND2_X1 \V4/V1/V4/V3/HA1/_0_  (.A1(\V4/V1/V4/V3/w2 ),
    .A2(\V4/V1/V4/V3/w1 ),
    .ZN(\V4/V1/V4/V3/w4 ));
 XOR2_X2 \V4/V1/V4/V3/HA1/_1_  (.A(\V4/V1/V4/V3/w2 ),
    .B(\V4/V1/V4/V3/w1 ),
    .Z(\V4/V1/V4/v3 [1]));
 AND2_X1 \V4/V1/V4/V3/HA2/_0_  (.A1(\V4/V1/V4/V3/w4 ),
    .A2(\V4/V1/V4/V3/w3 ),
    .ZN(\V4/V1/V4/v3 [3]));
 XOR2_X2 \V4/V1/V4/V3/HA2/_1_  (.A(\V4/V1/V4/V3/w4 ),
    .B(\V4/V1/V4/V3/w3 ),
    .Z(\V4/V1/V4/v3 [2]));
 AND2_X1 \V4/V1/V4/V3/_0_  (.A1(net37),
    .A2(net16),
    .ZN(\V4/V1/V4/v3 [0]));
 AND2_X1 \V4/V1/V4/V3/_1_  (.A1(net37),
    .A2(net15),
    .ZN(\V4/V1/V4/V3/w1 ));
 AND2_X1 \V4/V1/V4/V3/_2_  (.A1(net16),
    .A2(net36),
    .ZN(\V4/V1/V4/V3/w2 ));
 AND2_X1 \V4/V1/V4/V3/_3_  (.A1(net15),
    .A2(net36),
    .ZN(\V4/V1/V4/V3/w3 ));
 AND2_X1 \V4/V1/V4/V4/HA1/_0_  (.A1(\V4/V1/V4/V4/w2 ),
    .A2(\V4/V1/V4/V4/w1 ),
    .ZN(\V4/V1/V4/V4/w4 ));
 XOR2_X2 \V4/V1/V4/V4/HA1/_1_  (.A(\V4/V1/V4/V4/w2 ),
    .B(\V4/V1/V4/V4/w1 ),
    .Z(\V4/V1/V4/v4 [1]));
 AND2_X1 \V4/V1/V4/V4/HA2/_0_  (.A1(\V4/V1/V4/V4/w4 ),
    .A2(\V4/V1/V4/V4/w3 ),
    .ZN(\V4/V1/V4/v4 [3]));
 XOR2_X2 \V4/V1/V4/V4/HA2/_1_  (.A(\V4/V1/V4/V4/w4 ),
    .B(\V4/V1/V4/V4/w3 ),
    .Z(\V4/V1/V4/v4 [2]));
 AND2_X1 \V4/V1/V4/V4/_0_  (.A1(net35),
    .A2(net16),
    .ZN(\V4/V1/V4/v4 [0]));
 AND2_X1 \V4/V1/V4/V4/_1_  (.A1(net35),
    .A2(net15),
    .ZN(\V4/V1/V4/V4/w1 ));
 AND2_X1 \V4/V1/V4/V4/_2_  (.A1(net16),
    .A2(net34),
    .ZN(\V4/V1/V4/V4/w2 ));
 AND2_X1 \V4/V1/V4/V4/_3_  (.A1(net15),
    .A2(net34),
    .ZN(\V4/V1/V4/V4/w3 ));
 OR2_X1 \V4/V1/V4/_0_  (.A1(\V4/V1/V4/c1 ),
    .A2(\V4/V1/V4/c2 ),
    .ZN(\V4/V1/V4/c3 ));
 OR2_X1 \V4/V1/_0_  (.A1(\V4/V1/c1 ),
    .A2(\V4/V1/c2 ),
    .ZN(\V4/V1/c3 ));
 AND2_X1 \V4/V2/A1/A1/M1/M1/_0_  (.A1(\V4/V2/v2 [0]),
    .A2(\V4/V2/v3 [0]),
    .ZN(\V4/V2/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M1/M1/_1_  (.A(\V4/V2/v2 [0]),
    .B(\V4/V2/v3 [0]),
    .Z(\V4/V2/A1/A1/M1/s1 ));
 AND2_X1 \V4/V2/A1/A1/M1/M2/_0_  (.A1(\V4/V2/A1/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M1/M2/_1_  (.A(\V4/V2/A1/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/s1 [0]));
 OR2_X1 \V4/V2/A1/A1/M1/_0_  (.A1(\V4/V2/A1/A1/M1/c1 ),
    .A2(\V4/V2/A1/A1/M1/c2 ),
    .ZN(\V4/V2/A1/A1/c1 ));
 AND2_X1 \V4/V2/A1/A1/M2/M1/_0_  (.A1(\V4/V2/v2 [1]),
    .A2(\V4/V2/v3 [1]),
    .ZN(\V4/V2/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M2/M1/_1_  (.A(\V4/V2/v2 [1]),
    .B(\V4/V2/v3 [1]),
    .Z(\V4/V2/A1/A1/M2/s1 ));
 AND2_X1 \V4/V2/A1/A1/M2/M2/_0_  (.A1(\V4/V2/A1/A1/M2/s1 ),
    .A2(\V4/V2/A1/A1/c1 ),
    .ZN(\V4/V2/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M2/M2/_1_  (.A(\V4/V2/A1/A1/M2/s1 ),
    .B(\V4/V2/A1/A1/c1 ),
    .Z(\V4/V2/s1 [1]));
 OR2_X1 \V4/V2/A1/A1/M2/_0_  (.A1(\V4/V2/A1/A1/M2/c1 ),
    .A2(\V4/V2/A1/A1/M2/c2 ),
    .ZN(\V4/V2/A1/A1/c2 ));
 AND2_X1 \V4/V2/A1/A1/M3/M1/_0_  (.A1(\V4/V2/v2 [2]),
    .A2(\V4/V2/v3 [2]),
    .ZN(\V4/V2/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M3/M1/_1_  (.A(\V4/V2/v2 [2]),
    .B(\V4/V2/v3 [2]),
    .Z(\V4/V2/A1/A1/M3/s1 ));
 AND2_X1 \V4/V2/A1/A1/M3/M2/_0_  (.A1(\V4/V2/A1/A1/M3/s1 ),
    .A2(\V4/V2/A1/A1/c2 ),
    .ZN(\V4/V2/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M3/M2/_1_  (.A(\V4/V2/A1/A1/M3/s1 ),
    .B(\V4/V2/A1/A1/c2 ),
    .Z(\V4/V2/s1 [2]));
 OR2_X1 \V4/V2/A1/A1/M3/_0_  (.A1(\V4/V2/A1/A1/M3/c1 ),
    .A2(\V4/V2/A1/A1/M3/c2 ),
    .ZN(\V4/V2/A1/A1/c3 ));
 AND2_X1 \V4/V2/A1/A1/M4/M1/_0_  (.A1(\V4/V2/v2 [3]),
    .A2(\V4/V2/v3 [3]),
    .ZN(\V4/V2/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A1/A1/M4/M1/_1_  (.A(\V4/V2/v2 [3]),
    .B(\V4/V2/v3 [3]),
    .Z(\V4/V2/A1/A1/M4/s1 ));
 AND2_X1 \V4/V2/A1/A1/M4/M2/_0_  (.A1(\V4/V2/A1/A1/M4/s1 ),
    .A2(\V4/V2/A1/A1/c3 ),
    .ZN(\V4/V2/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A1/A1/M4/M2/_1_  (.A(\V4/V2/A1/A1/M4/s1 ),
    .B(\V4/V2/A1/A1/c3 ),
    .Z(\V4/V2/s1 [3]));
 OR2_X1 \V4/V2/A1/A1/M4/_0_  (.A1(\V4/V2/A1/A1/M4/c1 ),
    .A2(\V4/V2/A1/A1/M4/c2 ),
    .ZN(\V4/V2/A1/c1 ));
 AND2_X1 \V4/V2/A1/A2/M1/M1/_0_  (.A1(\V4/V2/v2 [4]),
    .A2(\V4/V2/v3 [4]),
    .ZN(\V4/V2/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M1/M1/_1_  (.A(\V4/V2/v2 [4]),
    .B(\V4/V2/v3 [4]),
    .Z(\V4/V2/A1/A2/M1/s1 ));
 AND2_X1 \V4/V2/A1/A2/M1/M2/_0_  (.A1(\V4/V2/A1/A2/M1/s1 ),
    .A2(\V4/V2/A1/c1 ),
    .ZN(\V4/V2/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M1/M2/_1_  (.A(\V4/V2/A1/A2/M1/s1 ),
    .B(\V4/V2/A1/c1 ),
    .Z(\V4/V2/s1 [4]));
 OR2_X1 \V4/V2/A1/A2/M1/_0_  (.A1(\V4/V2/A1/A2/M1/c1 ),
    .A2(\V4/V2/A1/A2/M1/c2 ),
    .ZN(\V4/V2/A1/A2/c1 ));
 AND2_X1 \V4/V2/A1/A2/M2/M1/_0_  (.A1(\V4/V2/v2 [5]),
    .A2(\V4/V2/v3 [5]),
    .ZN(\V4/V2/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M2/M1/_1_  (.A(\V4/V2/v2 [5]),
    .B(\V4/V2/v3 [5]),
    .Z(\V4/V2/A1/A2/M2/s1 ));
 AND2_X1 \V4/V2/A1/A2/M2/M2/_0_  (.A1(\V4/V2/A1/A2/M2/s1 ),
    .A2(\V4/V2/A1/A2/c1 ),
    .ZN(\V4/V2/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M2/M2/_1_  (.A(\V4/V2/A1/A2/M2/s1 ),
    .B(\V4/V2/A1/A2/c1 ),
    .Z(\V4/V2/s1 [5]));
 OR2_X1 \V4/V2/A1/A2/M2/_0_  (.A1(\V4/V2/A1/A2/M2/c1 ),
    .A2(\V4/V2/A1/A2/M2/c2 ),
    .ZN(\V4/V2/A1/A2/c2 ));
 AND2_X1 \V4/V2/A1/A2/M3/M1/_0_  (.A1(\V4/V2/v2 [6]),
    .A2(\V4/V2/v3 [6]),
    .ZN(\V4/V2/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M3/M1/_1_  (.A(\V4/V2/v2 [6]),
    .B(\V4/V2/v3 [6]),
    .Z(\V4/V2/A1/A2/M3/s1 ));
 AND2_X1 \V4/V2/A1/A2/M3/M2/_0_  (.A1(\V4/V2/A1/A2/M3/s1 ),
    .A2(\V4/V2/A1/A2/c2 ),
    .ZN(\V4/V2/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M3/M2/_1_  (.A(\V4/V2/A1/A2/M3/s1 ),
    .B(\V4/V2/A1/A2/c2 ),
    .Z(\V4/V2/s1 [6]));
 OR2_X1 \V4/V2/A1/A2/M3/_0_  (.A1(\V4/V2/A1/A2/M3/c1 ),
    .A2(\V4/V2/A1/A2/M3/c2 ),
    .ZN(\V4/V2/A1/A2/c3 ));
 AND2_X1 \V4/V2/A1/A2/M4/M1/_0_  (.A1(\V4/V2/v2 [7]),
    .A2(\V4/V2/v3 [7]),
    .ZN(\V4/V2/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A1/A2/M4/M1/_1_  (.A(\V4/V2/v2 [7]),
    .B(\V4/V2/v3 [7]),
    .Z(\V4/V2/A1/A2/M4/s1 ));
 AND2_X1 \V4/V2/A1/A2/M4/M2/_0_  (.A1(\V4/V2/A1/A2/M4/s1 ),
    .A2(\V4/V2/A1/A2/c3 ),
    .ZN(\V4/V2/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A1/A2/M4/M2/_1_  (.A(\V4/V2/A1/A2/M4/s1 ),
    .B(\V4/V2/A1/A2/c3 ),
    .Z(\V4/V2/s1 [7]));
 OR2_X1 \V4/V2/A1/A2/M4/_0_  (.A1(\V4/V2/A1/A2/M4/c1 ),
    .A2(\V4/V2/A1/A2/M4/c2 ),
    .ZN(\V4/V2/c1 ));
 AND2_X1 \V4/V2/A2/A1/M1/M1/_0_  (.A1(\V4/V2/s1 [0]),
    .A2(\V4/V2/v1 [4]),
    .ZN(\V4/V2/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M1/M1/_1_  (.A(\V4/V2/s1 [0]),
    .B(\V4/V2/v1 [4]),
    .Z(\V4/V2/A2/A1/M1/s1 ));
 AND2_X1 \V4/V2/A2/A1/M1/M2/_0_  (.A1(\V4/V2/A2/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M1/M2/_1_  (.A(\V4/V2/A2/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/v2 [4]));
 OR2_X1 \V4/V2/A2/A1/M1/_0_  (.A1(\V4/V2/A2/A1/M1/c1 ),
    .A2(\V4/V2/A2/A1/M1/c2 ),
    .ZN(\V4/V2/A2/A1/c1 ));
 AND2_X1 \V4/V2/A2/A1/M2/M1/_0_  (.A1(\V4/V2/s1 [1]),
    .A2(\V4/V2/v1 [5]),
    .ZN(\V4/V2/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M2/M1/_1_  (.A(\V4/V2/s1 [1]),
    .B(\V4/V2/v1 [5]),
    .Z(\V4/V2/A2/A1/M2/s1 ));
 AND2_X1 \V4/V2/A2/A1/M2/M2/_0_  (.A1(\V4/V2/A2/A1/M2/s1 ),
    .A2(\V4/V2/A2/A1/c1 ),
    .ZN(\V4/V2/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M2/M2/_1_  (.A(\V4/V2/A2/A1/M2/s1 ),
    .B(\V4/V2/A2/A1/c1 ),
    .Z(\V4/v2 [5]));
 OR2_X1 \V4/V2/A2/A1/M2/_0_  (.A1(\V4/V2/A2/A1/M2/c1 ),
    .A2(\V4/V2/A2/A1/M2/c2 ),
    .ZN(\V4/V2/A2/A1/c2 ));
 AND2_X1 \V4/V2/A2/A1/M3/M1/_0_  (.A1(\V4/V2/s1 [2]),
    .A2(\V4/V2/v1 [6]),
    .ZN(\V4/V2/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M3/M1/_1_  (.A(\V4/V2/s1 [2]),
    .B(\V4/V2/v1 [6]),
    .Z(\V4/V2/A2/A1/M3/s1 ));
 AND2_X1 \V4/V2/A2/A1/M3/M2/_0_  (.A1(\V4/V2/A2/A1/M3/s1 ),
    .A2(\V4/V2/A2/A1/c2 ),
    .ZN(\V4/V2/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M3/M2/_1_  (.A(\V4/V2/A2/A1/M3/s1 ),
    .B(\V4/V2/A2/A1/c2 ),
    .Z(\V4/v2 [6]));
 OR2_X1 \V4/V2/A2/A1/M3/_0_  (.A1(\V4/V2/A2/A1/M3/c1 ),
    .A2(\V4/V2/A2/A1/M3/c2 ),
    .ZN(\V4/V2/A2/A1/c3 ));
 AND2_X1 \V4/V2/A2/A1/M4/M1/_0_  (.A1(\V4/V2/s1 [3]),
    .A2(\V4/V2/v1 [7]),
    .ZN(\V4/V2/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A2/A1/M4/M1/_1_  (.A(\V4/V2/s1 [3]),
    .B(\V4/V2/v1 [7]),
    .Z(\V4/V2/A2/A1/M4/s1 ));
 AND2_X1 \V4/V2/A2/A1/M4/M2/_0_  (.A1(\V4/V2/A2/A1/M4/s1 ),
    .A2(\V4/V2/A2/A1/c3 ),
    .ZN(\V4/V2/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A2/A1/M4/M2/_1_  (.A(\V4/V2/A2/A1/M4/s1 ),
    .B(\V4/V2/A2/A1/c3 ),
    .Z(\V4/v2 [7]));
 OR2_X1 \V4/V2/A2/A1/M4/_0_  (.A1(\V4/V2/A2/A1/M4/c1 ),
    .A2(\V4/V2/A2/A1/M4/c2 ),
    .ZN(\V4/V2/A2/c1 ));
 AND2_X1 \V4/V2/A2/A2/M1/M1/_0_  (.A1(\V4/V2/s1 [4]),
    .A2(net1),
    .ZN(\V4/V2/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M1/M1/_1_  (.A(\V4/V2/s1 [4]),
    .B(net1),
    .Z(\V4/V2/A2/A2/M1/s1 ));
 AND2_X1 \V4/V2/A2/A2/M1/M2/_0_  (.A1(\V4/V2/A2/A2/M1/s1 ),
    .A2(\V4/V2/A2/c1 ),
    .ZN(\V4/V2/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M1/M2/_1_  (.A(\V4/V2/A2/A2/M1/s1 ),
    .B(\V4/V2/A2/c1 ),
    .Z(\V4/V2/s2 [4]));
 OR2_X1 \V4/V2/A2/A2/M1/_0_  (.A1(\V4/V2/A2/A2/M1/c1 ),
    .A2(\V4/V2/A2/A2/M1/c2 ),
    .ZN(\V4/V2/A2/A2/c1 ));
 AND2_X1 \V4/V2/A2/A2/M2/M1/_0_  (.A1(\V4/V2/s1 [5]),
    .A2(net1),
    .ZN(\V4/V2/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M2/M1/_1_  (.A(\V4/V2/s1 [5]),
    .B(net1),
    .Z(\V4/V2/A2/A2/M2/s1 ));
 AND2_X1 \V4/V2/A2/A2/M2/M2/_0_  (.A1(\V4/V2/A2/A2/M2/s1 ),
    .A2(\V4/V2/A2/A2/c1 ),
    .ZN(\V4/V2/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M2/M2/_1_  (.A(\V4/V2/A2/A2/M2/s1 ),
    .B(\V4/V2/A2/A2/c1 ),
    .Z(\V4/V2/s2 [5]));
 OR2_X1 \V4/V2/A2/A2/M2/_0_  (.A1(\V4/V2/A2/A2/M2/c1 ),
    .A2(\V4/V2/A2/A2/M2/c2 ),
    .ZN(\V4/V2/A2/A2/c2 ));
 AND2_X1 \V4/V2/A2/A2/M3/M1/_0_  (.A1(\V4/V2/s1 [6]),
    .A2(net1),
    .ZN(\V4/V2/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M3/M1/_1_  (.A(\V4/V2/s1 [6]),
    .B(net1),
    .Z(\V4/V2/A2/A2/M3/s1 ));
 AND2_X1 \V4/V2/A2/A2/M3/M2/_0_  (.A1(\V4/V2/A2/A2/M3/s1 ),
    .A2(\V4/V2/A2/A2/c2 ),
    .ZN(\V4/V2/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M3/M2/_1_  (.A(\V4/V2/A2/A2/M3/s1 ),
    .B(\V4/V2/A2/A2/c2 ),
    .Z(\V4/V2/s2 [6]));
 OR2_X1 \V4/V2/A2/A2/M3/_0_  (.A1(\V4/V2/A2/A2/M3/c1 ),
    .A2(\V4/V2/A2/A2/M3/c2 ),
    .ZN(\V4/V2/A2/A2/c3 ));
 AND2_X1 \V4/V2/A2/A2/M4/M1/_0_  (.A1(\V4/V2/s1 [7]),
    .A2(net1),
    .ZN(\V4/V2/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A2/A2/M4/M1/_1_  (.A(\V4/V2/s1 [7]),
    .B(net1),
    .Z(\V4/V2/A2/A2/M4/s1 ));
 AND2_X1 \V4/V2/A2/A2/M4/M2/_0_  (.A1(\V4/V2/A2/A2/M4/s1 ),
    .A2(\V4/V2/A2/A2/c3 ),
    .ZN(\V4/V2/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A2/A2/M4/M2/_1_  (.A(\V4/V2/A2/A2/M4/s1 ),
    .B(\V4/V2/A2/A2/c3 ),
    .Z(\V4/V2/s2 [7]));
 OR2_X1 \V4/V2/A2/A2/M4/_0_  (.A1(\V4/V2/A2/A2/M4/c1 ),
    .A2(\V4/V2/A2/A2/M4/c2 ),
    .ZN(\V4/V2/c2 ));
 AND2_X1 \V4/V2/A3/A1/M1/M1/_0_  (.A1(\V4/V2/v4 [0]),
    .A2(\V4/V2/s2 [4]),
    .ZN(\V4/V2/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M1/M1/_1_  (.A(\V4/V2/v4 [0]),
    .B(\V4/V2/s2 [4]),
    .Z(\V4/V2/A3/A1/M1/s1 ));
 AND2_X1 \V4/V2/A3/A1/M1/M2/_0_  (.A1(\V4/V2/A3/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M1/M2/_1_  (.A(\V4/V2/A3/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/v2 [8]));
 OR2_X1 \V4/V2/A3/A1/M1/_0_  (.A1(\V4/V2/A3/A1/M1/c1 ),
    .A2(\V4/V2/A3/A1/M1/c2 ),
    .ZN(\V4/V2/A3/A1/c1 ));
 AND2_X1 \V4/V2/A3/A1/M2/M1/_0_  (.A1(\V4/V2/v4 [1]),
    .A2(\V4/V2/s2 [5]),
    .ZN(\V4/V2/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M2/M1/_1_  (.A(\V4/V2/v4 [1]),
    .B(\V4/V2/s2 [5]),
    .Z(\V4/V2/A3/A1/M2/s1 ));
 AND2_X1 \V4/V2/A3/A1/M2/M2/_0_  (.A1(\V4/V2/A3/A1/M2/s1 ),
    .A2(\V4/V2/A3/A1/c1 ),
    .ZN(\V4/V2/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M2/M2/_1_  (.A(\V4/V2/A3/A1/M2/s1 ),
    .B(\V4/V2/A3/A1/c1 ),
    .Z(\V4/v2 [9]));
 OR2_X1 \V4/V2/A3/A1/M2/_0_  (.A1(\V4/V2/A3/A1/M2/c1 ),
    .A2(\V4/V2/A3/A1/M2/c2 ),
    .ZN(\V4/V2/A3/A1/c2 ));
 AND2_X1 \V4/V2/A3/A1/M3/M1/_0_  (.A1(\V4/V2/v4 [2]),
    .A2(\V4/V2/s2 [6]),
    .ZN(\V4/V2/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M3/M1/_1_  (.A(\V4/V2/v4 [2]),
    .B(\V4/V2/s2 [6]),
    .Z(\V4/V2/A3/A1/M3/s1 ));
 AND2_X1 \V4/V2/A3/A1/M3/M2/_0_  (.A1(\V4/V2/A3/A1/M3/s1 ),
    .A2(\V4/V2/A3/A1/c2 ),
    .ZN(\V4/V2/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M3/M2/_1_  (.A(\V4/V2/A3/A1/M3/s1 ),
    .B(\V4/V2/A3/A1/c2 ),
    .Z(\V4/v2 [10]));
 OR2_X1 \V4/V2/A3/A1/M3/_0_  (.A1(\V4/V2/A3/A1/M3/c1 ),
    .A2(\V4/V2/A3/A1/M3/c2 ),
    .ZN(\V4/V2/A3/A1/c3 ));
 AND2_X1 \V4/V2/A3/A1/M4/M1/_0_  (.A1(\V4/V2/v4 [3]),
    .A2(\V4/V2/s2 [7]),
    .ZN(\V4/V2/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V2/A3/A1/M4/M1/_1_  (.A(\V4/V2/v4 [3]),
    .B(\V4/V2/s2 [7]),
    .Z(\V4/V2/A3/A1/M4/s1 ));
 AND2_X1 \V4/V2/A3/A1/M4/M2/_0_  (.A1(\V4/V2/A3/A1/M4/s1 ),
    .A2(\V4/V2/A3/A1/c3 ),
    .ZN(\V4/V2/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V2/A3/A1/M4/M2/_1_  (.A(\V4/V2/A3/A1/M4/s1 ),
    .B(\V4/V2/A3/A1/c3 ),
    .Z(\V4/v2 [11]));
 OR2_X1 \V4/V2/A3/A1/M4/_0_  (.A1(\V4/V2/A3/A1/M4/c1 ),
    .A2(\V4/V2/A3/A1/M4/c2 ),
    .ZN(\V4/V2/A3/c1 ));
 AND2_X1 \V4/V2/A3/A2/M1/M1/_0_  (.A1(\V4/V2/v4 [4]),
    .A2(\V4/V2/c3 ),
    .ZN(\V4/V2/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M1/M1/_1_  (.A(\V4/V2/v4 [4]),
    .B(\V4/V2/c3 ),
    .Z(\V4/V2/A3/A2/M1/s1 ));
 AND2_X1 \V4/V2/A3/A2/M1/M2/_0_  (.A1(\V4/V2/A3/A2/M1/s1 ),
    .A2(\V4/V2/A3/c1 ),
    .ZN(\V4/V2/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M1/M2/_1_  (.A(\V4/V2/A3/A2/M1/s1 ),
    .B(\V4/V2/A3/c1 ),
    .Z(\V4/v2 [12]));
 OR2_X1 \V4/V2/A3/A2/M1/_0_  (.A1(\V4/V2/A3/A2/M1/c1 ),
    .A2(\V4/V2/A3/A2/M1/c2 ),
    .ZN(\V4/V2/A3/A2/c1 ));
 AND2_X1 \V4/V2/A3/A2/M2/M1/_0_  (.A1(\V4/V2/v4 [5]),
    .A2(net1),
    .ZN(\V4/V2/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M2/M1/_1_  (.A(\V4/V2/v4 [5]),
    .B(net1),
    .Z(\V4/V2/A3/A2/M2/s1 ));
 AND2_X1 \V4/V2/A3/A2/M2/M2/_0_  (.A1(\V4/V2/A3/A2/M2/s1 ),
    .A2(\V4/V2/A3/A2/c1 ),
    .ZN(\V4/V2/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M2/M2/_1_  (.A(\V4/V2/A3/A2/M2/s1 ),
    .B(\V4/V2/A3/A2/c1 ),
    .Z(\V4/v2 [13]));
 OR2_X1 \V4/V2/A3/A2/M2/_0_  (.A1(\V4/V2/A3/A2/M2/c1 ),
    .A2(\V4/V2/A3/A2/M2/c2 ),
    .ZN(\V4/V2/A3/A2/c2 ));
 AND2_X1 \V4/V2/A3/A2/M3/M1/_0_  (.A1(\V4/V2/v4 [6]),
    .A2(net1),
    .ZN(\V4/V2/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M3/M1/_1_  (.A(\V4/V2/v4 [6]),
    .B(net1),
    .Z(\V4/V2/A3/A2/M3/s1 ));
 AND2_X1 \V4/V2/A3/A2/M3/M2/_0_  (.A1(\V4/V2/A3/A2/M3/s1 ),
    .A2(\V4/V2/A3/A2/c2 ),
    .ZN(\V4/V2/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M3/M2/_1_  (.A(\V4/V2/A3/A2/M3/s1 ),
    .B(\V4/V2/A3/A2/c2 ),
    .Z(\V4/v2 [14]));
 OR2_X1 \V4/V2/A3/A2/M3/_0_  (.A1(\V4/V2/A3/A2/M3/c1 ),
    .A2(\V4/V2/A3/A2/M3/c2 ),
    .ZN(\V4/V2/A3/A2/c3 ));
 AND2_X1 \V4/V2/A3/A2/M4/M1/_0_  (.A1(\V4/V2/v4 [7]),
    .A2(net1),
    .ZN(\V4/V2/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V2/A3/A2/M4/M1/_1_  (.A(\V4/V2/v4 [7]),
    .B(net1),
    .Z(\V4/V2/A3/A2/M4/s1 ));
 AND2_X1 \V4/V2/A3/A2/M4/M2/_0_  (.A1(\V4/V2/A3/A2/M4/s1 ),
    .A2(\V4/V2/A3/A2/c3 ),
    .ZN(\V4/V2/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V2/A3/A2/M4/M2/_1_  (.A(\V4/V2/A3/A2/M4/s1 ),
    .B(\V4/V2/A3/A2/c3 ),
    .Z(\V4/v2 [15]));
 OR2_X1 \V4/V2/A3/A2/M4/_0_  (.A1(\V4/V2/A3/A2/M4/c1 ),
    .A2(\V4/V2/A3/A2/M4/c2 ),
    .ZN(\V4/V2/overflow ));
 AND2_X1 \V4/V2/V1/A1/M1/M1/_0_  (.A1(\V4/V2/V1/v2 [0]),
    .A2(\V4/V2/V1/v3 [0]),
    .ZN(\V4/V2/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M1/M1/_1_  (.A(\V4/V2/V1/v2 [0]),
    .B(\V4/V2/V1/v3 [0]),
    .Z(\V4/V2/V1/A1/M1/s1 ));
 AND2_X1 \V4/V2/V1/A1/M1/M2/_0_  (.A1(\V4/V2/V1/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M1/M2/_1_  (.A(\V4/V2/V1/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/V1/s1 [0]));
 OR2_X1 \V4/V2/V1/A1/M1/_0_  (.A1(\V4/V2/V1/A1/M1/c1 ),
    .A2(\V4/V2/V1/A1/M1/c2 ),
    .ZN(\V4/V2/V1/A1/c1 ));
 AND2_X1 \V4/V2/V1/A1/M2/M1/_0_  (.A1(\V4/V2/V1/v2 [1]),
    .A2(\V4/V2/V1/v3 [1]),
    .ZN(\V4/V2/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M2/M1/_1_  (.A(\V4/V2/V1/v2 [1]),
    .B(\V4/V2/V1/v3 [1]),
    .Z(\V4/V2/V1/A1/M2/s1 ));
 AND2_X1 \V4/V2/V1/A1/M2/M2/_0_  (.A1(\V4/V2/V1/A1/M2/s1 ),
    .A2(\V4/V2/V1/A1/c1 ),
    .ZN(\V4/V2/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M2/M2/_1_  (.A(\V4/V2/V1/A1/M2/s1 ),
    .B(\V4/V2/V1/A1/c1 ),
    .Z(\V4/V2/V1/s1 [1]));
 OR2_X1 \V4/V2/V1/A1/M2/_0_  (.A1(\V4/V2/V1/A1/M2/c1 ),
    .A2(\V4/V2/V1/A1/M2/c2 ),
    .ZN(\V4/V2/V1/A1/c2 ));
 AND2_X1 \V4/V2/V1/A1/M3/M1/_0_  (.A1(\V4/V2/V1/v2 [2]),
    .A2(\V4/V2/V1/v3 [2]),
    .ZN(\V4/V2/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M3/M1/_1_  (.A(\V4/V2/V1/v2 [2]),
    .B(\V4/V2/V1/v3 [2]),
    .Z(\V4/V2/V1/A1/M3/s1 ));
 AND2_X1 \V4/V2/V1/A1/M3/M2/_0_  (.A1(\V4/V2/V1/A1/M3/s1 ),
    .A2(\V4/V2/V1/A1/c2 ),
    .ZN(\V4/V2/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M3/M2/_1_  (.A(\V4/V2/V1/A1/M3/s1 ),
    .B(\V4/V2/V1/A1/c2 ),
    .Z(\V4/V2/V1/s1 [2]));
 OR2_X1 \V4/V2/V1/A1/M3/_0_  (.A1(\V4/V2/V1/A1/M3/c1 ),
    .A2(\V4/V2/V1/A1/M3/c2 ),
    .ZN(\V4/V2/V1/A1/c3 ));
 AND2_X1 \V4/V2/V1/A1/M4/M1/_0_  (.A1(\V4/V2/V1/v2 [3]),
    .A2(\V4/V2/V1/v3 [3]),
    .ZN(\V4/V2/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A1/M4/M1/_1_  (.A(\V4/V2/V1/v2 [3]),
    .B(\V4/V2/V1/v3 [3]),
    .Z(\V4/V2/V1/A1/M4/s1 ));
 AND2_X1 \V4/V2/V1/A1/M4/M2/_0_  (.A1(\V4/V2/V1/A1/M4/s1 ),
    .A2(\V4/V2/V1/A1/c3 ),
    .ZN(\V4/V2/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A1/M4/M2/_1_  (.A(\V4/V2/V1/A1/M4/s1 ),
    .B(\V4/V2/V1/A1/c3 ),
    .Z(\V4/V2/V1/s1 [3]));
 OR2_X1 \V4/V2/V1/A1/M4/_0_  (.A1(\V4/V2/V1/A1/M4/c1 ),
    .A2(\V4/V2/V1/A1/M4/c2 ),
    .ZN(\V4/V2/V1/c1 ));
 AND2_X1 \V4/V2/V1/A2/M1/M1/_0_  (.A1(\V4/V2/V1/s1 [0]),
    .A2(\V4/V2/V1/v1 [2]),
    .ZN(\V4/V2/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M1/M1/_1_  (.A(\V4/V2/V1/s1 [0]),
    .B(\V4/V2/V1/v1 [2]),
    .Z(\V4/V2/V1/A2/M1/s1 ));
 AND2_X1 \V4/V2/V1/A2/M1/M2/_0_  (.A1(\V4/V2/V1/A2/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M1/M2/_1_  (.A(\V4/V2/V1/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/v2 [2]));
 OR2_X1 \V4/V2/V1/A2/M1/_0_  (.A1(\V4/V2/V1/A2/M1/c1 ),
    .A2(\V4/V2/V1/A2/M1/c2 ),
    .ZN(\V4/V2/V1/A2/c1 ));
 AND2_X1 \V4/V2/V1/A2/M2/M1/_0_  (.A1(\V4/V2/V1/s1 [1]),
    .A2(\V4/V2/V1/v1 [3]),
    .ZN(\V4/V2/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M2/M1/_1_  (.A(\V4/V2/V1/s1 [1]),
    .B(\V4/V2/V1/v1 [3]),
    .Z(\V4/V2/V1/A2/M2/s1 ));
 AND2_X1 \V4/V2/V1/A2/M2/M2/_0_  (.A1(\V4/V2/V1/A2/M2/s1 ),
    .A2(\V4/V2/V1/A2/c1 ),
    .ZN(\V4/V2/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M2/M2/_1_  (.A(\V4/V2/V1/A2/M2/s1 ),
    .B(\V4/V2/V1/A2/c1 ),
    .Z(\V4/v2 [3]));
 OR2_X1 \V4/V2/V1/A2/M2/_0_  (.A1(\V4/V2/V1/A2/M2/c1 ),
    .A2(\V4/V2/V1/A2/M2/c2 ),
    .ZN(\V4/V2/V1/A2/c2 ));
 AND2_X1 \V4/V2/V1/A2/M3/M1/_0_  (.A1(\V4/V2/V1/s1 [2]),
    .A2(net1),
    .ZN(\V4/V2/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M3/M1/_1_  (.A(\V4/V2/V1/s1 [2]),
    .B(net1),
    .Z(\V4/V2/V1/A2/M3/s1 ));
 AND2_X1 \V4/V2/V1/A2/M3/M2/_0_  (.A1(\V4/V2/V1/A2/M3/s1 ),
    .A2(\V4/V2/V1/A2/c2 ),
    .ZN(\V4/V2/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M3/M2/_1_  (.A(\V4/V2/V1/A2/M3/s1 ),
    .B(\V4/V2/V1/A2/c2 ),
    .Z(\V4/V2/V1/s2 [2]));
 OR2_X1 \V4/V2/V1/A2/M3/_0_  (.A1(\V4/V2/V1/A2/M3/c1 ),
    .A2(\V4/V2/V1/A2/M3/c2 ),
    .ZN(\V4/V2/V1/A2/c3 ));
 AND2_X1 \V4/V2/V1/A2/M4/M1/_0_  (.A1(\V4/V2/V1/s1 [3]),
    .A2(net1),
    .ZN(\V4/V2/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A2/M4/M1/_1_  (.A(\V4/V2/V1/s1 [3]),
    .B(net1),
    .Z(\V4/V2/V1/A2/M4/s1 ));
 AND2_X1 \V4/V2/V1/A2/M4/M2/_0_  (.A1(\V4/V2/V1/A2/M4/s1 ),
    .A2(\V4/V2/V1/A2/c3 ),
    .ZN(\V4/V2/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A2/M4/M2/_1_  (.A(\V4/V2/V1/A2/M4/s1 ),
    .B(\V4/V2/V1/A2/c3 ),
    .Z(\V4/V2/V1/s2 [3]));
 OR2_X1 \V4/V2/V1/A2/M4/_0_  (.A1(\V4/V2/V1/A2/M4/c1 ),
    .A2(\V4/V2/V1/A2/M4/c2 ),
    .ZN(\V4/V2/V1/c2 ));
 AND2_X1 \V4/V2/V1/A3/M1/M1/_0_  (.A1(\V4/V2/V1/v4 [0]),
    .A2(\V4/V2/V1/s2 [2]),
    .ZN(\V4/V2/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M1/M1/_1_  (.A(\V4/V2/V1/v4 [0]),
    .B(\V4/V2/V1/s2 [2]),
    .Z(\V4/V2/V1/A3/M1/s1 ));
 AND2_X1 \V4/V2/V1/A3/M1/M2/_0_  (.A1(\V4/V2/V1/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M1/M2/_1_  (.A(\V4/V2/V1/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v1 [4]));
 OR2_X1 \V4/V2/V1/A3/M1/_0_  (.A1(\V4/V2/V1/A3/M1/c1 ),
    .A2(\V4/V2/V1/A3/M1/c2 ),
    .ZN(\V4/V2/V1/A3/c1 ));
 AND2_X1 \V4/V2/V1/A3/M2/M1/_0_  (.A1(\V4/V2/V1/v4 [1]),
    .A2(\V4/V2/V1/s2 [3]),
    .ZN(\V4/V2/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M2/M1/_1_  (.A(\V4/V2/V1/v4 [1]),
    .B(\V4/V2/V1/s2 [3]),
    .Z(\V4/V2/V1/A3/M2/s1 ));
 AND2_X1 \V4/V2/V1/A3/M2/M2/_0_  (.A1(\V4/V2/V1/A3/M2/s1 ),
    .A2(\V4/V2/V1/A3/c1 ),
    .ZN(\V4/V2/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M2/M2/_1_  (.A(\V4/V2/V1/A3/M2/s1 ),
    .B(\V4/V2/V1/A3/c1 ),
    .Z(\V4/V2/v1 [5]));
 OR2_X1 \V4/V2/V1/A3/M2/_0_  (.A1(\V4/V2/V1/A3/M2/c1 ),
    .A2(\V4/V2/V1/A3/M2/c2 ),
    .ZN(\V4/V2/V1/A3/c2 ));
 AND2_X1 \V4/V2/V1/A3/M3/M1/_0_  (.A1(\V4/V2/V1/v4 [2]),
    .A2(\V4/V2/V1/c3 ),
    .ZN(\V4/V2/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M3/M1/_1_  (.A(\V4/V2/V1/v4 [2]),
    .B(\V4/V2/V1/c3 ),
    .Z(\V4/V2/V1/A3/M3/s1 ));
 AND2_X1 \V4/V2/V1/A3/M3/M2/_0_  (.A1(\V4/V2/V1/A3/M3/s1 ),
    .A2(\V4/V2/V1/A3/c2 ),
    .ZN(\V4/V2/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M3/M2/_1_  (.A(\V4/V2/V1/A3/M3/s1 ),
    .B(\V4/V2/V1/A3/c2 ),
    .Z(\V4/V2/v1 [6]));
 OR2_X1 \V4/V2/V1/A3/M3/_0_  (.A1(\V4/V2/V1/A3/M3/c1 ),
    .A2(\V4/V2/V1/A3/M3/c2 ),
    .ZN(\V4/V2/V1/A3/c3 ));
 AND2_X1 \V4/V2/V1/A3/M4/M1/_0_  (.A1(\V4/V2/V1/v4 [3]),
    .A2(net1),
    .ZN(\V4/V2/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V1/A3/M4/M1/_1_  (.A(\V4/V2/V1/v4 [3]),
    .B(net1),
    .Z(\V4/V2/V1/A3/M4/s1 ));
 AND2_X1 \V4/V2/V1/A3/M4/M2/_0_  (.A1(\V4/V2/V1/A3/M4/s1 ),
    .A2(\V4/V2/V1/A3/c3 ),
    .ZN(\V4/V2/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V1/A3/M4/M2/_1_  (.A(\V4/V2/V1/A3/M4/s1 ),
    .B(\V4/V2/V1/A3/c3 ),
    .Z(\V4/V2/v1 [7]));
 OR2_X1 \V4/V2/V1/A3/M4/_0_  (.A1(\V4/V2/V1/A3/M4/c1 ),
    .A2(\V4/V2/V1/A3/M4/c2 ),
    .ZN(\V4/V2/V1/overflow ));
 AND2_X1 \V4/V2/V1/V1/HA1/_0_  (.A1(\V4/V2/V1/V1/w2 ),
    .A2(\V4/V2/V1/V1/w1 ),
    .ZN(\V4/V2/V1/V1/w4 ));
 XOR2_X2 \V4/V2/V1/V1/HA1/_1_  (.A(\V4/V2/V1/V1/w2 ),
    .B(\V4/V2/V1/V1/w1 ),
    .Z(\V4/v2 [1]));
 AND2_X1 \V4/V2/V1/V1/HA2/_0_  (.A1(\V4/V2/V1/V1/w4 ),
    .A2(\V4/V2/V1/V1/w3 ),
    .ZN(\V4/V2/V1/v1 [3]));
 XOR2_X2 \V4/V2/V1/V1/HA2/_1_  (.A(\V4/V2/V1/V1/w4 ),
    .B(\V4/V2/V1/V1/w3 ),
    .Z(\V4/V2/V1/v1 [2]));
 AND2_X1 \V4/V2/V1/V1/_0_  (.A1(net33),
    .A2(net22),
    .ZN(\V4/v2 [0]));
 AND2_X1 \V4/V2/V1/V1/_1_  (.A1(net33),
    .A2(net21),
    .ZN(\V4/V2/V1/V1/w1 ));
 AND2_X1 \V4/V2/V1/V1/_2_  (.A1(net22),
    .A2(net32),
    .ZN(\V4/V2/V1/V1/w2 ));
 AND2_X1 \V4/V2/V1/V1/_3_  (.A1(net21),
    .A2(net32),
    .ZN(\V4/V2/V1/V1/w3 ));
 AND2_X1 \V4/V2/V1/V2/HA1/_0_  (.A1(\V4/V2/V1/V2/w2 ),
    .A2(\V4/V2/V1/V2/w1 ),
    .ZN(\V4/V2/V1/V2/w4 ));
 XOR2_X2 \V4/V2/V1/V2/HA1/_1_  (.A(\V4/V2/V1/V2/w2 ),
    .B(\V4/V2/V1/V2/w1 ),
    .Z(\V4/V2/V1/v2 [1]));
 AND2_X1 \V4/V2/V1/V2/HA2/_0_  (.A1(\V4/V2/V1/V2/w4 ),
    .A2(\V4/V2/V1/V2/w3 ),
    .ZN(\V4/V2/V1/v2 [3]));
 XOR2_X2 \V4/V2/V1/V2/HA2/_1_  (.A(\V4/V2/V1/V2/w4 ),
    .B(\V4/V2/V1/V2/w3 ),
    .Z(\V4/V2/V1/v2 [2]));
 AND2_X1 \V4/V2/V1/V2/_0_  (.A1(net31),
    .A2(net22),
    .ZN(\V4/V2/V1/v2 [0]));
 AND2_X1 \V4/V2/V1/V2/_1_  (.A1(net31),
    .A2(net21),
    .ZN(\V4/V2/V1/V2/w1 ));
 AND2_X1 \V4/V2/V1/V2/_2_  (.A1(net22),
    .A2(net30),
    .ZN(\V4/V2/V1/V2/w2 ));
 AND2_X1 \V4/V2/V1/V2/_3_  (.A1(net21),
    .A2(net30),
    .ZN(\V4/V2/V1/V2/w3 ));
 AND2_X1 \V4/V2/V1/V3/HA1/_0_  (.A1(\V4/V2/V1/V3/w2 ),
    .A2(\V4/V2/V1/V3/w1 ),
    .ZN(\V4/V2/V1/V3/w4 ));
 XOR2_X2 \V4/V2/V1/V3/HA1/_1_  (.A(\V4/V2/V1/V3/w2 ),
    .B(\V4/V2/V1/V3/w1 ),
    .Z(\V4/V2/V1/v3 [1]));
 AND2_X1 \V4/V2/V1/V3/HA2/_0_  (.A1(\V4/V2/V1/V3/w4 ),
    .A2(\V4/V2/V1/V3/w3 ),
    .ZN(\V4/V2/V1/v3 [3]));
 XOR2_X2 \V4/V2/V1/V3/HA2/_1_  (.A(\V4/V2/V1/V3/w4 ),
    .B(\V4/V2/V1/V3/w3 ),
    .Z(\V4/V2/V1/v3 [2]));
 AND2_X1 \V4/V2/V1/V3/_0_  (.A1(net33),
    .A2(B[18]),
    .ZN(\V4/V2/V1/v3 [0]));
 AND2_X1 \V4/V2/V1/V3/_1_  (.A1(net33),
    .A2(B[19]),
    .ZN(\V4/V2/V1/V3/w1 ));
 AND2_X1 \V4/V2/V1/V3/_2_  (.A1(B[18]),
    .A2(net32),
    .ZN(\V4/V2/V1/V3/w2 ));
 AND2_X1 \V4/V2/V1/V3/_3_  (.A1(B[19]),
    .A2(net32),
    .ZN(\V4/V2/V1/V3/w3 ));
 AND2_X1 \V4/V2/V1/V4/HA1/_0_  (.A1(\V4/V2/V1/V4/w2 ),
    .A2(\V4/V2/V1/V4/w1 ),
    .ZN(\V4/V2/V1/V4/w4 ));
 XOR2_X2 \V4/V2/V1/V4/HA1/_1_  (.A(\V4/V2/V1/V4/w2 ),
    .B(\V4/V2/V1/V4/w1 ),
    .Z(\V4/V2/V1/v4 [1]));
 AND2_X1 \V4/V2/V1/V4/HA2/_0_  (.A1(\V4/V2/V1/V4/w4 ),
    .A2(\V4/V2/V1/V4/w3 ),
    .ZN(\V4/V2/V1/v4 [3]));
 XOR2_X2 \V4/V2/V1/V4/HA2/_1_  (.A(\V4/V2/V1/V4/w4 ),
    .B(\V4/V2/V1/V4/w3 ),
    .Z(\V4/V2/V1/v4 [2]));
 AND2_X1 \V4/V2/V1/V4/_0_  (.A1(net31),
    .A2(B[18]),
    .ZN(\V4/V2/V1/v4 [0]));
 AND2_X1 \V4/V2/V1/V4/_1_  (.A1(net31),
    .A2(B[19]),
    .ZN(\V4/V2/V1/V4/w1 ));
 AND2_X1 \V4/V2/V1/V4/_2_  (.A1(B[18]),
    .A2(net30),
    .ZN(\V4/V2/V1/V4/w2 ));
 AND2_X1 \V4/V2/V1/V4/_3_  (.A1(B[19]),
    .A2(net30),
    .ZN(\V4/V2/V1/V4/w3 ));
 OR2_X1 \V4/V2/V1/_0_  (.A1(\V4/V2/V1/c1 ),
    .A2(\V4/V2/V1/c2 ),
    .ZN(\V4/V2/V1/c3 ));
 AND2_X1 \V4/V2/V2/A1/M1/M1/_0_  (.A1(\V4/V2/V2/v2 [0]),
    .A2(\V4/V2/V2/v3 [0]),
    .ZN(\V4/V2/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M1/M1/_1_  (.A(\V4/V2/V2/v2 [0]),
    .B(\V4/V2/V2/v3 [0]),
    .Z(\V4/V2/V2/A1/M1/s1 ));
 AND2_X1 \V4/V2/V2/A1/M1/M2/_0_  (.A1(\V4/V2/V2/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M1/M2/_1_  (.A(\V4/V2/V2/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/V2/s1 [0]));
 OR2_X1 \V4/V2/V2/A1/M1/_0_  (.A1(\V4/V2/V2/A1/M1/c1 ),
    .A2(\V4/V2/V2/A1/M1/c2 ),
    .ZN(\V4/V2/V2/A1/c1 ));
 AND2_X1 \V4/V2/V2/A1/M2/M1/_0_  (.A1(\V4/V2/V2/v2 [1]),
    .A2(\V4/V2/V2/v3 [1]),
    .ZN(\V4/V2/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M2/M1/_1_  (.A(\V4/V2/V2/v2 [1]),
    .B(\V4/V2/V2/v3 [1]),
    .Z(\V4/V2/V2/A1/M2/s1 ));
 AND2_X1 \V4/V2/V2/A1/M2/M2/_0_  (.A1(\V4/V2/V2/A1/M2/s1 ),
    .A2(\V4/V2/V2/A1/c1 ),
    .ZN(\V4/V2/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M2/M2/_1_  (.A(\V4/V2/V2/A1/M2/s1 ),
    .B(\V4/V2/V2/A1/c1 ),
    .Z(\V4/V2/V2/s1 [1]));
 OR2_X1 \V4/V2/V2/A1/M2/_0_  (.A1(\V4/V2/V2/A1/M2/c1 ),
    .A2(\V4/V2/V2/A1/M2/c2 ),
    .ZN(\V4/V2/V2/A1/c2 ));
 AND2_X1 \V4/V2/V2/A1/M3/M1/_0_  (.A1(\V4/V2/V2/v2 [2]),
    .A2(\V4/V2/V2/v3 [2]),
    .ZN(\V4/V2/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M3/M1/_1_  (.A(\V4/V2/V2/v2 [2]),
    .B(\V4/V2/V2/v3 [2]),
    .Z(\V4/V2/V2/A1/M3/s1 ));
 AND2_X1 \V4/V2/V2/A1/M3/M2/_0_  (.A1(\V4/V2/V2/A1/M3/s1 ),
    .A2(\V4/V2/V2/A1/c2 ),
    .ZN(\V4/V2/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M3/M2/_1_  (.A(\V4/V2/V2/A1/M3/s1 ),
    .B(\V4/V2/V2/A1/c2 ),
    .Z(\V4/V2/V2/s1 [2]));
 OR2_X1 \V4/V2/V2/A1/M3/_0_  (.A1(\V4/V2/V2/A1/M3/c1 ),
    .A2(\V4/V2/V2/A1/M3/c2 ),
    .ZN(\V4/V2/V2/A1/c3 ));
 AND2_X1 \V4/V2/V2/A1/M4/M1/_0_  (.A1(\V4/V2/V2/v2 [3]),
    .A2(\V4/V2/V2/v3 [3]),
    .ZN(\V4/V2/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A1/M4/M1/_1_  (.A(\V4/V2/V2/v2 [3]),
    .B(\V4/V2/V2/v3 [3]),
    .Z(\V4/V2/V2/A1/M4/s1 ));
 AND2_X1 \V4/V2/V2/A1/M4/M2/_0_  (.A1(\V4/V2/V2/A1/M4/s1 ),
    .A2(\V4/V2/V2/A1/c3 ),
    .ZN(\V4/V2/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A1/M4/M2/_1_  (.A(\V4/V2/V2/A1/M4/s1 ),
    .B(\V4/V2/V2/A1/c3 ),
    .Z(\V4/V2/V2/s1 [3]));
 OR2_X1 \V4/V2/V2/A1/M4/_0_  (.A1(\V4/V2/V2/A1/M4/c1 ),
    .A2(\V4/V2/V2/A1/M4/c2 ),
    .ZN(\V4/V2/V2/c1 ));
 AND2_X1 \V4/V2/V2/A2/M1/M1/_0_  (.A1(\V4/V2/V2/s1 [0]),
    .A2(\V4/V2/V2/v1 [2]),
    .ZN(\V4/V2/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M1/M1/_1_  (.A(\V4/V2/V2/s1 [0]),
    .B(\V4/V2/V2/v1 [2]),
    .Z(\V4/V2/V2/A2/M1/s1 ));
 AND2_X1 \V4/V2/V2/A2/M1/M2/_0_  (.A1(\V4/V2/V2/A2/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M1/M2/_1_  (.A(\V4/V2/V2/A2/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v2 [2]));
 OR2_X1 \V4/V2/V2/A2/M1/_0_  (.A1(\V4/V2/V2/A2/M1/c1 ),
    .A2(\V4/V2/V2/A2/M1/c2 ),
    .ZN(\V4/V2/V2/A2/c1 ));
 AND2_X1 \V4/V2/V2/A2/M2/M1/_0_  (.A1(\V4/V2/V2/s1 [1]),
    .A2(\V4/V2/V2/v1 [3]),
    .ZN(\V4/V2/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M2/M1/_1_  (.A(\V4/V2/V2/s1 [1]),
    .B(\V4/V2/V2/v1 [3]),
    .Z(\V4/V2/V2/A2/M2/s1 ));
 AND2_X1 \V4/V2/V2/A2/M2/M2/_0_  (.A1(\V4/V2/V2/A2/M2/s1 ),
    .A2(\V4/V2/V2/A2/c1 ),
    .ZN(\V4/V2/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M2/M2/_1_  (.A(\V4/V2/V2/A2/M2/s1 ),
    .B(\V4/V2/V2/A2/c1 ),
    .Z(\V4/V2/v2 [3]));
 OR2_X1 \V4/V2/V2/A2/M2/_0_  (.A1(\V4/V2/V2/A2/M2/c1 ),
    .A2(\V4/V2/V2/A2/M2/c2 ),
    .ZN(\V4/V2/V2/A2/c2 ));
 AND2_X1 \V4/V2/V2/A2/M3/M1/_0_  (.A1(\V4/V2/V2/s1 [2]),
    .A2(net1),
    .ZN(\V4/V2/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M3/M1/_1_  (.A(\V4/V2/V2/s1 [2]),
    .B(net1),
    .Z(\V4/V2/V2/A2/M3/s1 ));
 AND2_X1 \V4/V2/V2/A2/M3/M2/_0_  (.A1(\V4/V2/V2/A2/M3/s1 ),
    .A2(\V4/V2/V2/A2/c2 ),
    .ZN(\V4/V2/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M3/M2/_1_  (.A(\V4/V2/V2/A2/M3/s1 ),
    .B(\V4/V2/V2/A2/c2 ),
    .Z(\V4/V2/V2/s2 [2]));
 OR2_X1 \V4/V2/V2/A2/M3/_0_  (.A1(\V4/V2/V2/A2/M3/c1 ),
    .A2(\V4/V2/V2/A2/M3/c2 ),
    .ZN(\V4/V2/V2/A2/c3 ));
 AND2_X1 \V4/V2/V2/A2/M4/M1/_0_  (.A1(\V4/V2/V2/s1 [3]),
    .A2(net1),
    .ZN(\V4/V2/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A2/M4/M1/_1_  (.A(\V4/V2/V2/s1 [3]),
    .B(net1),
    .Z(\V4/V2/V2/A2/M4/s1 ));
 AND2_X1 \V4/V2/V2/A2/M4/M2/_0_  (.A1(\V4/V2/V2/A2/M4/s1 ),
    .A2(\V4/V2/V2/A2/c3 ),
    .ZN(\V4/V2/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A2/M4/M2/_1_  (.A(\V4/V2/V2/A2/M4/s1 ),
    .B(\V4/V2/V2/A2/c3 ),
    .Z(\V4/V2/V2/s2 [3]));
 OR2_X1 \V4/V2/V2/A2/M4/_0_  (.A1(\V4/V2/V2/A2/M4/c1 ),
    .A2(\V4/V2/V2/A2/M4/c2 ),
    .ZN(\V4/V2/V2/c2 ));
 AND2_X1 \V4/V2/V2/A3/M1/M1/_0_  (.A1(\V4/V2/V2/v4 [0]),
    .A2(\V4/V2/V2/s2 [2]),
    .ZN(\V4/V2/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M1/M1/_1_  (.A(\V4/V2/V2/v4 [0]),
    .B(\V4/V2/V2/s2 [2]),
    .Z(\V4/V2/V2/A3/M1/s1 ));
 AND2_X1 \V4/V2/V2/A3/M1/M2/_0_  (.A1(\V4/V2/V2/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M1/M2/_1_  (.A(\V4/V2/V2/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v2 [4]));
 OR2_X1 \V4/V2/V2/A3/M1/_0_  (.A1(\V4/V2/V2/A3/M1/c1 ),
    .A2(\V4/V2/V2/A3/M1/c2 ),
    .ZN(\V4/V2/V2/A3/c1 ));
 AND2_X1 \V4/V2/V2/A3/M2/M1/_0_  (.A1(\V4/V2/V2/v4 [1]),
    .A2(\V4/V2/V2/s2 [3]),
    .ZN(\V4/V2/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M2/M1/_1_  (.A(\V4/V2/V2/v4 [1]),
    .B(\V4/V2/V2/s2 [3]),
    .Z(\V4/V2/V2/A3/M2/s1 ));
 AND2_X1 \V4/V2/V2/A3/M2/M2/_0_  (.A1(\V4/V2/V2/A3/M2/s1 ),
    .A2(\V4/V2/V2/A3/c1 ),
    .ZN(\V4/V2/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M2/M2/_1_  (.A(\V4/V2/V2/A3/M2/s1 ),
    .B(\V4/V2/V2/A3/c1 ),
    .Z(\V4/V2/v2 [5]));
 OR2_X1 \V4/V2/V2/A3/M2/_0_  (.A1(\V4/V2/V2/A3/M2/c1 ),
    .A2(\V4/V2/V2/A3/M2/c2 ),
    .ZN(\V4/V2/V2/A3/c2 ));
 AND2_X1 \V4/V2/V2/A3/M3/M1/_0_  (.A1(\V4/V2/V2/v4 [2]),
    .A2(\V4/V2/V2/c3 ),
    .ZN(\V4/V2/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M3/M1/_1_  (.A(\V4/V2/V2/v4 [2]),
    .B(\V4/V2/V2/c3 ),
    .Z(\V4/V2/V2/A3/M3/s1 ));
 AND2_X1 \V4/V2/V2/A3/M3/M2/_0_  (.A1(\V4/V2/V2/A3/M3/s1 ),
    .A2(\V4/V2/V2/A3/c2 ),
    .ZN(\V4/V2/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M3/M2/_1_  (.A(\V4/V2/V2/A3/M3/s1 ),
    .B(\V4/V2/V2/A3/c2 ),
    .Z(\V4/V2/v2 [6]));
 OR2_X1 \V4/V2/V2/A3/M3/_0_  (.A1(\V4/V2/V2/A3/M3/c1 ),
    .A2(\V4/V2/V2/A3/M3/c2 ),
    .ZN(\V4/V2/V2/A3/c3 ));
 AND2_X1 \V4/V2/V2/A3/M4/M1/_0_  (.A1(\V4/V2/V2/v4 [3]),
    .A2(net1),
    .ZN(\V4/V2/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V2/A3/M4/M1/_1_  (.A(\V4/V2/V2/v4 [3]),
    .B(net1),
    .Z(\V4/V2/V2/A3/M4/s1 ));
 AND2_X1 \V4/V2/V2/A3/M4/M2/_0_  (.A1(\V4/V2/V2/A3/M4/s1 ),
    .A2(\V4/V2/V2/A3/c3 ),
    .ZN(\V4/V2/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V2/A3/M4/M2/_1_  (.A(\V4/V2/V2/A3/M4/s1 ),
    .B(\V4/V2/V2/A3/c3 ),
    .Z(\V4/V2/v2 [7]));
 OR2_X1 \V4/V2/V2/A3/M4/_0_  (.A1(\V4/V2/V2/A3/M4/c1 ),
    .A2(\V4/V2/V2/A3/M4/c2 ),
    .ZN(\V4/V2/V2/overflow ));
 AND2_X1 \V4/V2/V2/V1/HA1/_0_  (.A1(\V4/V2/V2/V1/w2 ),
    .A2(\V4/V2/V2/V1/w1 ),
    .ZN(\V4/V2/V2/V1/w4 ));
 XOR2_X2 \V4/V2/V2/V1/HA1/_1_  (.A(\V4/V2/V2/V1/w2 ),
    .B(\V4/V2/V2/V1/w1 ),
    .Z(\V4/V2/v2 [1]));
 AND2_X1 \V4/V2/V2/V1/HA2/_0_  (.A1(\V4/V2/V2/V1/w4 ),
    .A2(\V4/V2/V2/V1/w3 ),
    .ZN(\V4/V2/V2/v1 [3]));
 XOR2_X2 \V4/V2/V2/V1/HA2/_1_  (.A(\V4/V2/V2/V1/w4 ),
    .B(\V4/V2/V2/V1/w3 ),
    .Z(\V4/V2/V2/v1 [2]));
 AND2_X1 \V4/V2/V2/V1/_0_  (.A1(net29),
    .A2(net22),
    .ZN(\V4/V2/v2 [0]));
 AND2_X1 \V4/V2/V2/V1/_1_  (.A1(net29),
    .A2(net21),
    .ZN(\V4/V2/V2/V1/w1 ));
 AND2_X1 \V4/V2/V2/V1/_2_  (.A1(net22),
    .A2(net28),
    .ZN(\V4/V2/V2/V1/w2 ));
 AND2_X1 \V4/V2/V2/V1/_3_  (.A1(net21),
    .A2(net28),
    .ZN(\V4/V2/V2/V1/w3 ));
 AND2_X1 \V4/V2/V2/V2/HA1/_0_  (.A1(\V4/V2/V2/V2/w2 ),
    .A2(\V4/V2/V2/V2/w1 ),
    .ZN(\V4/V2/V2/V2/w4 ));
 XOR2_X2 \V4/V2/V2/V2/HA1/_1_  (.A(\V4/V2/V2/V2/w2 ),
    .B(\V4/V2/V2/V2/w1 ),
    .Z(\V4/V2/V2/v2 [1]));
 AND2_X1 \V4/V2/V2/V2/HA2/_0_  (.A1(\V4/V2/V2/V2/w4 ),
    .A2(\V4/V2/V2/V2/w3 ),
    .ZN(\V4/V2/V2/v2 [3]));
 XOR2_X2 \V4/V2/V2/V2/HA2/_1_  (.A(\V4/V2/V2/V2/w4 ),
    .B(\V4/V2/V2/V2/w3 ),
    .Z(\V4/V2/V2/v2 [2]));
 AND2_X1 \V4/V2/V2/V2/_0_  (.A1(net27),
    .A2(net22),
    .ZN(\V4/V2/V2/v2 [0]));
 AND2_X1 \V4/V2/V2/V2/_1_  (.A1(net27),
    .A2(net21),
    .ZN(\V4/V2/V2/V2/w1 ));
 AND2_X1 \V4/V2/V2/V2/_2_  (.A1(net22),
    .A2(net26),
    .ZN(\V4/V2/V2/V2/w2 ));
 AND2_X1 \V4/V2/V2/V2/_3_  (.A1(net21),
    .A2(net26),
    .ZN(\V4/V2/V2/V2/w3 ));
 AND2_X1 \V4/V2/V2/V3/HA1/_0_  (.A1(\V4/V2/V2/V3/w2 ),
    .A2(\V4/V2/V2/V3/w1 ),
    .ZN(\V4/V2/V2/V3/w4 ));
 XOR2_X2 \V4/V2/V2/V3/HA1/_1_  (.A(\V4/V2/V2/V3/w2 ),
    .B(\V4/V2/V2/V3/w1 ),
    .Z(\V4/V2/V2/v3 [1]));
 AND2_X1 \V4/V2/V2/V3/HA2/_0_  (.A1(\V4/V2/V2/V3/w4 ),
    .A2(\V4/V2/V2/V3/w3 ),
    .ZN(\V4/V2/V2/v3 [3]));
 XOR2_X2 \V4/V2/V2/V3/HA2/_1_  (.A(\V4/V2/V2/V3/w4 ),
    .B(\V4/V2/V2/V3/w3 ),
    .Z(\V4/V2/V2/v3 [2]));
 AND2_X1 \V4/V2/V2/V3/_0_  (.A1(net29),
    .A2(B[18]),
    .ZN(\V4/V2/V2/v3 [0]));
 AND2_X1 \V4/V2/V2/V3/_1_  (.A1(net29),
    .A2(B[19]),
    .ZN(\V4/V2/V2/V3/w1 ));
 AND2_X1 \V4/V2/V2/V3/_2_  (.A1(B[18]),
    .A2(net28),
    .ZN(\V4/V2/V2/V3/w2 ));
 AND2_X1 \V4/V2/V2/V3/_3_  (.A1(B[19]),
    .A2(net28),
    .ZN(\V4/V2/V2/V3/w3 ));
 AND2_X1 \V4/V2/V2/V4/HA1/_0_  (.A1(\V4/V2/V2/V4/w2 ),
    .A2(\V4/V2/V2/V4/w1 ),
    .ZN(\V4/V2/V2/V4/w4 ));
 XOR2_X2 \V4/V2/V2/V4/HA1/_1_  (.A(\V4/V2/V2/V4/w2 ),
    .B(\V4/V2/V2/V4/w1 ),
    .Z(\V4/V2/V2/v4 [1]));
 AND2_X1 \V4/V2/V2/V4/HA2/_0_  (.A1(\V4/V2/V2/V4/w4 ),
    .A2(\V4/V2/V2/V4/w3 ),
    .ZN(\V4/V2/V2/v4 [3]));
 XOR2_X2 \V4/V2/V2/V4/HA2/_1_  (.A(\V4/V2/V2/V4/w4 ),
    .B(\V4/V2/V2/V4/w3 ),
    .Z(\V4/V2/V2/v4 [2]));
 AND2_X1 \V4/V2/V2/V4/_0_  (.A1(net27),
    .A2(B[18]),
    .ZN(\V4/V2/V2/v4 [0]));
 AND2_X1 \V4/V2/V2/V4/_1_  (.A1(net27),
    .A2(B[19]),
    .ZN(\V4/V2/V2/V4/w1 ));
 AND2_X1 \V4/V2/V2/V4/_2_  (.A1(B[18]),
    .A2(net26),
    .ZN(\V4/V2/V2/V4/w2 ));
 AND2_X1 \V4/V2/V2/V4/_3_  (.A1(B[19]),
    .A2(net26),
    .ZN(\V4/V2/V2/V4/w3 ));
 OR2_X1 \V4/V2/V2/_0_  (.A1(\V4/V2/V2/c1 ),
    .A2(\V4/V2/V2/c2 ),
    .ZN(\V4/V2/V2/c3 ));
 AND2_X1 \V4/V2/V3/A1/M1/M1/_0_  (.A1(\V4/V2/V3/v2 [0]),
    .A2(\V4/V2/V3/v3 [0]),
    .ZN(\V4/V2/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M1/M1/_1_  (.A(\V4/V2/V3/v2 [0]),
    .B(\V4/V2/V3/v3 [0]),
    .Z(\V4/V2/V3/A1/M1/s1 ));
 AND2_X1 \V4/V2/V3/A1/M1/M2/_0_  (.A1(\V4/V2/V3/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M1/M2/_1_  (.A(\V4/V2/V3/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/V3/s1 [0]));
 OR2_X1 \V4/V2/V3/A1/M1/_0_  (.A1(\V4/V2/V3/A1/M1/c1 ),
    .A2(\V4/V2/V3/A1/M1/c2 ),
    .ZN(\V4/V2/V3/A1/c1 ));
 AND2_X1 \V4/V2/V3/A1/M2/M1/_0_  (.A1(\V4/V2/V3/v2 [1]),
    .A2(\V4/V2/V3/v3 [1]),
    .ZN(\V4/V2/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M2/M1/_1_  (.A(\V4/V2/V3/v2 [1]),
    .B(\V4/V2/V3/v3 [1]),
    .Z(\V4/V2/V3/A1/M2/s1 ));
 AND2_X1 \V4/V2/V3/A1/M2/M2/_0_  (.A1(\V4/V2/V3/A1/M2/s1 ),
    .A2(\V4/V2/V3/A1/c1 ),
    .ZN(\V4/V2/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M2/M2/_1_  (.A(\V4/V2/V3/A1/M2/s1 ),
    .B(\V4/V2/V3/A1/c1 ),
    .Z(\V4/V2/V3/s1 [1]));
 OR2_X1 \V4/V2/V3/A1/M2/_0_  (.A1(\V4/V2/V3/A1/M2/c1 ),
    .A2(\V4/V2/V3/A1/M2/c2 ),
    .ZN(\V4/V2/V3/A1/c2 ));
 AND2_X1 \V4/V2/V3/A1/M3/M1/_0_  (.A1(\V4/V2/V3/v2 [2]),
    .A2(\V4/V2/V3/v3 [2]),
    .ZN(\V4/V2/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M3/M1/_1_  (.A(\V4/V2/V3/v2 [2]),
    .B(\V4/V2/V3/v3 [2]),
    .Z(\V4/V2/V3/A1/M3/s1 ));
 AND2_X1 \V4/V2/V3/A1/M3/M2/_0_  (.A1(\V4/V2/V3/A1/M3/s1 ),
    .A2(\V4/V2/V3/A1/c2 ),
    .ZN(\V4/V2/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M3/M2/_1_  (.A(\V4/V2/V3/A1/M3/s1 ),
    .B(\V4/V2/V3/A1/c2 ),
    .Z(\V4/V2/V3/s1 [2]));
 OR2_X1 \V4/V2/V3/A1/M3/_0_  (.A1(\V4/V2/V3/A1/M3/c1 ),
    .A2(\V4/V2/V3/A1/M3/c2 ),
    .ZN(\V4/V2/V3/A1/c3 ));
 AND2_X1 \V4/V2/V3/A1/M4/M1/_0_  (.A1(\V4/V2/V3/v2 [3]),
    .A2(\V4/V2/V3/v3 [3]),
    .ZN(\V4/V2/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A1/M4/M1/_1_  (.A(\V4/V2/V3/v2 [3]),
    .B(\V4/V2/V3/v3 [3]),
    .Z(\V4/V2/V3/A1/M4/s1 ));
 AND2_X1 \V4/V2/V3/A1/M4/M2/_0_  (.A1(\V4/V2/V3/A1/M4/s1 ),
    .A2(\V4/V2/V3/A1/c3 ),
    .ZN(\V4/V2/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A1/M4/M2/_1_  (.A(\V4/V2/V3/A1/M4/s1 ),
    .B(\V4/V2/V3/A1/c3 ),
    .Z(\V4/V2/V3/s1 [3]));
 OR2_X1 \V4/V2/V3/A1/M4/_0_  (.A1(\V4/V2/V3/A1/M4/c1 ),
    .A2(\V4/V2/V3/A1/M4/c2 ),
    .ZN(\V4/V2/V3/c1 ));
 AND2_X1 \V4/V2/V3/A2/M1/M1/_0_  (.A1(\V4/V2/V3/s1 [0]),
    .A2(\V4/V2/V3/v1 [2]),
    .ZN(\V4/V2/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M1/M1/_1_  (.A(\V4/V2/V3/s1 [0]),
    .B(\V4/V2/V3/v1 [2]),
    .Z(\V4/V2/V3/A2/M1/s1 ));
 AND2_X1 \V4/V2/V3/A2/M1/M2/_0_  (.A1(\V4/V2/V3/A2/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M1/M2/_1_  (.A(\V4/V2/V3/A2/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v3 [2]));
 OR2_X1 \V4/V2/V3/A2/M1/_0_  (.A1(\V4/V2/V3/A2/M1/c1 ),
    .A2(\V4/V2/V3/A2/M1/c2 ),
    .ZN(\V4/V2/V3/A2/c1 ));
 AND2_X1 \V4/V2/V3/A2/M2/M1/_0_  (.A1(\V4/V2/V3/s1 [1]),
    .A2(\V4/V2/V3/v1 [3]),
    .ZN(\V4/V2/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M2/M1/_1_  (.A(\V4/V2/V3/s1 [1]),
    .B(\V4/V2/V3/v1 [3]),
    .Z(\V4/V2/V3/A2/M2/s1 ));
 AND2_X1 \V4/V2/V3/A2/M2/M2/_0_  (.A1(\V4/V2/V3/A2/M2/s1 ),
    .A2(\V4/V2/V3/A2/c1 ),
    .ZN(\V4/V2/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M2/M2/_1_  (.A(\V4/V2/V3/A2/M2/s1 ),
    .B(\V4/V2/V3/A2/c1 ),
    .Z(\V4/V2/v3 [3]));
 OR2_X1 \V4/V2/V3/A2/M2/_0_  (.A1(\V4/V2/V3/A2/M2/c1 ),
    .A2(\V4/V2/V3/A2/M2/c2 ),
    .ZN(\V4/V2/V3/A2/c2 ));
 AND2_X1 \V4/V2/V3/A2/M3/M1/_0_  (.A1(\V4/V2/V3/s1 [2]),
    .A2(net1),
    .ZN(\V4/V2/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M3/M1/_1_  (.A(\V4/V2/V3/s1 [2]),
    .B(net1),
    .Z(\V4/V2/V3/A2/M3/s1 ));
 AND2_X1 \V4/V2/V3/A2/M3/M2/_0_  (.A1(\V4/V2/V3/A2/M3/s1 ),
    .A2(\V4/V2/V3/A2/c2 ),
    .ZN(\V4/V2/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M3/M2/_1_  (.A(\V4/V2/V3/A2/M3/s1 ),
    .B(\V4/V2/V3/A2/c2 ),
    .Z(\V4/V2/V3/s2 [2]));
 OR2_X1 \V4/V2/V3/A2/M3/_0_  (.A1(\V4/V2/V3/A2/M3/c1 ),
    .A2(\V4/V2/V3/A2/M3/c2 ),
    .ZN(\V4/V2/V3/A2/c3 ));
 AND2_X1 \V4/V2/V3/A2/M4/M1/_0_  (.A1(\V4/V2/V3/s1 [3]),
    .A2(net1),
    .ZN(\V4/V2/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A2/M4/M1/_1_  (.A(\V4/V2/V3/s1 [3]),
    .B(net1),
    .Z(\V4/V2/V3/A2/M4/s1 ));
 AND2_X1 \V4/V2/V3/A2/M4/M2/_0_  (.A1(\V4/V2/V3/A2/M4/s1 ),
    .A2(\V4/V2/V3/A2/c3 ),
    .ZN(\V4/V2/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A2/M4/M2/_1_  (.A(\V4/V2/V3/A2/M4/s1 ),
    .B(\V4/V2/V3/A2/c3 ),
    .Z(\V4/V2/V3/s2 [3]));
 OR2_X1 \V4/V2/V3/A2/M4/_0_  (.A1(\V4/V2/V3/A2/M4/c1 ),
    .A2(\V4/V2/V3/A2/M4/c2 ),
    .ZN(\V4/V2/V3/c2 ));
 AND2_X1 \V4/V2/V3/A3/M1/M1/_0_  (.A1(\V4/V2/V3/v4 [0]),
    .A2(\V4/V2/V3/s2 [2]),
    .ZN(\V4/V2/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M1/M1/_1_  (.A(\V4/V2/V3/v4 [0]),
    .B(\V4/V2/V3/s2 [2]),
    .Z(\V4/V2/V3/A3/M1/s1 ));
 AND2_X1 \V4/V2/V3/A3/M1/M2/_0_  (.A1(\V4/V2/V3/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M1/M2/_1_  (.A(\V4/V2/V3/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v3 [4]));
 OR2_X1 \V4/V2/V3/A3/M1/_0_  (.A1(\V4/V2/V3/A3/M1/c1 ),
    .A2(\V4/V2/V3/A3/M1/c2 ),
    .ZN(\V4/V2/V3/A3/c1 ));
 AND2_X1 \V4/V2/V3/A3/M2/M1/_0_  (.A1(\V4/V2/V3/v4 [1]),
    .A2(\V4/V2/V3/s2 [3]),
    .ZN(\V4/V2/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M2/M1/_1_  (.A(\V4/V2/V3/v4 [1]),
    .B(\V4/V2/V3/s2 [3]),
    .Z(\V4/V2/V3/A3/M2/s1 ));
 AND2_X1 \V4/V2/V3/A3/M2/M2/_0_  (.A1(\V4/V2/V3/A3/M2/s1 ),
    .A2(\V4/V2/V3/A3/c1 ),
    .ZN(\V4/V2/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M2/M2/_1_  (.A(\V4/V2/V3/A3/M2/s1 ),
    .B(\V4/V2/V3/A3/c1 ),
    .Z(\V4/V2/v3 [5]));
 OR2_X1 \V4/V2/V3/A3/M2/_0_  (.A1(\V4/V2/V3/A3/M2/c1 ),
    .A2(\V4/V2/V3/A3/M2/c2 ),
    .ZN(\V4/V2/V3/A3/c2 ));
 AND2_X1 \V4/V2/V3/A3/M3/M1/_0_  (.A1(\V4/V2/V3/v4 [2]),
    .A2(\V4/V2/V3/c3 ),
    .ZN(\V4/V2/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M3/M1/_1_  (.A(\V4/V2/V3/v4 [2]),
    .B(\V4/V2/V3/c3 ),
    .Z(\V4/V2/V3/A3/M3/s1 ));
 AND2_X1 \V4/V2/V3/A3/M3/M2/_0_  (.A1(\V4/V2/V3/A3/M3/s1 ),
    .A2(\V4/V2/V3/A3/c2 ),
    .ZN(\V4/V2/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M3/M2/_1_  (.A(\V4/V2/V3/A3/M3/s1 ),
    .B(\V4/V2/V3/A3/c2 ),
    .Z(\V4/V2/v3 [6]));
 OR2_X1 \V4/V2/V3/A3/M3/_0_  (.A1(\V4/V2/V3/A3/M3/c1 ),
    .A2(\V4/V2/V3/A3/M3/c2 ),
    .ZN(\V4/V2/V3/A3/c3 ));
 AND2_X1 \V4/V2/V3/A3/M4/M1/_0_  (.A1(\V4/V2/V3/v4 [3]),
    .A2(net1),
    .ZN(\V4/V2/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V3/A3/M4/M1/_1_  (.A(\V4/V2/V3/v4 [3]),
    .B(net1),
    .Z(\V4/V2/V3/A3/M4/s1 ));
 AND2_X1 \V4/V2/V3/A3/M4/M2/_0_  (.A1(\V4/V2/V3/A3/M4/s1 ),
    .A2(\V4/V2/V3/A3/c3 ),
    .ZN(\V4/V2/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V3/A3/M4/M2/_1_  (.A(\V4/V2/V3/A3/M4/s1 ),
    .B(\V4/V2/V3/A3/c3 ),
    .Z(\V4/V2/v3 [7]));
 OR2_X1 \V4/V2/V3/A3/M4/_0_  (.A1(\V4/V2/V3/A3/M4/c1 ),
    .A2(\V4/V2/V3/A3/M4/c2 ),
    .ZN(\V4/V2/V3/overflow ));
 AND2_X1 \V4/V2/V3/V1/HA1/_0_  (.A1(\V4/V2/V3/V1/w2 ),
    .A2(\V4/V2/V3/V1/w1 ),
    .ZN(\V4/V2/V3/V1/w4 ));
 XOR2_X2 \V4/V2/V3/V1/HA1/_1_  (.A(\V4/V2/V3/V1/w2 ),
    .B(\V4/V2/V3/V1/w1 ),
    .Z(\V4/V2/v3 [1]));
 AND2_X1 \V4/V2/V3/V1/HA2/_0_  (.A1(\V4/V2/V3/V1/w4 ),
    .A2(\V4/V2/V3/V1/w3 ),
    .ZN(\V4/V2/V3/v1 [3]));
 XOR2_X2 \V4/V2/V3/V1/HA2/_1_  (.A(\V4/V2/V3/V1/w4 ),
    .B(\V4/V2/V3/V1/w3 ),
    .Z(\V4/V2/V3/v1 [2]));
 AND2_X1 \V4/V2/V3/V1/_0_  (.A1(net33),
    .A2(net18),
    .ZN(\V4/V2/v3 [0]));
 AND2_X1 \V4/V2/V3/V1/_1_  (.A1(net33),
    .A2(net17),
    .ZN(\V4/V2/V3/V1/w1 ));
 AND2_X1 \V4/V2/V3/V1/_2_  (.A1(net18),
    .A2(net32),
    .ZN(\V4/V2/V3/V1/w2 ));
 AND2_X1 \V4/V2/V3/V1/_3_  (.A1(net17),
    .A2(net32),
    .ZN(\V4/V2/V3/V1/w3 ));
 AND2_X1 \V4/V2/V3/V2/HA1/_0_  (.A1(\V4/V2/V3/V2/w2 ),
    .A2(\V4/V2/V3/V2/w1 ),
    .ZN(\V4/V2/V3/V2/w4 ));
 XOR2_X2 \V4/V2/V3/V2/HA1/_1_  (.A(\V4/V2/V3/V2/w2 ),
    .B(\V4/V2/V3/V2/w1 ),
    .Z(\V4/V2/V3/v2 [1]));
 AND2_X1 \V4/V2/V3/V2/HA2/_0_  (.A1(\V4/V2/V3/V2/w4 ),
    .A2(\V4/V2/V3/V2/w3 ),
    .ZN(\V4/V2/V3/v2 [3]));
 XOR2_X2 \V4/V2/V3/V2/HA2/_1_  (.A(\V4/V2/V3/V2/w4 ),
    .B(\V4/V2/V3/V2/w3 ),
    .Z(\V4/V2/V3/v2 [2]));
 AND2_X1 \V4/V2/V3/V2/_0_  (.A1(net31),
    .A2(net18),
    .ZN(\V4/V2/V3/v2 [0]));
 AND2_X1 \V4/V2/V3/V2/_1_  (.A1(net31),
    .A2(net17),
    .ZN(\V4/V2/V3/V2/w1 ));
 AND2_X1 \V4/V2/V3/V2/_2_  (.A1(net18),
    .A2(net30),
    .ZN(\V4/V2/V3/V2/w2 ));
 AND2_X1 \V4/V2/V3/V2/_3_  (.A1(net17),
    .A2(net30),
    .ZN(\V4/V2/V3/V2/w3 ));
 AND2_X1 \V4/V2/V3/V3/HA1/_0_  (.A1(\V4/V2/V3/V3/w2 ),
    .A2(\V4/V2/V3/V3/w1 ),
    .ZN(\V4/V2/V3/V3/w4 ));
 XOR2_X2 \V4/V2/V3/V3/HA1/_1_  (.A(\V4/V2/V3/V3/w2 ),
    .B(\V4/V2/V3/V3/w1 ),
    .Z(\V4/V2/V3/v3 [1]));
 AND2_X1 \V4/V2/V3/V3/HA2/_0_  (.A1(\V4/V2/V3/V3/w4 ),
    .A2(\V4/V2/V3/V3/w3 ),
    .ZN(\V4/V2/V3/v3 [3]));
 XOR2_X2 \V4/V2/V3/V3/HA2/_1_  (.A(\V4/V2/V3/V3/w4 ),
    .B(\V4/V2/V3/V3/w3 ),
    .Z(\V4/V2/V3/v3 [2]));
 AND2_X1 \V4/V2/V3/V3/_0_  (.A1(net33),
    .A2(net16),
    .ZN(\V4/V2/V3/v3 [0]));
 AND2_X1 \V4/V2/V3/V3/_1_  (.A1(net33),
    .A2(net15),
    .ZN(\V4/V2/V3/V3/w1 ));
 AND2_X1 \V4/V2/V3/V3/_2_  (.A1(net16),
    .A2(net32),
    .ZN(\V4/V2/V3/V3/w2 ));
 AND2_X1 \V4/V2/V3/V3/_3_  (.A1(net15),
    .A2(net32),
    .ZN(\V4/V2/V3/V3/w3 ));
 AND2_X1 \V4/V2/V3/V4/HA1/_0_  (.A1(\V4/V2/V3/V4/w2 ),
    .A2(\V4/V2/V3/V4/w1 ),
    .ZN(\V4/V2/V3/V4/w4 ));
 XOR2_X2 \V4/V2/V3/V4/HA1/_1_  (.A(\V4/V2/V3/V4/w2 ),
    .B(\V4/V2/V3/V4/w1 ),
    .Z(\V4/V2/V3/v4 [1]));
 AND2_X1 \V4/V2/V3/V4/HA2/_0_  (.A1(\V4/V2/V3/V4/w4 ),
    .A2(\V4/V2/V3/V4/w3 ),
    .ZN(\V4/V2/V3/v4 [3]));
 XOR2_X2 \V4/V2/V3/V4/HA2/_1_  (.A(\V4/V2/V3/V4/w4 ),
    .B(\V4/V2/V3/V4/w3 ),
    .Z(\V4/V2/V3/v4 [2]));
 AND2_X1 \V4/V2/V3/V4/_0_  (.A1(net31),
    .A2(net16),
    .ZN(\V4/V2/V3/v4 [0]));
 AND2_X1 \V4/V2/V3/V4/_1_  (.A1(net31),
    .A2(net15),
    .ZN(\V4/V2/V3/V4/w1 ));
 AND2_X1 \V4/V2/V3/V4/_2_  (.A1(net16),
    .A2(net30),
    .ZN(\V4/V2/V3/V4/w2 ));
 AND2_X1 \V4/V2/V3/V4/_3_  (.A1(net15),
    .A2(net30),
    .ZN(\V4/V2/V3/V4/w3 ));
 OR2_X1 \V4/V2/V3/_0_  (.A1(\V4/V2/V3/c1 ),
    .A2(\V4/V2/V3/c2 ),
    .ZN(\V4/V2/V3/c3 ));
 AND2_X1 \V4/V2/V4/A1/M1/M1/_0_  (.A1(\V4/V2/V4/v2 [0]),
    .A2(\V4/V2/V4/v3 [0]),
    .ZN(\V4/V2/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M1/M1/_1_  (.A(\V4/V2/V4/v2 [0]),
    .B(\V4/V2/V4/v3 [0]),
    .Z(\V4/V2/V4/A1/M1/s1 ));
 AND2_X1 \V4/V2/V4/A1/M1/M2/_0_  (.A1(\V4/V2/V4/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M1/M2/_1_  (.A(\V4/V2/V4/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/V4/s1 [0]));
 OR2_X1 \V4/V2/V4/A1/M1/_0_  (.A1(\V4/V2/V4/A1/M1/c1 ),
    .A2(\V4/V2/V4/A1/M1/c2 ),
    .ZN(\V4/V2/V4/A1/c1 ));
 AND2_X1 \V4/V2/V4/A1/M2/M1/_0_  (.A1(\V4/V2/V4/v2 [1]),
    .A2(\V4/V2/V4/v3 [1]),
    .ZN(\V4/V2/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M2/M1/_1_  (.A(\V4/V2/V4/v2 [1]),
    .B(\V4/V2/V4/v3 [1]),
    .Z(\V4/V2/V4/A1/M2/s1 ));
 AND2_X1 \V4/V2/V4/A1/M2/M2/_0_  (.A1(\V4/V2/V4/A1/M2/s1 ),
    .A2(\V4/V2/V4/A1/c1 ),
    .ZN(\V4/V2/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M2/M2/_1_  (.A(\V4/V2/V4/A1/M2/s1 ),
    .B(\V4/V2/V4/A1/c1 ),
    .Z(\V4/V2/V4/s1 [1]));
 OR2_X1 \V4/V2/V4/A1/M2/_0_  (.A1(\V4/V2/V4/A1/M2/c1 ),
    .A2(\V4/V2/V4/A1/M2/c2 ),
    .ZN(\V4/V2/V4/A1/c2 ));
 AND2_X1 \V4/V2/V4/A1/M3/M1/_0_  (.A1(\V4/V2/V4/v2 [2]),
    .A2(\V4/V2/V4/v3 [2]),
    .ZN(\V4/V2/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M3/M1/_1_  (.A(\V4/V2/V4/v2 [2]),
    .B(\V4/V2/V4/v3 [2]),
    .Z(\V4/V2/V4/A1/M3/s1 ));
 AND2_X1 \V4/V2/V4/A1/M3/M2/_0_  (.A1(\V4/V2/V4/A1/M3/s1 ),
    .A2(\V4/V2/V4/A1/c2 ),
    .ZN(\V4/V2/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M3/M2/_1_  (.A(\V4/V2/V4/A1/M3/s1 ),
    .B(\V4/V2/V4/A1/c2 ),
    .Z(\V4/V2/V4/s1 [2]));
 OR2_X1 \V4/V2/V4/A1/M3/_0_  (.A1(\V4/V2/V4/A1/M3/c1 ),
    .A2(\V4/V2/V4/A1/M3/c2 ),
    .ZN(\V4/V2/V4/A1/c3 ));
 AND2_X1 \V4/V2/V4/A1/M4/M1/_0_  (.A1(\V4/V2/V4/v2 [3]),
    .A2(\V4/V2/V4/v3 [3]),
    .ZN(\V4/V2/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A1/M4/M1/_1_  (.A(\V4/V2/V4/v2 [3]),
    .B(\V4/V2/V4/v3 [3]),
    .Z(\V4/V2/V4/A1/M4/s1 ));
 AND2_X1 \V4/V2/V4/A1/M4/M2/_0_  (.A1(\V4/V2/V4/A1/M4/s1 ),
    .A2(\V4/V2/V4/A1/c3 ),
    .ZN(\V4/V2/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A1/M4/M2/_1_  (.A(\V4/V2/V4/A1/M4/s1 ),
    .B(\V4/V2/V4/A1/c3 ),
    .Z(\V4/V2/V4/s1 [3]));
 OR2_X1 \V4/V2/V4/A1/M4/_0_  (.A1(\V4/V2/V4/A1/M4/c1 ),
    .A2(\V4/V2/V4/A1/M4/c2 ),
    .ZN(\V4/V2/V4/c1 ));
 AND2_X1 \V4/V2/V4/A2/M1/M1/_0_  (.A1(\V4/V2/V4/s1 [0]),
    .A2(\V4/V2/V4/v1 [2]),
    .ZN(\V4/V2/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M1/M1/_1_  (.A(\V4/V2/V4/s1 [0]),
    .B(\V4/V2/V4/v1 [2]),
    .Z(\V4/V2/V4/A2/M1/s1 ));
 AND2_X1 \V4/V2/V4/A2/M1/M2/_0_  (.A1(\V4/V2/V4/A2/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M1/M2/_1_  (.A(\V4/V2/V4/A2/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v4 [2]));
 OR2_X1 \V4/V2/V4/A2/M1/_0_  (.A1(\V4/V2/V4/A2/M1/c1 ),
    .A2(\V4/V2/V4/A2/M1/c2 ),
    .ZN(\V4/V2/V4/A2/c1 ));
 AND2_X1 \V4/V2/V4/A2/M2/M1/_0_  (.A1(\V4/V2/V4/s1 [1]),
    .A2(\V4/V2/V4/v1 [3]),
    .ZN(\V4/V2/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M2/M1/_1_  (.A(\V4/V2/V4/s1 [1]),
    .B(\V4/V2/V4/v1 [3]),
    .Z(\V4/V2/V4/A2/M2/s1 ));
 AND2_X1 \V4/V2/V4/A2/M2/M2/_0_  (.A1(\V4/V2/V4/A2/M2/s1 ),
    .A2(\V4/V2/V4/A2/c1 ),
    .ZN(\V4/V2/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M2/M2/_1_  (.A(\V4/V2/V4/A2/M2/s1 ),
    .B(\V4/V2/V4/A2/c1 ),
    .Z(\V4/V2/v4 [3]));
 OR2_X1 \V4/V2/V4/A2/M2/_0_  (.A1(\V4/V2/V4/A2/M2/c1 ),
    .A2(\V4/V2/V4/A2/M2/c2 ),
    .ZN(\V4/V2/V4/A2/c2 ));
 AND2_X1 \V4/V2/V4/A2/M3/M1/_0_  (.A1(\V4/V2/V4/s1 [2]),
    .A2(net1),
    .ZN(\V4/V2/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M3/M1/_1_  (.A(\V4/V2/V4/s1 [2]),
    .B(net1),
    .Z(\V4/V2/V4/A2/M3/s1 ));
 AND2_X1 \V4/V2/V4/A2/M3/M2/_0_  (.A1(\V4/V2/V4/A2/M3/s1 ),
    .A2(\V4/V2/V4/A2/c2 ),
    .ZN(\V4/V2/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M3/M2/_1_  (.A(\V4/V2/V4/A2/M3/s1 ),
    .B(\V4/V2/V4/A2/c2 ),
    .Z(\V4/V2/V4/s2 [2]));
 OR2_X1 \V4/V2/V4/A2/M3/_0_  (.A1(\V4/V2/V4/A2/M3/c1 ),
    .A2(\V4/V2/V4/A2/M3/c2 ),
    .ZN(\V4/V2/V4/A2/c3 ));
 AND2_X1 \V4/V2/V4/A2/M4/M1/_0_  (.A1(\V4/V2/V4/s1 [3]),
    .A2(net1),
    .ZN(\V4/V2/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A2/M4/M1/_1_  (.A(\V4/V2/V4/s1 [3]),
    .B(net1),
    .Z(\V4/V2/V4/A2/M4/s1 ));
 AND2_X1 \V4/V2/V4/A2/M4/M2/_0_  (.A1(\V4/V2/V4/A2/M4/s1 ),
    .A2(\V4/V2/V4/A2/c3 ),
    .ZN(\V4/V2/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A2/M4/M2/_1_  (.A(\V4/V2/V4/A2/M4/s1 ),
    .B(\V4/V2/V4/A2/c3 ),
    .Z(\V4/V2/V4/s2 [3]));
 OR2_X1 \V4/V2/V4/A2/M4/_0_  (.A1(\V4/V2/V4/A2/M4/c1 ),
    .A2(\V4/V2/V4/A2/M4/c2 ),
    .ZN(\V4/V2/V4/c2 ));
 AND2_X1 \V4/V2/V4/A3/M1/M1/_0_  (.A1(\V4/V2/V4/v4 [0]),
    .A2(\V4/V2/V4/s2 [2]),
    .ZN(\V4/V2/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M1/M1/_1_  (.A(\V4/V2/V4/v4 [0]),
    .B(\V4/V2/V4/s2 [2]),
    .Z(\V4/V2/V4/A3/M1/s1 ));
 AND2_X1 \V4/V2/V4/A3/M1/M2/_0_  (.A1(\V4/V2/V4/A3/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V2/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M1/M2/_1_  (.A(\V4/V2/V4/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V2/v4 [4]));
 OR2_X1 \V4/V2/V4/A3/M1/_0_  (.A1(\V4/V2/V4/A3/M1/c1 ),
    .A2(\V4/V2/V4/A3/M1/c2 ),
    .ZN(\V4/V2/V4/A3/c1 ));
 AND2_X1 \V4/V2/V4/A3/M2/M1/_0_  (.A1(\V4/V2/V4/v4 [1]),
    .A2(\V4/V2/V4/s2 [3]),
    .ZN(\V4/V2/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M2/M1/_1_  (.A(\V4/V2/V4/v4 [1]),
    .B(\V4/V2/V4/s2 [3]),
    .Z(\V4/V2/V4/A3/M2/s1 ));
 AND2_X1 \V4/V2/V4/A3/M2/M2/_0_  (.A1(\V4/V2/V4/A3/M2/s1 ),
    .A2(\V4/V2/V4/A3/c1 ),
    .ZN(\V4/V2/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M2/M2/_1_  (.A(\V4/V2/V4/A3/M2/s1 ),
    .B(\V4/V2/V4/A3/c1 ),
    .Z(\V4/V2/v4 [5]));
 OR2_X1 \V4/V2/V4/A3/M2/_0_  (.A1(\V4/V2/V4/A3/M2/c1 ),
    .A2(\V4/V2/V4/A3/M2/c2 ),
    .ZN(\V4/V2/V4/A3/c2 ));
 AND2_X1 \V4/V2/V4/A3/M3/M1/_0_  (.A1(\V4/V2/V4/v4 [2]),
    .A2(\V4/V2/V4/c3 ),
    .ZN(\V4/V2/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M3/M1/_1_  (.A(\V4/V2/V4/v4 [2]),
    .B(\V4/V2/V4/c3 ),
    .Z(\V4/V2/V4/A3/M3/s1 ));
 AND2_X1 \V4/V2/V4/A3/M3/M2/_0_  (.A1(\V4/V2/V4/A3/M3/s1 ),
    .A2(\V4/V2/V4/A3/c2 ),
    .ZN(\V4/V2/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M3/M2/_1_  (.A(\V4/V2/V4/A3/M3/s1 ),
    .B(\V4/V2/V4/A3/c2 ),
    .Z(\V4/V2/v4 [6]));
 OR2_X1 \V4/V2/V4/A3/M3/_0_  (.A1(\V4/V2/V4/A3/M3/c1 ),
    .A2(\V4/V2/V4/A3/M3/c2 ),
    .ZN(\V4/V2/V4/A3/c3 ));
 AND2_X1 \V4/V2/V4/A3/M4/M1/_0_  (.A1(\V4/V2/V4/v4 [3]),
    .A2(net1),
    .ZN(\V4/V2/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V2/V4/A3/M4/M1/_1_  (.A(\V4/V2/V4/v4 [3]),
    .B(net1),
    .Z(\V4/V2/V4/A3/M4/s1 ));
 AND2_X1 \V4/V2/V4/A3/M4/M2/_0_  (.A1(\V4/V2/V4/A3/M4/s1 ),
    .A2(\V4/V2/V4/A3/c3 ),
    .ZN(\V4/V2/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V2/V4/A3/M4/M2/_1_  (.A(\V4/V2/V4/A3/M4/s1 ),
    .B(\V4/V2/V4/A3/c3 ),
    .Z(\V4/V2/v4 [7]));
 OR2_X1 \V4/V2/V4/A3/M4/_0_  (.A1(\V4/V2/V4/A3/M4/c1 ),
    .A2(\V4/V2/V4/A3/M4/c2 ),
    .ZN(\V4/V2/V4/overflow ));
 AND2_X1 \V4/V2/V4/V1/HA1/_0_  (.A1(\V4/V2/V4/V1/w2 ),
    .A2(\V4/V2/V4/V1/w1 ),
    .ZN(\V4/V2/V4/V1/w4 ));
 XOR2_X2 \V4/V2/V4/V1/HA1/_1_  (.A(\V4/V2/V4/V1/w2 ),
    .B(\V4/V2/V4/V1/w1 ),
    .Z(\V4/V2/v4 [1]));
 AND2_X1 \V4/V2/V4/V1/HA2/_0_  (.A1(\V4/V2/V4/V1/w4 ),
    .A2(\V4/V2/V4/V1/w3 ),
    .ZN(\V4/V2/V4/v1 [3]));
 XOR2_X2 \V4/V2/V4/V1/HA2/_1_  (.A(\V4/V2/V4/V1/w4 ),
    .B(\V4/V2/V4/V1/w3 ),
    .Z(\V4/V2/V4/v1 [2]));
 AND2_X1 \V4/V2/V4/V1/_0_  (.A1(net29),
    .A2(net18),
    .ZN(\V4/V2/v4 [0]));
 AND2_X1 \V4/V2/V4/V1/_1_  (.A1(net29),
    .A2(net17),
    .ZN(\V4/V2/V4/V1/w1 ));
 AND2_X1 \V4/V2/V4/V1/_2_  (.A1(net18),
    .A2(net28),
    .ZN(\V4/V2/V4/V1/w2 ));
 AND2_X1 \V4/V2/V4/V1/_3_  (.A1(net17),
    .A2(net28),
    .ZN(\V4/V2/V4/V1/w3 ));
 AND2_X1 \V4/V2/V4/V2/HA1/_0_  (.A1(\V4/V2/V4/V2/w2 ),
    .A2(\V4/V2/V4/V2/w1 ),
    .ZN(\V4/V2/V4/V2/w4 ));
 XOR2_X2 \V4/V2/V4/V2/HA1/_1_  (.A(\V4/V2/V4/V2/w2 ),
    .B(\V4/V2/V4/V2/w1 ),
    .Z(\V4/V2/V4/v2 [1]));
 AND2_X1 \V4/V2/V4/V2/HA2/_0_  (.A1(\V4/V2/V4/V2/w4 ),
    .A2(\V4/V2/V4/V2/w3 ),
    .ZN(\V4/V2/V4/v2 [3]));
 XOR2_X2 \V4/V2/V4/V2/HA2/_1_  (.A(\V4/V2/V4/V2/w4 ),
    .B(\V4/V2/V4/V2/w3 ),
    .Z(\V4/V2/V4/v2 [2]));
 AND2_X1 \V4/V2/V4/V2/_0_  (.A1(net27),
    .A2(net18),
    .ZN(\V4/V2/V4/v2 [0]));
 AND2_X1 \V4/V2/V4/V2/_1_  (.A1(net27),
    .A2(net17),
    .ZN(\V4/V2/V4/V2/w1 ));
 AND2_X1 \V4/V2/V4/V2/_2_  (.A1(net18),
    .A2(net26),
    .ZN(\V4/V2/V4/V2/w2 ));
 AND2_X1 \V4/V2/V4/V2/_3_  (.A1(net17),
    .A2(net26),
    .ZN(\V4/V2/V4/V2/w3 ));
 AND2_X1 \V4/V2/V4/V3/HA1/_0_  (.A1(\V4/V2/V4/V3/w2 ),
    .A2(\V4/V2/V4/V3/w1 ),
    .ZN(\V4/V2/V4/V3/w4 ));
 XOR2_X2 \V4/V2/V4/V3/HA1/_1_  (.A(\V4/V2/V4/V3/w2 ),
    .B(\V4/V2/V4/V3/w1 ),
    .Z(\V4/V2/V4/v3 [1]));
 AND2_X1 \V4/V2/V4/V3/HA2/_0_  (.A1(\V4/V2/V4/V3/w4 ),
    .A2(\V4/V2/V4/V3/w3 ),
    .ZN(\V4/V2/V4/v3 [3]));
 XOR2_X2 \V4/V2/V4/V3/HA2/_1_  (.A(\V4/V2/V4/V3/w4 ),
    .B(\V4/V2/V4/V3/w3 ),
    .Z(\V4/V2/V4/v3 [2]));
 AND2_X1 \V4/V2/V4/V3/_0_  (.A1(net29),
    .A2(net16),
    .ZN(\V4/V2/V4/v3 [0]));
 AND2_X1 \V4/V2/V4/V3/_1_  (.A1(net29),
    .A2(net15),
    .ZN(\V4/V2/V4/V3/w1 ));
 AND2_X1 \V4/V2/V4/V3/_2_  (.A1(net16),
    .A2(net28),
    .ZN(\V4/V2/V4/V3/w2 ));
 AND2_X1 \V4/V2/V4/V3/_3_  (.A1(net15),
    .A2(net28),
    .ZN(\V4/V2/V4/V3/w3 ));
 AND2_X1 \V4/V2/V4/V4/HA1/_0_  (.A1(\V4/V2/V4/V4/w2 ),
    .A2(\V4/V2/V4/V4/w1 ),
    .ZN(\V4/V2/V4/V4/w4 ));
 XOR2_X2 \V4/V2/V4/V4/HA1/_1_  (.A(\V4/V2/V4/V4/w2 ),
    .B(\V4/V2/V4/V4/w1 ),
    .Z(\V4/V2/V4/v4 [1]));
 AND2_X1 \V4/V2/V4/V4/HA2/_0_  (.A1(\V4/V2/V4/V4/w4 ),
    .A2(\V4/V2/V4/V4/w3 ),
    .ZN(\V4/V2/V4/v4 [3]));
 XOR2_X2 \V4/V2/V4/V4/HA2/_1_  (.A(\V4/V2/V4/V4/w4 ),
    .B(\V4/V2/V4/V4/w3 ),
    .Z(\V4/V2/V4/v4 [2]));
 AND2_X1 \V4/V2/V4/V4/_0_  (.A1(net27),
    .A2(net16),
    .ZN(\V4/V2/V4/v4 [0]));
 AND2_X1 \V4/V2/V4/V4/_1_  (.A1(net27),
    .A2(net15),
    .ZN(\V4/V2/V4/V4/w1 ));
 AND2_X1 \V4/V2/V4/V4/_2_  (.A1(net16),
    .A2(net26),
    .ZN(\V4/V2/V4/V4/w2 ));
 AND2_X1 \V4/V2/V4/V4/_3_  (.A1(net15),
    .A2(net26),
    .ZN(\V4/V2/V4/V4/w3 ));
 OR2_X1 \V4/V2/V4/_0_  (.A1(\V4/V2/V4/c1 ),
    .A2(\V4/V2/V4/c2 ),
    .ZN(\V4/V2/V4/c3 ));
 OR2_X1 \V4/V2/_0_  (.A1(\V4/V2/c1 ),
    .A2(\V4/V2/c2 ),
    .ZN(\V4/V2/c3 ));
 AND2_X1 \V4/V3/A1/A1/M1/M1/_0_  (.A1(\V4/V3/v2 [0]),
    .A2(\V4/V3/v3 [0]),
    .ZN(\V4/V3/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M1/M1/_1_  (.A(\V4/V3/v2 [0]),
    .B(\V4/V3/v3 [0]),
    .Z(\V4/V3/A1/A1/M1/s1 ));
 AND2_X1 \V4/V3/A1/A1/M1/M2/_0_  (.A1(\V4/V3/A1/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M1/M2/_1_  (.A(\V4/V3/A1/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/s1 [0]));
 OR2_X1 \V4/V3/A1/A1/M1/_0_  (.A1(\V4/V3/A1/A1/M1/c1 ),
    .A2(\V4/V3/A1/A1/M1/c2 ),
    .ZN(\V4/V3/A1/A1/c1 ));
 AND2_X1 \V4/V3/A1/A1/M2/M1/_0_  (.A1(\V4/V3/v2 [1]),
    .A2(\V4/V3/v3 [1]),
    .ZN(\V4/V3/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M2/M1/_1_  (.A(\V4/V3/v2 [1]),
    .B(\V4/V3/v3 [1]),
    .Z(\V4/V3/A1/A1/M2/s1 ));
 AND2_X1 \V4/V3/A1/A1/M2/M2/_0_  (.A1(\V4/V3/A1/A1/M2/s1 ),
    .A2(\V4/V3/A1/A1/c1 ),
    .ZN(\V4/V3/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M2/M2/_1_  (.A(\V4/V3/A1/A1/M2/s1 ),
    .B(\V4/V3/A1/A1/c1 ),
    .Z(\V4/V3/s1 [1]));
 OR2_X1 \V4/V3/A1/A1/M2/_0_  (.A1(\V4/V3/A1/A1/M2/c1 ),
    .A2(\V4/V3/A1/A1/M2/c2 ),
    .ZN(\V4/V3/A1/A1/c2 ));
 AND2_X1 \V4/V3/A1/A1/M3/M1/_0_  (.A1(\V4/V3/v2 [2]),
    .A2(\V4/V3/v3 [2]),
    .ZN(\V4/V3/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M3/M1/_1_  (.A(\V4/V3/v2 [2]),
    .B(\V4/V3/v3 [2]),
    .Z(\V4/V3/A1/A1/M3/s1 ));
 AND2_X1 \V4/V3/A1/A1/M3/M2/_0_  (.A1(\V4/V3/A1/A1/M3/s1 ),
    .A2(\V4/V3/A1/A1/c2 ),
    .ZN(\V4/V3/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M3/M2/_1_  (.A(\V4/V3/A1/A1/M3/s1 ),
    .B(\V4/V3/A1/A1/c2 ),
    .Z(\V4/V3/s1 [2]));
 OR2_X1 \V4/V3/A1/A1/M3/_0_  (.A1(\V4/V3/A1/A1/M3/c1 ),
    .A2(\V4/V3/A1/A1/M3/c2 ),
    .ZN(\V4/V3/A1/A1/c3 ));
 AND2_X1 \V4/V3/A1/A1/M4/M1/_0_  (.A1(\V4/V3/v2 [3]),
    .A2(\V4/V3/v3 [3]),
    .ZN(\V4/V3/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A1/A1/M4/M1/_1_  (.A(\V4/V3/v2 [3]),
    .B(\V4/V3/v3 [3]),
    .Z(\V4/V3/A1/A1/M4/s1 ));
 AND2_X1 \V4/V3/A1/A1/M4/M2/_0_  (.A1(\V4/V3/A1/A1/M4/s1 ),
    .A2(\V4/V3/A1/A1/c3 ),
    .ZN(\V4/V3/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A1/A1/M4/M2/_1_  (.A(\V4/V3/A1/A1/M4/s1 ),
    .B(\V4/V3/A1/A1/c3 ),
    .Z(\V4/V3/s1 [3]));
 OR2_X1 \V4/V3/A1/A1/M4/_0_  (.A1(\V4/V3/A1/A1/M4/c1 ),
    .A2(\V4/V3/A1/A1/M4/c2 ),
    .ZN(\V4/V3/A1/c1 ));
 AND2_X1 \V4/V3/A1/A2/M1/M1/_0_  (.A1(\V4/V3/v2 [4]),
    .A2(\V4/V3/v3 [4]),
    .ZN(\V4/V3/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M1/M1/_1_  (.A(\V4/V3/v2 [4]),
    .B(\V4/V3/v3 [4]),
    .Z(\V4/V3/A1/A2/M1/s1 ));
 AND2_X1 \V4/V3/A1/A2/M1/M2/_0_  (.A1(\V4/V3/A1/A2/M1/s1 ),
    .A2(\V4/V3/A1/c1 ),
    .ZN(\V4/V3/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M1/M2/_1_  (.A(\V4/V3/A1/A2/M1/s1 ),
    .B(\V4/V3/A1/c1 ),
    .Z(\V4/V3/s1 [4]));
 OR2_X1 \V4/V3/A1/A2/M1/_0_  (.A1(\V4/V3/A1/A2/M1/c1 ),
    .A2(\V4/V3/A1/A2/M1/c2 ),
    .ZN(\V4/V3/A1/A2/c1 ));
 AND2_X1 \V4/V3/A1/A2/M2/M1/_0_  (.A1(\V4/V3/v2 [5]),
    .A2(\V4/V3/v3 [5]),
    .ZN(\V4/V3/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M2/M1/_1_  (.A(\V4/V3/v2 [5]),
    .B(\V4/V3/v3 [5]),
    .Z(\V4/V3/A1/A2/M2/s1 ));
 AND2_X1 \V4/V3/A1/A2/M2/M2/_0_  (.A1(\V4/V3/A1/A2/M2/s1 ),
    .A2(\V4/V3/A1/A2/c1 ),
    .ZN(\V4/V3/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M2/M2/_1_  (.A(\V4/V3/A1/A2/M2/s1 ),
    .B(\V4/V3/A1/A2/c1 ),
    .Z(\V4/V3/s1 [5]));
 OR2_X1 \V4/V3/A1/A2/M2/_0_  (.A1(\V4/V3/A1/A2/M2/c1 ),
    .A2(\V4/V3/A1/A2/M2/c2 ),
    .ZN(\V4/V3/A1/A2/c2 ));
 AND2_X1 \V4/V3/A1/A2/M3/M1/_0_  (.A1(\V4/V3/v2 [6]),
    .A2(\V4/V3/v3 [6]),
    .ZN(\V4/V3/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M3/M1/_1_  (.A(\V4/V3/v2 [6]),
    .B(\V4/V3/v3 [6]),
    .Z(\V4/V3/A1/A2/M3/s1 ));
 AND2_X1 \V4/V3/A1/A2/M3/M2/_0_  (.A1(\V4/V3/A1/A2/M3/s1 ),
    .A2(\V4/V3/A1/A2/c2 ),
    .ZN(\V4/V3/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M3/M2/_1_  (.A(\V4/V3/A1/A2/M3/s1 ),
    .B(\V4/V3/A1/A2/c2 ),
    .Z(\V4/V3/s1 [6]));
 OR2_X1 \V4/V3/A1/A2/M3/_0_  (.A1(\V4/V3/A1/A2/M3/c1 ),
    .A2(\V4/V3/A1/A2/M3/c2 ),
    .ZN(\V4/V3/A1/A2/c3 ));
 AND2_X1 \V4/V3/A1/A2/M4/M1/_0_  (.A1(\V4/V3/v2 [7]),
    .A2(\V4/V3/v3 [7]),
    .ZN(\V4/V3/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A1/A2/M4/M1/_1_  (.A(\V4/V3/v2 [7]),
    .B(\V4/V3/v3 [7]),
    .Z(\V4/V3/A1/A2/M4/s1 ));
 AND2_X1 \V4/V3/A1/A2/M4/M2/_0_  (.A1(\V4/V3/A1/A2/M4/s1 ),
    .A2(\V4/V3/A1/A2/c3 ),
    .ZN(\V4/V3/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A1/A2/M4/M2/_1_  (.A(\V4/V3/A1/A2/M4/s1 ),
    .B(\V4/V3/A1/A2/c3 ),
    .Z(\V4/V3/s1 [7]));
 OR2_X1 \V4/V3/A1/A2/M4/_0_  (.A1(\V4/V3/A1/A2/M4/c1 ),
    .A2(\V4/V3/A1/A2/M4/c2 ),
    .ZN(\V4/V3/c1 ));
 AND2_X1 \V4/V3/A2/A1/M1/M1/_0_  (.A1(\V4/V3/s1 [0]),
    .A2(\V4/V3/v1 [4]),
    .ZN(\V4/V3/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M1/M1/_1_  (.A(\V4/V3/s1 [0]),
    .B(\V4/V3/v1 [4]),
    .Z(\V4/V3/A2/A1/M1/s1 ));
 AND2_X1 \V4/V3/A2/A1/M1/M2/_0_  (.A1(\V4/V3/A2/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M1/M2/_1_  (.A(\V4/V3/A2/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/v3 [4]));
 OR2_X1 \V4/V3/A2/A1/M1/_0_  (.A1(\V4/V3/A2/A1/M1/c1 ),
    .A2(\V4/V3/A2/A1/M1/c2 ),
    .ZN(\V4/V3/A2/A1/c1 ));
 AND2_X1 \V4/V3/A2/A1/M2/M1/_0_  (.A1(\V4/V3/s1 [1]),
    .A2(\V4/V3/v1 [5]),
    .ZN(\V4/V3/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M2/M1/_1_  (.A(\V4/V3/s1 [1]),
    .B(\V4/V3/v1 [5]),
    .Z(\V4/V3/A2/A1/M2/s1 ));
 AND2_X1 \V4/V3/A2/A1/M2/M2/_0_  (.A1(\V4/V3/A2/A1/M2/s1 ),
    .A2(\V4/V3/A2/A1/c1 ),
    .ZN(\V4/V3/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M2/M2/_1_  (.A(\V4/V3/A2/A1/M2/s1 ),
    .B(\V4/V3/A2/A1/c1 ),
    .Z(\V4/v3 [5]));
 OR2_X1 \V4/V3/A2/A1/M2/_0_  (.A1(\V4/V3/A2/A1/M2/c1 ),
    .A2(\V4/V3/A2/A1/M2/c2 ),
    .ZN(\V4/V3/A2/A1/c2 ));
 AND2_X1 \V4/V3/A2/A1/M3/M1/_0_  (.A1(\V4/V3/s1 [2]),
    .A2(\V4/V3/v1 [6]),
    .ZN(\V4/V3/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M3/M1/_1_  (.A(\V4/V3/s1 [2]),
    .B(\V4/V3/v1 [6]),
    .Z(\V4/V3/A2/A1/M3/s1 ));
 AND2_X1 \V4/V3/A2/A1/M3/M2/_0_  (.A1(\V4/V3/A2/A1/M3/s1 ),
    .A2(\V4/V3/A2/A1/c2 ),
    .ZN(\V4/V3/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M3/M2/_1_  (.A(\V4/V3/A2/A1/M3/s1 ),
    .B(\V4/V3/A2/A1/c2 ),
    .Z(\V4/v3 [6]));
 OR2_X1 \V4/V3/A2/A1/M3/_0_  (.A1(\V4/V3/A2/A1/M3/c1 ),
    .A2(\V4/V3/A2/A1/M3/c2 ),
    .ZN(\V4/V3/A2/A1/c3 ));
 AND2_X1 \V4/V3/A2/A1/M4/M1/_0_  (.A1(\V4/V3/s1 [3]),
    .A2(\V4/V3/v1 [7]),
    .ZN(\V4/V3/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A2/A1/M4/M1/_1_  (.A(\V4/V3/s1 [3]),
    .B(\V4/V3/v1 [7]),
    .Z(\V4/V3/A2/A1/M4/s1 ));
 AND2_X1 \V4/V3/A2/A1/M4/M2/_0_  (.A1(\V4/V3/A2/A1/M4/s1 ),
    .A2(\V4/V3/A2/A1/c3 ),
    .ZN(\V4/V3/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A2/A1/M4/M2/_1_  (.A(\V4/V3/A2/A1/M4/s1 ),
    .B(\V4/V3/A2/A1/c3 ),
    .Z(\V4/v3 [7]));
 OR2_X1 \V4/V3/A2/A1/M4/_0_  (.A1(\V4/V3/A2/A1/M4/c1 ),
    .A2(\V4/V3/A2/A1/M4/c2 ),
    .ZN(\V4/V3/A2/c1 ));
 AND2_X1 \V4/V3/A2/A2/M1/M1/_0_  (.A1(\V4/V3/s1 [4]),
    .A2(net10),
    .ZN(\V4/V3/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M1/M1/_1_  (.A(\V4/V3/s1 [4]),
    .B(net10),
    .Z(\V4/V3/A2/A2/M1/s1 ));
 AND2_X1 \V4/V3/A2/A2/M1/M2/_0_  (.A1(\V4/V3/A2/A2/M1/s1 ),
    .A2(\V4/V3/A2/c1 ),
    .ZN(\V4/V3/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M1/M2/_1_  (.A(\V4/V3/A2/A2/M1/s1 ),
    .B(\V4/V3/A2/c1 ),
    .Z(\V4/V3/s2 [4]));
 OR2_X1 \V4/V3/A2/A2/M1/_0_  (.A1(\V4/V3/A2/A2/M1/c1 ),
    .A2(\V4/V3/A2/A2/M1/c2 ),
    .ZN(\V4/V3/A2/A2/c1 ));
 AND2_X1 \V4/V3/A2/A2/M2/M1/_0_  (.A1(\V4/V3/s1 [5]),
    .A2(net10),
    .ZN(\V4/V3/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M2/M1/_1_  (.A(\V4/V3/s1 [5]),
    .B(net10),
    .Z(\V4/V3/A2/A2/M2/s1 ));
 AND2_X1 \V4/V3/A2/A2/M2/M2/_0_  (.A1(\V4/V3/A2/A2/M2/s1 ),
    .A2(\V4/V3/A2/A2/c1 ),
    .ZN(\V4/V3/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M2/M2/_1_  (.A(\V4/V3/A2/A2/M2/s1 ),
    .B(\V4/V3/A2/A2/c1 ),
    .Z(\V4/V3/s2 [5]));
 OR2_X1 \V4/V3/A2/A2/M2/_0_  (.A1(\V4/V3/A2/A2/M2/c1 ),
    .A2(\V4/V3/A2/A2/M2/c2 ),
    .ZN(\V4/V3/A2/A2/c2 ));
 AND2_X1 \V4/V3/A2/A2/M3/M1/_0_  (.A1(\V4/V3/s1 [6]),
    .A2(net10),
    .ZN(\V4/V3/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M3/M1/_1_  (.A(\V4/V3/s1 [6]),
    .B(net10),
    .Z(\V4/V3/A2/A2/M3/s1 ));
 AND2_X1 \V4/V3/A2/A2/M3/M2/_0_  (.A1(\V4/V3/A2/A2/M3/s1 ),
    .A2(\V4/V3/A2/A2/c2 ),
    .ZN(\V4/V3/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M3/M2/_1_  (.A(\V4/V3/A2/A2/M3/s1 ),
    .B(\V4/V3/A2/A2/c2 ),
    .Z(\V4/V3/s2 [6]));
 OR2_X1 \V4/V3/A2/A2/M3/_0_  (.A1(\V4/V3/A2/A2/M3/c1 ),
    .A2(\V4/V3/A2/A2/M3/c2 ),
    .ZN(\V4/V3/A2/A2/c3 ));
 AND2_X1 \V4/V3/A2/A2/M4/M1/_0_  (.A1(\V4/V3/s1 [7]),
    .A2(net10),
    .ZN(\V4/V3/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A2/A2/M4/M1/_1_  (.A(\V4/V3/s1 [7]),
    .B(net10),
    .Z(\V4/V3/A2/A2/M4/s1 ));
 AND2_X1 \V4/V3/A2/A2/M4/M2/_0_  (.A1(\V4/V3/A2/A2/M4/s1 ),
    .A2(\V4/V3/A2/A2/c3 ),
    .ZN(\V4/V3/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A2/A2/M4/M2/_1_  (.A(\V4/V3/A2/A2/M4/s1 ),
    .B(\V4/V3/A2/A2/c3 ),
    .Z(\V4/V3/s2 [7]));
 OR2_X1 \V4/V3/A2/A2/M4/_0_  (.A1(\V4/V3/A2/A2/M4/c1 ),
    .A2(\V4/V3/A2/A2/M4/c2 ),
    .ZN(\V4/V3/c2 ));
 AND2_X1 \V4/V3/A3/A1/M1/M1/_0_  (.A1(\V4/V3/v4 [0]),
    .A2(\V4/V3/s2 [4]),
    .ZN(\V4/V3/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M1/M1/_1_  (.A(\V4/V3/v4 [0]),
    .B(\V4/V3/s2 [4]),
    .Z(\V4/V3/A3/A1/M1/s1 ));
 AND2_X1 \V4/V3/A3/A1/M1/M2/_0_  (.A1(\V4/V3/A3/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M1/M2/_1_  (.A(\V4/V3/A3/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/v3 [8]));
 OR2_X1 \V4/V3/A3/A1/M1/_0_  (.A1(\V4/V3/A3/A1/M1/c1 ),
    .A2(\V4/V3/A3/A1/M1/c2 ),
    .ZN(\V4/V3/A3/A1/c1 ));
 AND2_X1 \V4/V3/A3/A1/M2/M1/_0_  (.A1(\V4/V3/v4 [1]),
    .A2(\V4/V3/s2 [5]),
    .ZN(\V4/V3/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M2/M1/_1_  (.A(\V4/V3/v4 [1]),
    .B(\V4/V3/s2 [5]),
    .Z(\V4/V3/A3/A1/M2/s1 ));
 AND2_X1 \V4/V3/A3/A1/M2/M2/_0_  (.A1(\V4/V3/A3/A1/M2/s1 ),
    .A2(\V4/V3/A3/A1/c1 ),
    .ZN(\V4/V3/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M2/M2/_1_  (.A(\V4/V3/A3/A1/M2/s1 ),
    .B(\V4/V3/A3/A1/c1 ),
    .Z(\V4/v3 [9]));
 OR2_X1 \V4/V3/A3/A1/M2/_0_  (.A1(\V4/V3/A3/A1/M2/c1 ),
    .A2(\V4/V3/A3/A1/M2/c2 ),
    .ZN(\V4/V3/A3/A1/c2 ));
 AND2_X1 \V4/V3/A3/A1/M3/M1/_0_  (.A1(\V4/V3/v4 [2]),
    .A2(\V4/V3/s2 [6]),
    .ZN(\V4/V3/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M3/M1/_1_  (.A(\V4/V3/v4 [2]),
    .B(\V4/V3/s2 [6]),
    .Z(\V4/V3/A3/A1/M3/s1 ));
 AND2_X1 \V4/V3/A3/A1/M3/M2/_0_  (.A1(\V4/V3/A3/A1/M3/s1 ),
    .A2(\V4/V3/A3/A1/c2 ),
    .ZN(\V4/V3/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M3/M2/_1_  (.A(\V4/V3/A3/A1/M3/s1 ),
    .B(\V4/V3/A3/A1/c2 ),
    .Z(\V4/v3 [10]));
 OR2_X1 \V4/V3/A3/A1/M3/_0_  (.A1(\V4/V3/A3/A1/M3/c1 ),
    .A2(\V4/V3/A3/A1/M3/c2 ),
    .ZN(\V4/V3/A3/A1/c3 ));
 AND2_X1 \V4/V3/A3/A1/M4/M1/_0_  (.A1(\V4/V3/v4 [3]),
    .A2(\V4/V3/s2 [7]),
    .ZN(\V4/V3/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V3/A3/A1/M4/M1/_1_  (.A(\V4/V3/v4 [3]),
    .B(\V4/V3/s2 [7]),
    .Z(\V4/V3/A3/A1/M4/s1 ));
 AND2_X1 \V4/V3/A3/A1/M4/M2/_0_  (.A1(\V4/V3/A3/A1/M4/s1 ),
    .A2(\V4/V3/A3/A1/c3 ),
    .ZN(\V4/V3/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V3/A3/A1/M4/M2/_1_  (.A(\V4/V3/A3/A1/M4/s1 ),
    .B(\V4/V3/A3/A1/c3 ),
    .Z(\V4/v3 [11]));
 OR2_X1 \V4/V3/A3/A1/M4/_0_  (.A1(\V4/V3/A3/A1/M4/c1 ),
    .A2(\V4/V3/A3/A1/M4/c2 ),
    .ZN(\V4/V3/A3/c1 ));
 AND2_X1 \V4/V3/A3/A2/M1/M1/_0_  (.A1(\V4/V3/v4 [4]),
    .A2(\V4/V3/c3 ),
    .ZN(\V4/V3/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M1/M1/_1_  (.A(\V4/V3/v4 [4]),
    .B(\V4/V3/c3 ),
    .Z(\V4/V3/A3/A2/M1/s1 ));
 AND2_X1 \V4/V3/A3/A2/M1/M2/_0_  (.A1(\V4/V3/A3/A2/M1/s1 ),
    .A2(\V4/V3/A3/c1 ),
    .ZN(\V4/V3/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M1/M2/_1_  (.A(\V4/V3/A3/A2/M1/s1 ),
    .B(\V4/V3/A3/c1 ),
    .Z(\V4/v3 [12]));
 OR2_X1 \V4/V3/A3/A2/M1/_0_  (.A1(\V4/V3/A3/A2/M1/c1 ),
    .A2(\V4/V3/A3/A2/M1/c2 ),
    .ZN(\V4/V3/A3/A2/c1 ));
 AND2_X1 \V4/V3/A3/A2/M2/M1/_0_  (.A1(\V4/V3/v4 [5]),
    .A2(net10),
    .ZN(\V4/V3/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M2/M1/_1_  (.A(\V4/V3/v4 [5]),
    .B(net10),
    .Z(\V4/V3/A3/A2/M2/s1 ));
 AND2_X1 \V4/V3/A3/A2/M2/M2/_0_  (.A1(\V4/V3/A3/A2/M2/s1 ),
    .A2(\V4/V3/A3/A2/c1 ),
    .ZN(\V4/V3/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M2/M2/_1_  (.A(\V4/V3/A3/A2/M2/s1 ),
    .B(\V4/V3/A3/A2/c1 ),
    .Z(\V4/v3 [13]));
 OR2_X1 \V4/V3/A3/A2/M2/_0_  (.A1(\V4/V3/A3/A2/M2/c1 ),
    .A2(\V4/V3/A3/A2/M2/c2 ),
    .ZN(\V4/V3/A3/A2/c2 ));
 AND2_X1 \V4/V3/A3/A2/M3/M1/_0_  (.A1(\V4/V3/v4 [6]),
    .A2(net10),
    .ZN(\V4/V3/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M3/M1/_1_  (.A(\V4/V3/v4 [6]),
    .B(net10),
    .Z(\V4/V3/A3/A2/M3/s1 ));
 AND2_X1 \V4/V3/A3/A2/M3/M2/_0_  (.A1(\V4/V3/A3/A2/M3/s1 ),
    .A2(\V4/V3/A3/A2/c2 ),
    .ZN(\V4/V3/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M3/M2/_1_  (.A(\V4/V3/A3/A2/M3/s1 ),
    .B(\V4/V3/A3/A2/c2 ),
    .Z(\V4/v3 [14]));
 OR2_X1 \V4/V3/A3/A2/M3/_0_  (.A1(\V4/V3/A3/A2/M3/c1 ),
    .A2(\V4/V3/A3/A2/M3/c2 ),
    .ZN(\V4/V3/A3/A2/c3 ));
 AND2_X1 \V4/V3/A3/A2/M4/M1/_0_  (.A1(\V4/V3/v4 [7]),
    .A2(net10),
    .ZN(\V4/V3/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V3/A3/A2/M4/M1/_1_  (.A(\V4/V3/v4 [7]),
    .B(net10),
    .Z(\V4/V3/A3/A2/M4/s1 ));
 AND2_X1 \V4/V3/A3/A2/M4/M2/_0_  (.A1(\V4/V3/A3/A2/M4/s1 ),
    .A2(\V4/V3/A3/A2/c3 ),
    .ZN(\V4/V3/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V3/A3/A2/M4/M2/_1_  (.A(\V4/V3/A3/A2/M4/s1 ),
    .B(\V4/V3/A3/A2/c3 ),
    .Z(\V4/v3 [15]));
 OR2_X1 \V4/V3/A3/A2/M4/_0_  (.A1(\V4/V3/A3/A2/M4/c1 ),
    .A2(\V4/V3/A3/A2/M4/c2 ),
    .ZN(\V4/V3/overflow ));
 AND2_X1 \V4/V3/V1/A1/M1/M1/_0_  (.A1(\V4/V3/V1/v2 [0]),
    .A2(\V4/V3/V1/v3 [0]),
    .ZN(\V4/V3/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M1/M1/_1_  (.A(\V4/V3/V1/v2 [0]),
    .B(\V4/V3/V1/v3 [0]),
    .Z(\V4/V3/V1/A1/M1/s1 ));
 AND2_X1 \V4/V3/V1/A1/M1/M2/_0_  (.A1(\V4/V3/V1/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M1/M2/_1_  (.A(\V4/V3/V1/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/V1/s1 [0]));
 OR2_X1 \V4/V3/V1/A1/M1/_0_  (.A1(\V4/V3/V1/A1/M1/c1 ),
    .A2(\V4/V3/V1/A1/M1/c2 ),
    .ZN(\V4/V3/V1/A1/c1 ));
 AND2_X1 \V4/V3/V1/A1/M2/M1/_0_  (.A1(\V4/V3/V1/v2 [1]),
    .A2(\V4/V3/V1/v3 [1]),
    .ZN(\V4/V3/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M2/M1/_1_  (.A(\V4/V3/V1/v2 [1]),
    .B(\V4/V3/V1/v3 [1]),
    .Z(\V4/V3/V1/A1/M2/s1 ));
 AND2_X1 \V4/V3/V1/A1/M2/M2/_0_  (.A1(\V4/V3/V1/A1/M2/s1 ),
    .A2(\V4/V3/V1/A1/c1 ),
    .ZN(\V4/V3/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M2/M2/_1_  (.A(\V4/V3/V1/A1/M2/s1 ),
    .B(\V4/V3/V1/A1/c1 ),
    .Z(\V4/V3/V1/s1 [1]));
 OR2_X1 \V4/V3/V1/A1/M2/_0_  (.A1(\V4/V3/V1/A1/M2/c1 ),
    .A2(\V4/V3/V1/A1/M2/c2 ),
    .ZN(\V4/V3/V1/A1/c2 ));
 AND2_X1 \V4/V3/V1/A1/M3/M1/_0_  (.A1(\V4/V3/V1/v2 [2]),
    .A2(\V4/V3/V1/v3 [2]),
    .ZN(\V4/V3/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M3/M1/_1_  (.A(\V4/V3/V1/v2 [2]),
    .B(\V4/V3/V1/v3 [2]),
    .Z(\V4/V3/V1/A1/M3/s1 ));
 AND2_X1 \V4/V3/V1/A1/M3/M2/_0_  (.A1(\V4/V3/V1/A1/M3/s1 ),
    .A2(\V4/V3/V1/A1/c2 ),
    .ZN(\V4/V3/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M3/M2/_1_  (.A(\V4/V3/V1/A1/M3/s1 ),
    .B(\V4/V3/V1/A1/c2 ),
    .Z(\V4/V3/V1/s1 [2]));
 OR2_X1 \V4/V3/V1/A1/M3/_0_  (.A1(\V4/V3/V1/A1/M3/c1 ),
    .A2(\V4/V3/V1/A1/M3/c2 ),
    .ZN(\V4/V3/V1/A1/c3 ));
 AND2_X1 \V4/V3/V1/A1/M4/M1/_0_  (.A1(\V4/V3/V1/v2 [3]),
    .A2(\V4/V3/V1/v3 [3]),
    .ZN(\V4/V3/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A1/M4/M1/_1_  (.A(\V4/V3/V1/v2 [3]),
    .B(\V4/V3/V1/v3 [3]),
    .Z(\V4/V3/V1/A1/M4/s1 ));
 AND2_X1 \V4/V3/V1/A1/M4/M2/_0_  (.A1(\V4/V3/V1/A1/M4/s1 ),
    .A2(\V4/V3/V1/A1/c3 ),
    .ZN(\V4/V3/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A1/M4/M2/_1_  (.A(\V4/V3/V1/A1/M4/s1 ),
    .B(\V4/V3/V1/A1/c3 ),
    .Z(\V4/V3/V1/s1 [3]));
 OR2_X1 \V4/V3/V1/A1/M4/_0_  (.A1(\V4/V3/V1/A1/M4/c1 ),
    .A2(\V4/V3/V1/A1/M4/c2 ),
    .ZN(\V4/V3/V1/c1 ));
 AND2_X1 \V4/V3/V1/A2/M1/M1/_0_  (.A1(\V4/V3/V1/s1 [0]),
    .A2(\V4/V3/V1/v1 [2]),
    .ZN(\V4/V3/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M1/M1/_1_  (.A(\V4/V3/V1/s1 [0]),
    .B(\V4/V3/V1/v1 [2]),
    .Z(\V4/V3/V1/A2/M1/s1 ));
 AND2_X1 \V4/V3/V1/A2/M1/M2/_0_  (.A1(\V4/V3/V1/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M1/M2/_1_  (.A(\V4/V3/V1/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/v3 [2]));
 OR2_X1 \V4/V3/V1/A2/M1/_0_  (.A1(\V4/V3/V1/A2/M1/c1 ),
    .A2(\V4/V3/V1/A2/M1/c2 ),
    .ZN(\V4/V3/V1/A2/c1 ));
 AND2_X1 \V4/V3/V1/A2/M2/M1/_0_  (.A1(\V4/V3/V1/s1 [1]),
    .A2(\V4/V3/V1/v1 [3]),
    .ZN(\V4/V3/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M2/M1/_1_  (.A(\V4/V3/V1/s1 [1]),
    .B(\V4/V3/V1/v1 [3]),
    .Z(\V4/V3/V1/A2/M2/s1 ));
 AND2_X1 \V4/V3/V1/A2/M2/M2/_0_  (.A1(\V4/V3/V1/A2/M2/s1 ),
    .A2(\V4/V3/V1/A2/c1 ),
    .ZN(\V4/V3/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M2/M2/_1_  (.A(\V4/V3/V1/A2/M2/s1 ),
    .B(\V4/V3/V1/A2/c1 ),
    .Z(\V4/v3 [3]));
 OR2_X1 \V4/V3/V1/A2/M2/_0_  (.A1(\V4/V3/V1/A2/M2/c1 ),
    .A2(\V4/V3/V1/A2/M2/c2 ),
    .ZN(\V4/V3/V1/A2/c2 ));
 AND2_X1 \V4/V3/V1/A2/M3/M1/_0_  (.A1(\V4/V3/V1/s1 [2]),
    .A2(net10),
    .ZN(\V4/V3/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M3/M1/_1_  (.A(\V4/V3/V1/s1 [2]),
    .B(net10),
    .Z(\V4/V3/V1/A2/M3/s1 ));
 AND2_X1 \V4/V3/V1/A2/M3/M2/_0_  (.A1(\V4/V3/V1/A2/M3/s1 ),
    .A2(\V4/V3/V1/A2/c2 ),
    .ZN(\V4/V3/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M3/M2/_1_  (.A(\V4/V3/V1/A2/M3/s1 ),
    .B(\V4/V3/V1/A2/c2 ),
    .Z(\V4/V3/V1/s2 [2]));
 OR2_X1 \V4/V3/V1/A2/M3/_0_  (.A1(\V4/V3/V1/A2/M3/c1 ),
    .A2(\V4/V3/V1/A2/M3/c2 ),
    .ZN(\V4/V3/V1/A2/c3 ));
 AND2_X1 \V4/V3/V1/A2/M4/M1/_0_  (.A1(\V4/V3/V1/s1 [3]),
    .A2(net10),
    .ZN(\V4/V3/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A2/M4/M1/_1_  (.A(\V4/V3/V1/s1 [3]),
    .B(net10),
    .Z(\V4/V3/V1/A2/M4/s1 ));
 AND2_X1 \V4/V3/V1/A2/M4/M2/_0_  (.A1(\V4/V3/V1/A2/M4/s1 ),
    .A2(\V4/V3/V1/A2/c3 ),
    .ZN(\V4/V3/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A2/M4/M2/_1_  (.A(\V4/V3/V1/A2/M4/s1 ),
    .B(\V4/V3/V1/A2/c3 ),
    .Z(\V4/V3/V1/s2 [3]));
 OR2_X1 \V4/V3/V1/A2/M4/_0_  (.A1(\V4/V3/V1/A2/M4/c1 ),
    .A2(\V4/V3/V1/A2/M4/c2 ),
    .ZN(\V4/V3/V1/c2 ));
 AND2_X1 \V4/V3/V1/A3/M1/M1/_0_  (.A1(\V4/V3/V1/v4 [0]),
    .A2(\V4/V3/V1/s2 [2]),
    .ZN(\V4/V3/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M1/M1/_1_  (.A(\V4/V3/V1/v4 [0]),
    .B(\V4/V3/V1/s2 [2]),
    .Z(\V4/V3/V1/A3/M1/s1 ));
 AND2_X1 \V4/V3/V1/A3/M1/M2/_0_  (.A1(\V4/V3/V1/A3/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M1/M2/_1_  (.A(\V4/V3/V1/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v1 [4]));
 OR2_X1 \V4/V3/V1/A3/M1/_0_  (.A1(\V4/V3/V1/A3/M1/c1 ),
    .A2(\V4/V3/V1/A3/M1/c2 ),
    .ZN(\V4/V3/V1/A3/c1 ));
 AND2_X1 \V4/V3/V1/A3/M2/M1/_0_  (.A1(\V4/V3/V1/v4 [1]),
    .A2(\V4/V3/V1/s2 [3]),
    .ZN(\V4/V3/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M2/M1/_1_  (.A(\V4/V3/V1/v4 [1]),
    .B(\V4/V3/V1/s2 [3]),
    .Z(\V4/V3/V1/A3/M2/s1 ));
 AND2_X1 \V4/V3/V1/A3/M2/M2/_0_  (.A1(\V4/V3/V1/A3/M2/s1 ),
    .A2(\V4/V3/V1/A3/c1 ),
    .ZN(\V4/V3/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M2/M2/_1_  (.A(\V4/V3/V1/A3/M2/s1 ),
    .B(\V4/V3/V1/A3/c1 ),
    .Z(\V4/V3/v1 [5]));
 OR2_X1 \V4/V3/V1/A3/M2/_0_  (.A1(\V4/V3/V1/A3/M2/c1 ),
    .A2(\V4/V3/V1/A3/M2/c2 ),
    .ZN(\V4/V3/V1/A3/c2 ));
 AND2_X1 \V4/V3/V1/A3/M3/M1/_0_  (.A1(\V4/V3/V1/v4 [2]),
    .A2(\V4/V3/V1/c3 ),
    .ZN(\V4/V3/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M3/M1/_1_  (.A(\V4/V3/V1/v4 [2]),
    .B(\V4/V3/V1/c3 ),
    .Z(\V4/V3/V1/A3/M3/s1 ));
 AND2_X1 \V4/V3/V1/A3/M3/M2/_0_  (.A1(\V4/V3/V1/A3/M3/s1 ),
    .A2(\V4/V3/V1/A3/c2 ),
    .ZN(\V4/V3/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M3/M2/_1_  (.A(\V4/V3/V1/A3/M3/s1 ),
    .B(\V4/V3/V1/A3/c2 ),
    .Z(\V4/V3/v1 [6]));
 OR2_X1 \V4/V3/V1/A3/M3/_0_  (.A1(\V4/V3/V1/A3/M3/c1 ),
    .A2(\V4/V3/V1/A3/M3/c2 ),
    .ZN(\V4/V3/V1/A3/c3 ));
 AND2_X1 \V4/V3/V1/A3/M4/M1/_0_  (.A1(\V4/V3/V1/v4 [3]),
    .A2(net10),
    .ZN(\V4/V3/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V1/A3/M4/M1/_1_  (.A(\V4/V3/V1/v4 [3]),
    .B(net10),
    .Z(\V4/V3/V1/A3/M4/s1 ));
 AND2_X1 \V4/V3/V1/A3/M4/M2/_0_  (.A1(\V4/V3/V1/A3/M4/s1 ),
    .A2(\V4/V3/V1/A3/c3 ),
    .ZN(\V4/V3/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V1/A3/M4/M2/_1_  (.A(\V4/V3/V1/A3/M4/s1 ),
    .B(\V4/V3/V1/A3/c3 ),
    .Z(\V4/V3/v1 [7]));
 OR2_X1 \V4/V3/V1/A3/M4/_0_  (.A1(\V4/V3/V1/A3/M4/c1 ),
    .A2(\V4/V3/V1/A3/M4/c2 ),
    .ZN(\V4/V3/V1/overflow ));
 AND2_X1 \V4/V3/V1/V1/HA1/_0_  (.A1(\V4/V3/V1/V1/w2 ),
    .A2(\V4/V3/V1/V1/w1 ),
    .ZN(\V4/V3/V1/V1/w4 ));
 XOR2_X2 \V4/V3/V1/V1/HA1/_1_  (.A(\V4/V3/V1/V1/w2 ),
    .B(\V4/V3/V1/V1/w1 ),
    .Z(\V4/v3 [1]));
 AND2_X1 \V4/V3/V1/V1/HA2/_0_  (.A1(\V4/V3/V1/V1/w4 ),
    .A2(\V4/V3/V1/V1/w3 ),
    .ZN(\V4/V3/V1/v1 [3]));
 XOR2_X2 \V4/V3/V1/V1/HA2/_1_  (.A(\V4/V3/V1/V1/w4 ),
    .B(\V4/V3/V1/V1/w3 ),
    .Z(\V4/V3/V1/v1 [2]));
 AND2_X1 \V4/V3/V1/V1/_0_  (.A1(net41),
    .A2(net14),
    .ZN(\V4/v3 [0]));
 AND2_X1 \V4/V3/V1/V1/_1_  (.A1(net41),
    .A2(B[25]),
    .ZN(\V4/V3/V1/V1/w1 ));
 AND2_X1 \V4/V3/V1/V1/_2_  (.A1(net14),
    .A2(net40),
    .ZN(\V4/V3/V1/V1/w2 ));
 AND2_X1 \V4/V3/V1/V1/_3_  (.A1(B[25]),
    .A2(net40),
    .ZN(\V4/V3/V1/V1/w3 ));
 AND2_X1 \V4/V3/V1/V2/HA1/_0_  (.A1(\V4/V3/V1/V2/w2 ),
    .A2(\V4/V3/V1/V2/w1 ),
    .ZN(\V4/V3/V1/V2/w4 ));
 XOR2_X2 \V4/V3/V1/V2/HA1/_1_  (.A(\V4/V3/V1/V2/w2 ),
    .B(\V4/V3/V1/V2/w1 ),
    .Z(\V4/V3/V1/v2 [1]));
 AND2_X1 \V4/V3/V1/V2/HA2/_0_  (.A1(\V4/V3/V1/V2/w4 ),
    .A2(\V4/V3/V1/V2/w3 ),
    .ZN(\V4/V3/V1/v2 [3]));
 XOR2_X2 \V4/V3/V1/V2/HA2/_1_  (.A(\V4/V3/V1/V2/w4 ),
    .B(\V4/V3/V1/V2/w3 ),
    .Z(\V4/V3/V1/v2 [2]));
 AND2_X1 \V4/V3/V1/V2/_0_  (.A1(net39),
    .A2(net14),
    .ZN(\V4/V3/V1/v2 [0]));
 AND2_X1 \V4/V3/V1/V2/_1_  (.A1(net39),
    .A2(B[25]),
    .ZN(\V4/V3/V1/V2/w1 ));
 AND2_X1 \V4/V3/V1/V2/_2_  (.A1(net14),
    .A2(net38),
    .ZN(\V4/V3/V1/V2/w2 ));
 AND2_X1 \V4/V3/V1/V2/_3_  (.A1(B[25]),
    .A2(net38),
    .ZN(\V4/V3/V1/V2/w3 ));
 AND2_X1 \V4/V3/V1/V3/HA1/_0_  (.A1(\V4/V3/V1/V3/w2 ),
    .A2(\V4/V3/V1/V3/w1 ),
    .ZN(\V4/V3/V1/V3/w4 ));
 XOR2_X2 \V4/V3/V1/V3/HA1/_1_  (.A(\V4/V3/V1/V3/w2 ),
    .B(\V4/V3/V1/V3/w1 ),
    .Z(\V4/V3/V1/v3 [1]));
 AND2_X1 \V4/V3/V1/V3/HA2/_0_  (.A1(\V4/V3/V1/V3/w4 ),
    .A2(\V4/V3/V1/V3/w3 ),
    .ZN(\V4/V3/V1/v3 [3]));
 XOR2_X2 \V4/V3/V1/V3/HA2/_1_  (.A(\V4/V3/V1/V3/w4 ),
    .B(\V4/V3/V1/V3/w3 ),
    .Z(\V4/V3/V1/v3 [2]));
 AND2_X1 \V4/V3/V1/V3/_0_  (.A1(net41),
    .A2(net13),
    .ZN(\V4/V3/V1/v3 [0]));
 AND2_X1 \V4/V3/V1/V3/_1_  (.A1(net41),
    .A2(B[27]),
    .ZN(\V4/V3/V1/V3/w1 ));
 AND2_X1 \V4/V3/V1/V3/_2_  (.A1(net13),
    .A2(net40),
    .ZN(\V4/V3/V1/V3/w2 ));
 AND2_X1 \V4/V3/V1/V3/_3_  (.A1(B[27]),
    .A2(net40),
    .ZN(\V4/V3/V1/V3/w3 ));
 AND2_X1 \V4/V3/V1/V4/HA1/_0_  (.A1(\V4/V3/V1/V4/w2 ),
    .A2(\V4/V3/V1/V4/w1 ),
    .ZN(\V4/V3/V1/V4/w4 ));
 XOR2_X2 \V4/V3/V1/V4/HA1/_1_  (.A(\V4/V3/V1/V4/w2 ),
    .B(\V4/V3/V1/V4/w1 ),
    .Z(\V4/V3/V1/v4 [1]));
 AND2_X1 \V4/V3/V1/V4/HA2/_0_  (.A1(\V4/V3/V1/V4/w4 ),
    .A2(\V4/V3/V1/V4/w3 ),
    .ZN(\V4/V3/V1/v4 [3]));
 XOR2_X2 \V4/V3/V1/V4/HA2/_1_  (.A(\V4/V3/V1/V4/w4 ),
    .B(\V4/V3/V1/V4/w3 ),
    .Z(\V4/V3/V1/v4 [2]));
 AND2_X1 \V4/V3/V1/V4/_0_  (.A1(net39),
    .A2(net13),
    .ZN(\V4/V3/V1/v4 [0]));
 AND2_X1 \V4/V3/V1/V4/_1_  (.A1(net39),
    .A2(B[27]),
    .ZN(\V4/V3/V1/V4/w1 ));
 AND2_X1 \V4/V3/V1/V4/_2_  (.A1(net13),
    .A2(net38),
    .ZN(\V4/V3/V1/V4/w2 ));
 AND2_X1 \V4/V3/V1/V4/_3_  (.A1(B[27]),
    .A2(net38),
    .ZN(\V4/V3/V1/V4/w3 ));
 OR2_X1 \V4/V3/V1/_0_  (.A1(\V4/V3/V1/c1 ),
    .A2(\V4/V3/V1/c2 ),
    .ZN(\V4/V3/V1/c3 ));
 AND2_X1 \V4/V3/V2/A1/M1/M1/_0_  (.A1(\V4/V3/V2/v2 [0]),
    .A2(\V4/V3/V2/v3 [0]),
    .ZN(\V4/V3/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M1/M1/_1_  (.A(\V4/V3/V2/v2 [0]),
    .B(\V4/V3/V2/v3 [0]),
    .Z(\V4/V3/V2/A1/M1/s1 ));
 AND2_X1 \V4/V3/V2/A1/M1/M2/_0_  (.A1(\V4/V3/V2/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V3/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M1/M2/_1_  (.A(\V4/V3/V2/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/V3/V2/s1 [0]));
 OR2_X1 \V4/V3/V2/A1/M1/_0_  (.A1(\V4/V3/V2/A1/M1/c1 ),
    .A2(\V4/V3/V2/A1/M1/c2 ),
    .ZN(\V4/V3/V2/A1/c1 ));
 AND2_X1 \V4/V3/V2/A1/M2/M1/_0_  (.A1(\V4/V3/V2/v2 [1]),
    .A2(\V4/V3/V2/v3 [1]),
    .ZN(\V4/V3/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M2/M1/_1_  (.A(\V4/V3/V2/v2 [1]),
    .B(\V4/V3/V2/v3 [1]),
    .Z(\V4/V3/V2/A1/M2/s1 ));
 AND2_X1 \V4/V3/V2/A1/M2/M2/_0_  (.A1(\V4/V3/V2/A1/M2/s1 ),
    .A2(\V4/V3/V2/A1/c1 ),
    .ZN(\V4/V3/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M2/M2/_1_  (.A(\V4/V3/V2/A1/M2/s1 ),
    .B(\V4/V3/V2/A1/c1 ),
    .Z(\V4/V3/V2/s1 [1]));
 OR2_X1 \V4/V3/V2/A1/M2/_0_  (.A1(\V4/V3/V2/A1/M2/c1 ),
    .A2(\V4/V3/V2/A1/M2/c2 ),
    .ZN(\V4/V3/V2/A1/c2 ));
 AND2_X1 \V4/V3/V2/A1/M3/M1/_0_  (.A1(\V4/V3/V2/v2 [2]),
    .A2(\V4/V3/V2/v3 [2]),
    .ZN(\V4/V3/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M3/M1/_1_  (.A(\V4/V3/V2/v2 [2]),
    .B(\V4/V3/V2/v3 [2]),
    .Z(\V4/V3/V2/A1/M3/s1 ));
 AND2_X1 \V4/V3/V2/A1/M3/M2/_0_  (.A1(\V4/V3/V2/A1/M3/s1 ),
    .A2(\V4/V3/V2/A1/c2 ),
    .ZN(\V4/V3/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M3/M2/_1_  (.A(\V4/V3/V2/A1/M3/s1 ),
    .B(\V4/V3/V2/A1/c2 ),
    .Z(\V4/V3/V2/s1 [2]));
 OR2_X1 \V4/V3/V2/A1/M3/_0_  (.A1(\V4/V3/V2/A1/M3/c1 ),
    .A2(\V4/V3/V2/A1/M3/c2 ),
    .ZN(\V4/V3/V2/A1/c3 ));
 AND2_X1 \V4/V3/V2/A1/M4/M1/_0_  (.A1(\V4/V3/V2/v2 [3]),
    .A2(\V4/V3/V2/v3 [3]),
    .ZN(\V4/V3/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A1/M4/M1/_1_  (.A(\V4/V3/V2/v2 [3]),
    .B(\V4/V3/V2/v3 [3]),
    .Z(\V4/V3/V2/A1/M4/s1 ));
 AND2_X1 \V4/V3/V2/A1/M4/M2/_0_  (.A1(\V4/V3/V2/A1/M4/s1 ),
    .A2(\V4/V3/V2/A1/c3 ),
    .ZN(\V4/V3/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A1/M4/M2/_1_  (.A(\V4/V3/V2/A1/M4/s1 ),
    .B(\V4/V3/V2/A1/c3 ),
    .Z(\V4/V3/V2/s1 [3]));
 OR2_X1 \V4/V3/V2/A1/M4/_0_  (.A1(\V4/V3/V2/A1/M4/c1 ),
    .A2(\V4/V3/V2/A1/M4/c2 ),
    .ZN(\V4/V3/V2/c1 ));
 AND2_X1 \V4/V3/V2/A2/M1/M1/_0_  (.A1(\V4/V3/V2/s1 [0]),
    .A2(\V4/V3/V2/v1 [2]),
    .ZN(\V4/V3/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M1/M1/_1_  (.A(\V4/V3/V2/s1 [0]),
    .B(\V4/V3/V2/v1 [2]),
    .Z(\V4/V3/V2/A2/M1/s1 ));
 AND2_X1 \V4/V3/V2/A2/M1/M2/_0_  (.A1(\V4/V3/V2/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M1/M2/_1_  (.A(\V4/V3/V2/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v2 [2]));
 OR2_X1 \V4/V3/V2/A2/M1/_0_  (.A1(\V4/V3/V2/A2/M1/c1 ),
    .A2(\V4/V3/V2/A2/M1/c2 ),
    .ZN(\V4/V3/V2/A2/c1 ));
 AND2_X1 \V4/V3/V2/A2/M2/M1/_0_  (.A1(\V4/V3/V2/s1 [1]),
    .A2(\V4/V3/V2/v1 [3]),
    .ZN(\V4/V3/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M2/M1/_1_  (.A(\V4/V3/V2/s1 [1]),
    .B(\V4/V3/V2/v1 [3]),
    .Z(\V4/V3/V2/A2/M2/s1 ));
 AND2_X1 \V4/V3/V2/A2/M2/M2/_0_  (.A1(\V4/V3/V2/A2/M2/s1 ),
    .A2(\V4/V3/V2/A2/c1 ),
    .ZN(\V4/V3/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M2/M2/_1_  (.A(\V4/V3/V2/A2/M2/s1 ),
    .B(\V4/V3/V2/A2/c1 ),
    .Z(\V4/V3/v2 [3]));
 OR2_X1 \V4/V3/V2/A2/M2/_0_  (.A1(\V4/V3/V2/A2/M2/c1 ),
    .A2(\V4/V3/V2/A2/M2/c2 ),
    .ZN(\V4/V3/V2/A2/c2 ));
 AND2_X1 \V4/V3/V2/A2/M3/M1/_0_  (.A1(\V4/V3/V2/s1 [2]),
    .A2(net9),
    .ZN(\V4/V3/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M3/M1/_1_  (.A(\V4/V3/V2/s1 [2]),
    .B(net9),
    .Z(\V4/V3/V2/A2/M3/s1 ));
 AND2_X1 \V4/V3/V2/A2/M3/M2/_0_  (.A1(\V4/V3/V2/A2/M3/s1 ),
    .A2(\V4/V3/V2/A2/c2 ),
    .ZN(\V4/V3/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M3/M2/_1_  (.A(\V4/V3/V2/A2/M3/s1 ),
    .B(\V4/V3/V2/A2/c2 ),
    .Z(\V4/V3/V2/s2 [2]));
 OR2_X1 \V4/V3/V2/A2/M3/_0_  (.A1(\V4/V3/V2/A2/M3/c1 ),
    .A2(\V4/V3/V2/A2/M3/c2 ),
    .ZN(\V4/V3/V2/A2/c3 ));
 AND2_X1 \V4/V3/V2/A2/M4/M1/_0_  (.A1(\V4/V3/V2/s1 [3]),
    .A2(net8),
    .ZN(\V4/V3/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A2/M4/M1/_1_  (.A(\V4/V3/V2/s1 [3]),
    .B(net8),
    .Z(\V4/V3/V2/A2/M4/s1 ));
 AND2_X1 \V4/V3/V2/A2/M4/M2/_0_  (.A1(\V4/V3/V2/A2/M4/s1 ),
    .A2(\V4/V3/V2/A2/c3 ),
    .ZN(\V4/V3/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A2/M4/M2/_1_  (.A(\V4/V3/V2/A2/M4/s1 ),
    .B(\V4/V3/V2/A2/c3 ),
    .Z(\V4/V3/V2/s2 [3]));
 OR2_X1 \V4/V3/V2/A2/M4/_0_  (.A1(\V4/V3/V2/A2/M4/c1 ),
    .A2(\V4/V3/V2/A2/M4/c2 ),
    .ZN(\V4/V3/V2/c2 ));
 AND2_X1 \V4/V3/V2/A3/M1/M1/_0_  (.A1(\V4/V3/V2/v4 [0]),
    .A2(\V4/V3/V2/s2 [2]),
    .ZN(\V4/V3/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M1/M1/_1_  (.A(\V4/V3/V2/v4 [0]),
    .B(\V4/V3/V2/s2 [2]),
    .Z(\V4/V3/V2/A3/M1/s1 ));
 AND2_X1 \V4/V3/V2/A3/M1/M2/_0_  (.A1(\V4/V3/V2/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V3/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M1/M2/_1_  (.A(\V4/V3/V2/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v2 [4]));
 OR2_X1 \V4/V3/V2/A3/M1/_0_  (.A1(\V4/V3/V2/A3/M1/c1 ),
    .A2(\V4/V3/V2/A3/M1/c2 ),
    .ZN(\V4/V3/V2/A3/c1 ));
 AND2_X1 \V4/V3/V2/A3/M2/M1/_0_  (.A1(\V4/V3/V2/v4 [1]),
    .A2(\V4/V3/V2/s2 [3]),
    .ZN(\V4/V3/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M2/M1/_1_  (.A(\V4/V3/V2/v4 [1]),
    .B(\V4/V3/V2/s2 [3]),
    .Z(\V4/V3/V2/A3/M2/s1 ));
 AND2_X1 \V4/V3/V2/A3/M2/M2/_0_  (.A1(\V4/V3/V2/A3/M2/s1 ),
    .A2(\V4/V3/V2/A3/c1 ),
    .ZN(\V4/V3/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M2/M2/_1_  (.A(\V4/V3/V2/A3/M2/s1 ),
    .B(\V4/V3/V2/A3/c1 ),
    .Z(\V4/V3/v2 [5]));
 OR2_X1 \V4/V3/V2/A3/M2/_0_  (.A1(\V4/V3/V2/A3/M2/c1 ),
    .A2(\V4/V3/V2/A3/M2/c2 ),
    .ZN(\V4/V3/V2/A3/c2 ));
 AND2_X1 \V4/V3/V2/A3/M3/M1/_0_  (.A1(\V4/V3/V2/v4 [2]),
    .A2(\V4/V3/V2/c3 ),
    .ZN(\V4/V3/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M3/M1/_1_  (.A(\V4/V3/V2/v4 [2]),
    .B(\V4/V3/V2/c3 ),
    .Z(\V4/V3/V2/A3/M3/s1 ));
 AND2_X1 \V4/V3/V2/A3/M3/M2/_0_  (.A1(\V4/V3/V2/A3/M3/s1 ),
    .A2(\V4/V3/V2/A3/c2 ),
    .ZN(\V4/V3/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M3/M2/_1_  (.A(\V4/V3/V2/A3/M3/s1 ),
    .B(\V4/V3/V2/A3/c2 ),
    .Z(\V4/V3/v2 [6]));
 OR2_X1 \V4/V3/V2/A3/M3/_0_  (.A1(\V4/V3/V2/A3/M3/c1 ),
    .A2(\V4/V3/V2/A3/M3/c2 ),
    .ZN(\V4/V3/V2/A3/c3 ));
 AND2_X1 \V4/V3/V2/A3/M4/M1/_0_  (.A1(\V4/V3/V2/v4 [3]),
    .A2(net9),
    .ZN(\V4/V3/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V2/A3/M4/M1/_1_  (.A(\V4/V3/V2/v4 [3]),
    .B(net9),
    .Z(\V4/V3/V2/A3/M4/s1 ));
 AND2_X1 \V4/V3/V2/A3/M4/M2/_0_  (.A1(\V4/V3/V2/A3/M4/s1 ),
    .A2(\V4/V3/V2/A3/c3 ),
    .ZN(\V4/V3/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V2/A3/M4/M2/_1_  (.A(\V4/V3/V2/A3/M4/s1 ),
    .B(\V4/V3/V2/A3/c3 ),
    .Z(\V4/V3/v2 [7]));
 OR2_X1 \V4/V3/V2/A3/M4/_0_  (.A1(\V4/V3/V2/A3/M4/c1 ),
    .A2(\V4/V3/V2/A3/M4/c2 ),
    .ZN(\V4/V3/V2/overflow ));
 AND2_X1 \V4/V3/V2/V1/HA1/_0_  (.A1(\V4/V3/V2/V1/w2 ),
    .A2(\V4/V3/V2/V1/w1 ),
    .ZN(\V4/V3/V2/V1/w4 ));
 XOR2_X2 \V4/V3/V2/V1/HA1/_1_  (.A(\V4/V3/V2/V1/w2 ),
    .B(\V4/V3/V2/V1/w1 ),
    .Z(\V4/V3/v2 [1]));
 AND2_X1 \V4/V3/V2/V1/HA2/_0_  (.A1(\V4/V3/V2/V1/w4 ),
    .A2(\V4/V3/V2/V1/w3 ),
    .ZN(\V4/V3/V2/v1 [3]));
 XOR2_X2 \V4/V3/V2/V1/HA2/_1_  (.A(\V4/V3/V2/V1/w4 ),
    .B(\V4/V3/V2/V1/w3 ),
    .Z(\V4/V3/V2/v1 [2]));
 AND2_X1 \V4/V3/V2/V1/_0_  (.A1(net37),
    .A2(net14),
    .ZN(\V4/V3/v2 [0]));
 AND2_X1 \V4/V3/V2/V1/_1_  (.A1(net37),
    .A2(B[25]),
    .ZN(\V4/V3/V2/V1/w1 ));
 AND2_X1 \V4/V3/V2/V1/_2_  (.A1(net14),
    .A2(net36),
    .ZN(\V4/V3/V2/V1/w2 ));
 AND2_X1 \V4/V3/V2/V1/_3_  (.A1(B[25]),
    .A2(net36),
    .ZN(\V4/V3/V2/V1/w3 ));
 AND2_X1 \V4/V3/V2/V2/HA1/_0_  (.A1(\V4/V3/V2/V2/w2 ),
    .A2(\V4/V3/V2/V2/w1 ),
    .ZN(\V4/V3/V2/V2/w4 ));
 XOR2_X2 \V4/V3/V2/V2/HA1/_1_  (.A(\V4/V3/V2/V2/w2 ),
    .B(\V4/V3/V2/V2/w1 ),
    .Z(\V4/V3/V2/v2 [1]));
 AND2_X1 \V4/V3/V2/V2/HA2/_0_  (.A1(\V4/V3/V2/V2/w4 ),
    .A2(\V4/V3/V2/V2/w3 ),
    .ZN(\V4/V3/V2/v2 [3]));
 XOR2_X2 \V4/V3/V2/V2/HA2/_1_  (.A(\V4/V3/V2/V2/w4 ),
    .B(\V4/V3/V2/V2/w3 ),
    .Z(\V4/V3/V2/v2 [2]));
 AND2_X1 \V4/V3/V2/V2/_0_  (.A1(net35),
    .A2(net14),
    .ZN(\V4/V3/V2/v2 [0]));
 AND2_X1 \V4/V3/V2/V2/_1_  (.A1(net35),
    .A2(B[25]),
    .ZN(\V4/V3/V2/V2/w1 ));
 AND2_X1 \V4/V3/V2/V2/_2_  (.A1(net14),
    .A2(net34),
    .ZN(\V4/V3/V2/V2/w2 ));
 AND2_X1 \V4/V3/V2/V2/_3_  (.A1(B[25]),
    .A2(net34),
    .ZN(\V4/V3/V2/V2/w3 ));
 AND2_X1 \V4/V3/V2/V3/HA1/_0_  (.A1(\V4/V3/V2/V3/w2 ),
    .A2(\V4/V3/V2/V3/w1 ),
    .ZN(\V4/V3/V2/V3/w4 ));
 XOR2_X2 \V4/V3/V2/V3/HA1/_1_  (.A(\V4/V3/V2/V3/w2 ),
    .B(\V4/V3/V2/V3/w1 ),
    .Z(\V4/V3/V2/v3 [1]));
 AND2_X1 \V4/V3/V2/V3/HA2/_0_  (.A1(\V4/V3/V2/V3/w4 ),
    .A2(\V4/V3/V2/V3/w3 ),
    .ZN(\V4/V3/V2/v3 [3]));
 XOR2_X2 \V4/V3/V2/V3/HA2/_1_  (.A(\V4/V3/V2/V3/w4 ),
    .B(\V4/V3/V2/V3/w3 ),
    .Z(\V4/V3/V2/v3 [2]));
 AND2_X1 \V4/V3/V2/V3/_0_  (.A1(net37),
    .A2(net13),
    .ZN(\V4/V3/V2/v3 [0]));
 AND2_X1 \V4/V3/V2/V3/_1_  (.A1(net37),
    .A2(B[27]),
    .ZN(\V4/V3/V2/V3/w1 ));
 AND2_X1 \V4/V3/V2/V3/_2_  (.A1(net13),
    .A2(net36),
    .ZN(\V4/V3/V2/V3/w2 ));
 AND2_X1 \V4/V3/V2/V3/_3_  (.A1(B[27]),
    .A2(net36),
    .ZN(\V4/V3/V2/V3/w3 ));
 AND2_X1 \V4/V3/V2/V4/HA1/_0_  (.A1(\V4/V3/V2/V4/w2 ),
    .A2(\V4/V3/V2/V4/w1 ),
    .ZN(\V4/V3/V2/V4/w4 ));
 XOR2_X2 \V4/V3/V2/V4/HA1/_1_  (.A(\V4/V3/V2/V4/w2 ),
    .B(\V4/V3/V2/V4/w1 ),
    .Z(\V4/V3/V2/v4 [1]));
 AND2_X1 \V4/V3/V2/V4/HA2/_0_  (.A1(\V4/V3/V2/V4/w4 ),
    .A2(\V4/V3/V2/V4/w3 ),
    .ZN(\V4/V3/V2/v4 [3]));
 XOR2_X2 \V4/V3/V2/V4/HA2/_1_  (.A(\V4/V3/V2/V4/w4 ),
    .B(\V4/V3/V2/V4/w3 ),
    .Z(\V4/V3/V2/v4 [2]));
 AND2_X1 \V4/V3/V2/V4/_0_  (.A1(net35),
    .A2(net13),
    .ZN(\V4/V3/V2/v4 [0]));
 AND2_X1 \V4/V3/V2/V4/_1_  (.A1(net35),
    .A2(B[27]),
    .ZN(\V4/V3/V2/V4/w1 ));
 AND2_X1 \V4/V3/V2/V4/_2_  (.A1(net13),
    .A2(net34),
    .ZN(\V4/V3/V2/V4/w2 ));
 AND2_X1 \V4/V3/V2/V4/_3_  (.A1(B[27]),
    .A2(net34),
    .ZN(\V4/V3/V2/V4/w3 ));
 OR2_X1 \V4/V3/V2/_0_  (.A1(\V4/V3/V2/c1 ),
    .A2(\V4/V3/V2/c2 ),
    .ZN(\V4/V3/V2/c3 ));
 AND2_X1 \V4/V3/V3/A1/M1/M1/_0_  (.A1(\V4/V3/V3/v2 [0]),
    .A2(\V4/V3/V3/v3 [0]),
    .ZN(\V4/V3/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M1/M1/_1_  (.A(\V4/V3/V3/v2 [0]),
    .B(\V4/V3/V3/v3 [0]),
    .Z(\V4/V3/V3/A1/M1/s1 ));
 AND2_X1 \V4/V3/V3/A1/M1/M2/_0_  (.A1(\V4/V3/V3/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M1/M2/_1_  (.A(\V4/V3/V3/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/V3/s1 [0]));
 OR2_X1 \V4/V3/V3/A1/M1/_0_  (.A1(\V4/V3/V3/A1/M1/c1 ),
    .A2(\V4/V3/V3/A1/M1/c2 ),
    .ZN(\V4/V3/V3/A1/c1 ));
 AND2_X1 \V4/V3/V3/A1/M2/M1/_0_  (.A1(\V4/V3/V3/v2 [1]),
    .A2(\V4/V3/V3/v3 [1]),
    .ZN(\V4/V3/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M2/M1/_1_  (.A(\V4/V3/V3/v2 [1]),
    .B(\V4/V3/V3/v3 [1]),
    .Z(\V4/V3/V3/A1/M2/s1 ));
 AND2_X1 \V4/V3/V3/A1/M2/M2/_0_  (.A1(\V4/V3/V3/A1/M2/s1 ),
    .A2(\V4/V3/V3/A1/c1 ),
    .ZN(\V4/V3/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M2/M2/_1_  (.A(\V4/V3/V3/A1/M2/s1 ),
    .B(\V4/V3/V3/A1/c1 ),
    .Z(\V4/V3/V3/s1 [1]));
 OR2_X1 \V4/V3/V3/A1/M2/_0_  (.A1(\V4/V3/V3/A1/M2/c1 ),
    .A2(\V4/V3/V3/A1/M2/c2 ),
    .ZN(\V4/V3/V3/A1/c2 ));
 AND2_X1 \V4/V3/V3/A1/M3/M1/_0_  (.A1(\V4/V3/V3/v2 [2]),
    .A2(\V4/V3/V3/v3 [2]),
    .ZN(\V4/V3/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M3/M1/_1_  (.A(\V4/V3/V3/v2 [2]),
    .B(\V4/V3/V3/v3 [2]),
    .Z(\V4/V3/V3/A1/M3/s1 ));
 AND2_X1 \V4/V3/V3/A1/M3/M2/_0_  (.A1(\V4/V3/V3/A1/M3/s1 ),
    .A2(\V4/V3/V3/A1/c2 ),
    .ZN(\V4/V3/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M3/M2/_1_  (.A(\V4/V3/V3/A1/M3/s1 ),
    .B(\V4/V3/V3/A1/c2 ),
    .Z(\V4/V3/V3/s1 [2]));
 OR2_X1 \V4/V3/V3/A1/M3/_0_  (.A1(\V4/V3/V3/A1/M3/c1 ),
    .A2(\V4/V3/V3/A1/M3/c2 ),
    .ZN(\V4/V3/V3/A1/c3 ));
 AND2_X1 \V4/V3/V3/A1/M4/M1/_0_  (.A1(\V4/V3/V3/v2 [3]),
    .A2(\V4/V3/V3/v3 [3]),
    .ZN(\V4/V3/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A1/M4/M1/_1_  (.A(\V4/V3/V3/v2 [3]),
    .B(\V4/V3/V3/v3 [3]),
    .Z(\V4/V3/V3/A1/M4/s1 ));
 AND2_X1 \V4/V3/V3/A1/M4/M2/_0_  (.A1(\V4/V3/V3/A1/M4/s1 ),
    .A2(\V4/V3/V3/A1/c3 ),
    .ZN(\V4/V3/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A1/M4/M2/_1_  (.A(\V4/V3/V3/A1/M4/s1 ),
    .B(\V4/V3/V3/A1/c3 ),
    .Z(\V4/V3/V3/s1 [3]));
 OR2_X1 \V4/V3/V3/A1/M4/_0_  (.A1(\V4/V3/V3/A1/M4/c1 ),
    .A2(\V4/V3/V3/A1/M4/c2 ),
    .ZN(\V4/V3/V3/c1 ));
 AND2_X1 \V4/V3/V3/A2/M1/M1/_0_  (.A1(\V4/V3/V3/s1 [0]),
    .A2(\V4/V3/V3/v1 [2]),
    .ZN(\V4/V3/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M1/M1/_1_  (.A(\V4/V3/V3/s1 [0]),
    .B(\V4/V3/V3/v1 [2]),
    .Z(\V4/V3/V3/A2/M1/s1 ));
 AND2_X1 \V4/V3/V3/A2/M1/M2/_0_  (.A1(\V4/V3/V3/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M1/M2/_1_  (.A(\V4/V3/V3/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v3 [2]));
 OR2_X1 \V4/V3/V3/A2/M1/_0_  (.A1(\V4/V3/V3/A2/M1/c1 ),
    .A2(\V4/V3/V3/A2/M1/c2 ),
    .ZN(\V4/V3/V3/A2/c1 ));
 AND2_X1 \V4/V3/V3/A2/M2/M1/_0_  (.A1(\V4/V3/V3/s1 [1]),
    .A2(\V4/V3/V3/v1 [3]),
    .ZN(\V4/V3/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M2/M1/_1_  (.A(\V4/V3/V3/s1 [1]),
    .B(\V4/V3/V3/v1 [3]),
    .Z(\V4/V3/V3/A2/M2/s1 ));
 AND2_X1 \V4/V3/V3/A2/M2/M2/_0_  (.A1(\V4/V3/V3/A2/M2/s1 ),
    .A2(\V4/V3/V3/A2/c1 ),
    .ZN(\V4/V3/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M2/M2/_1_  (.A(\V4/V3/V3/A2/M2/s1 ),
    .B(\V4/V3/V3/A2/c1 ),
    .Z(\V4/V3/v3 [3]));
 OR2_X1 \V4/V3/V3/A2/M2/_0_  (.A1(\V4/V3/V3/A2/M2/c1 ),
    .A2(\V4/V3/V3/A2/M2/c2 ),
    .ZN(\V4/V3/V3/A2/c2 ));
 AND2_X1 \V4/V3/V3/A2/M3/M1/_0_  (.A1(\V4/V3/V3/s1 [2]),
    .A2(net10),
    .ZN(\V4/V3/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M3/M1/_1_  (.A(\V4/V3/V3/s1 [2]),
    .B(net10),
    .Z(\V4/V3/V3/A2/M3/s1 ));
 AND2_X1 \V4/V3/V3/A2/M3/M2/_0_  (.A1(\V4/V3/V3/A2/M3/s1 ),
    .A2(\V4/V3/V3/A2/c2 ),
    .ZN(\V4/V3/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M3/M2/_1_  (.A(\V4/V3/V3/A2/M3/s1 ),
    .B(\V4/V3/V3/A2/c2 ),
    .Z(\V4/V3/V3/s2 [2]));
 OR2_X1 \V4/V3/V3/A2/M3/_0_  (.A1(\V4/V3/V3/A2/M3/c1 ),
    .A2(\V4/V3/V3/A2/M3/c2 ),
    .ZN(\V4/V3/V3/A2/c3 ));
 AND2_X1 \V4/V3/V3/A2/M4/M1/_0_  (.A1(\V4/V3/V3/s1 [3]),
    .A2(net9),
    .ZN(\V4/V3/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A2/M4/M1/_1_  (.A(\V4/V3/V3/s1 [3]),
    .B(net9),
    .Z(\V4/V3/V3/A2/M4/s1 ));
 AND2_X1 \V4/V3/V3/A2/M4/M2/_0_  (.A1(\V4/V3/V3/A2/M4/s1 ),
    .A2(\V4/V3/V3/A2/c3 ),
    .ZN(\V4/V3/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A2/M4/M2/_1_  (.A(\V4/V3/V3/A2/M4/s1 ),
    .B(\V4/V3/V3/A2/c3 ),
    .Z(\V4/V3/V3/s2 [3]));
 OR2_X1 \V4/V3/V3/A2/M4/_0_  (.A1(\V4/V3/V3/A2/M4/c1 ),
    .A2(\V4/V3/V3/A2/M4/c2 ),
    .ZN(\V4/V3/V3/c2 ));
 AND2_X1 \V4/V3/V3/A3/M1/M1/_0_  (.A1(\V4/V3/V3/v4 [0]),
    .A2(\V4/V3/V3/s2 [2]),
    .ZN(\V4/V3/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M1/M1/_1_  (.A(\V4/V3/V3/v4 [0]),
    .B(\V4/V3/V3/s2 [2]),
    .Z(\V4/V3/V3/A3/M1/s1 ));
 AND2_X1 \V4/V3/V3/A3/M1/M2/_0_  (.A1(\V4/V3/V3/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V3/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M1/M2/_1_  (.A(\V4/V3/V3/A3/M1/s1 ),
    .B(net9),
    .Z(\V4/V3/v3 [4]));
 OR2_X1 \V4/V3/V3/A3/M1/_0_  (.A1(\V4/V3/V3/A3/M1/c1 ),
    .A2(\V4/V3/V3/A3/M1/c2 ),
    .ZN(\V4/V3/V3/A3/c1 ));
 AND2_X1 \V4/V3/V3/A3/M2/M1/_0_  (.A1(\V4/V3/V3/v4 [1]),
    .A2(\V4/V3/V3/s2 [3]),
    .ZN(\V4/V3/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M2/M1/_1_  (.A(\V4/V3/V3/v4 [1]),
    .B(\V4/V3/V3/s2 [3]),
    .Z(\V4/V3/V3/A3/M2/s1 ));
 AND2_X1 \V4/V3/V3/A3/M2/M2/_0_  (.A1(\V4/V3/V3/A3/M2/s1 ),
    .A2(\V4/V3/V3/A3/c1 ),
    .ZN(\V4/V3/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M2/M2/_1_  (.A(\V4/V3/V3/A3/M2/s1 ),
    .B(\V4/V3/V3/A3/c1 ),
    .Z(\V4/V3/v3 [5]));
 OR2_X1 \V4/V3/V3/A3/M2/_0_  (.A1(\V4/V3/V3/A3/M2/c1 ),
    .A2(\V4/V3/V3/A3/M2/c2 ),
    .ZN(\V4/V3/V3/A3/c2 ));
 AND2_X1 \V4/V3/V3/A3/M3/M1/_0_  (.A1(\V4/V3/V3/v4 [2]),
    .A2(\V4/V3/V3/c3 ),
    .ZN(\V4/V3/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M3/M1/_1_  (.A(\V4/V3/V3/v4 [2]),
    .B(\V4/V3/V3/c3 ),
    .Z(\V4/V3/V3/A3/M3/s1 ));
 AND2_X1 \V4/V3/V3/A3/M3/M2/_0_  (.A1(\V4/V3/V3/A3/M3/s1 ),
    .A2(\V4/V3/V3/A3/c2 ),
    .ZN(\V4/V3/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M3/M2/_1_  (.A(\V4/V3/V3/A3/M3/s1 ),
    .B(\V4/V3/V3/A3/c2 ),
    .Z(\V4/V3/v3 [6]));
 OR2_X1 \V4/V3/V3/A3/M3/_0_  (.A1(\V4/V3/V3/A3/M3/c1 ),
    .A2(\V4/V3/V3/A3/M3/c2 ),
    .ZN(\V4/V3/V3/A3/c3 ));
 AND2_X1 \V4/V3/V3/A3/M4/M1/_0_  (.A1(\V4/V3/V3/v4 [3]),
    .A2(net7),
    .ZN(\V4/V3/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V3/A3/M4/M1/_1_  (.A(\V4/V3/V3/v4 [3]),
    .B(net7),
    .Z(\V4/V3/V3/A3/M4/s1 ));
 AND2_X1 \V4/V3/V3/A3/M4/M2/_0_  (.A1(\V4/V3/V3/A3/M4/s1 ),
    .A2(\V4/V3/V3/A3/c3 ),
    .ZN(\V4/V3/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V3/A3/M4/M2/_1_  (.A(\V4/V3/V3/A3/M4/s1 ),
    .B(\V4/V3/V3/A3/c3 ),
    .Z(\V4/V3/v3 [7]));
 OR2_X1 \V4/V3/V3/A3/M4/_0_  (.A1(\V4/V3/V3/A3/M4/c1 ),
    .A2(\V4/V3/V3/A3/M4/c2 ),
    .ZN(\V4/V3/V3/overflow ));
 AND2_X1 \V4/V3/V3/V1/HA1/_0_  (.A1(\V4/V3/V3/V1/w2 ),
    .A2(\V4/V3/V3/V1/w1 ),
    .ZN(\V4/V3/V3/V1/w4 ));
 XOR2_X2 \V4/V3/V3/V1/HA1/_1_  (.A(\V4/V3/V3/V1/w2 ),
    .B(\V4/V3/V3/V1/w1 ),
    .Z(\V4/V3/v3 [1]));
 AND2_X1 \V4/V3/V3/V1/HA2/_0_  (.A1(\V4/V3/V3/V1/w4 ),
    .A2(\V4/V3/V3/V1/w3 ),
    .ZN(\V4/V3/V3/v1 [3]));
 XOR2_X2 \V4/V3/V3/V1/HA2/_1_  (.A(\V4/V3/V3/V1/w4 ),
    .B(\V4/V3/V3/V1/w3 ),
    .Z(\V4/V3/V3/v1 [2]));
 AND2_X1 \V4/V3/V3/V1/_0_  (.A1(net41),
    .A2(B[28]),
    .ZN(\V4/V3/v3 [0]));
 AND2_X1 \V4/V3/V3/V1/_1_  (.A1(net41),
    .A2(B[29]),
    .ZN(\V4/V3/V3/V1/w1 ));
 AND2_X1 \V4/V3/V3/V1/_2_  (.A1(B[28]),
    .A2(net40),
    .ZN(\V4/V3/V3/V1/w2 ));
 AND2_X1 \V4/V3/V3/V1/_3_  (.A1(B[29]),
    .A2(net40),
    .ZN(\V4/V3/V3/V1/w3 ));
 AND2_X1 \V4/V3/V3/V2/HA1/_0_  (.A1(\V4/V3/V3/V2/w2 ),
    .A2(\V4/V3/V3/V2/w1 ),
    .ZN(\V4/V3/V3/V2/w4 ));
 XOR2_X2 \V4/V3/V3/V2/HA1/_1_  (.A(\V4/V3/V3/V2/w2 ),
    .B(\V4/V3/V3/V2/w1 ),
    .Z(\V4/V3/V3/v2 [1]));
 AND2_X1 \V4/V3/V3/V2/HA2/_0_  (.A1(\V4/V3/V3/V2/w4 ),
    .A2(\V4/V3/V3/V2/w3 ),
    .ZN(\V4/V3/V3/v2 [3]));
 XOR2_X2 \V4/V3/V3/V2/HA2/_1_  (.A(\V4/V3/V3/V2/w4 ),
    .B(\V4/V3/V3/V2/w3 ),
    .Z(\V4/V3/V3/v2 [2]));
 AND2_X1 \V4/V3/V3/V2/_0_  (.A1(net39),
    .A2(B[28]),
    .ZN(\V4/V3/V3/v2 [0]));
 AND2_X1 \V4/V3/V3/V2/_1_  (.A1(net39),
    .A2(B[29]),
    .ZN(\V4/V3/V3/V2/w1 ));
 AND2_X1 \V4/V3/V3/V2/_2_  (.A1(B[28]),
    .A2(net38),
    .ZN(\V4/V3/V3/V2/w2 ));
 AND2_X1 \V4/V3/V3/V2/_3_  (.A1(B[29]),
    .A2(net38),
    .ZN(\V4/V3/V3/V2/w3 ));
 AND2_X1 \V4/V3/V3/V3/HA1/_0_  (.A1(\V4/V3/V3/V3/w2 ),
    .A2(\V4/V3/V3/V3/w1 ),
    .ZN(\V4/V3/V3/V3/w4 ));
 XOR2_X2 \V4/V3/V3/V3/HA1/_1_  (.A(\V4/V3/V3/V3/w2 ),
    .B(\V4/V3/V3/V3/w1 ),
    .Z(\V4/V3/V3/v3 [1]));
 AND2_X1 \V4/V3/V3/V3/HA2/_0_  (.A1(\V4/V3/V3/V3/w4 ),
    .A2(\V4/V3/V3/V3/w3 ),
    .ZN(\V4/V3/V3/v3 [3]));
 XOR2_X2 \V4/V3/V3/V3/HA2/_1_  (.A(\V4/V3/V3/V3/w4 ),
    .B(\V4/V3/V3/V3/w3 ),
    .Z(\V4/V3/V3/v3 [2]));
 AND2_X1 \V4/V3/V3/V3/_0_  (.A1(net41),
    .A2(B[30]),
    .ZN(\V4/V3/V3/v3 [0]));
 AND2_X1 \V4/V3/V3/V3/_1_  (.A1(net41),
    .A2(B[31]),
    .ZN(\V4/V3/V3/V3/w1 ));
 AND2_X1 \V4/V3/V3/V3/_2_  (.A1(B[30]),
    .A2(net40),
    .ZN(\V4/V3/V3/V3/w2 ));
 AND2_X1 \V4/V3/V3/V3/_3_  (.A1(B[31]),
    .A2(net40),
    .ZN(\V4/V3/V3/V3/w3 ));
 AND2_X1 \V4/V3/V3/V4/HA1/_0_  (.A1(\V4/V3/V3/V4/w2 ),
    .A2(\V4/V3/V3/V4/w1 ),
    .ZN(\V4/V3/V3/V4/w4 ));
 XOR2_X2 \V4/V3/V3/V4/HA1/_1_  (.A(\V4/V3/V3/V4/w2 ),
    .B(\V4/V3/V3/V4/w1 ),
    .Z(\V4/V3/V3/v4 [1]));
 AND2_X1 \V4/V3/V3/V4/HA2/_0_  (.A1(\V4/V3/V3/V4/w4 ),
    .A2(\V4/V3/V3/V4/w3 ),
    .ZN(\V4/V3/V3/v4 [3]));
 XOR2_X2 \V4/V3/V3/V4/HA2/_1_  (.A(\V4/V3/V3/V4/w4 ),
    .B(\V4/V3/V3/V4/w3 ),
    .Z(\V4/V3/V3/v4 [2]));
 AND2_X1 \V4/V3/V3/V4/_0_  (.A1(net39),
    .A2(B[30]),
    .ZN(\V4/V3/V3/v4 [0]));
 AND2_X1 \V4/V3/V3/V4/_1_  (.A1(net39),
    .A2(B[31]),
    .ZN(\V4/V3/V3/V4/w1 ));
 AND2_X1 \V4/V3/V3/V4/_2_  (.A1(B[30]),
    .A2(net38),
    .ZN(\V4/V3/V3/V4/w2 ));
 AND2_X1 \V4/V3/V3/V4/_3_  (.A1(B[31]),
    .A2(net38),
    .ZN(\V4/V3/V3/V4/w3 ));
 OR2_X1 \V4/V3/V3/_0_  (.A1(\V4/V3/V3/c1 ),
    .A2(\V4/V3/V3/c2 ),
    .ZN(\V4/V3/V3/c3 ));
 AND2_X1 \V4/V3/V4/A1/M1/M1/_0_  (.A1(\V4/V3/V4/v2 [0]),
    .A2(\V4/V3/V4/v3 [0]),
    .ZN(\V4/V3/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M1/M1/_1_  (.A(\V4/V3/V4/v2 [0]),
    .B(\V4/V3/V4/v3 [0]),
    .Z(\V4/V3/V4/A1/M1/s1 ));
 AND2_X1 \V4/V3/V4/A1/M1/M2/_0_  (.A1(\V4/V3/V4/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M1/M2/_1_  (.A(\V4/V3/V4/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/V4/s1 [0]));
 OR2_X1 \V4/V3/V4/A1/M1/_0_  (.A1(\V4/V3/V4/A1/M1/c1 ),
    .A2(\V4/V3/V4/A1/M1/c2 ),
    .ZN(\V4/V3/V4/A1/c1 ));
 AND2_X1 \V4/V3/V4/A1/M2/M1/_0_  (.A1(\V4/V3/V4/v2 [1]),
    .A2(\V4/V3/V4/v3 [1]),
    .ZN(\V4/V3/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M2/M1/_1_  (.A(\V4/V3/V4/v2 [1]),
    .B(\V4/V3/V4/v3 [1]),
    .Z(\V4/V3/V4/A1/M2/s1 ));
 AND2_X1 \V4/V3/V4/A1/M2/M2/_0_  (.A1(\V4/V3/V4/A1/M2/s1 ),
    .A2(\V4/V3/V4/A1/c1 ),
    .ZN(\V4/V3/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M2/M2/_1_  (.A(\V4/V3/V4/A1/M2/s1 ),
    .B(\V4/V3/V4/A1/c1 ),
    .Z(\V4/V3/V4/s1 [1]));
 OR2_X1 \V4/V3/V4/A1/M2/_0_  (.A1(\V4/V3/V4/A1/M2/c1 ),
    .A2(\V4/V3/V4/A1/M2/c2 ),
    .ZN(\V4/V3/V4/A1/c2 ));
 AND2_X1 \V4/V3/V4/A1/M3/M1/_0_  (.A1(\V4/V3/V4/v2 [2]),
    .A2(\V4/V3/V4/v3 [2]),
    .ZN(\V4/V3/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M3/M1/_1_  (.A(\V4/V3/V4/v2 [2]),
    .B(\V4/V3/V4/v3 [2]),
    .Z(\V4/V3/V4/A1/M3/s1 ));
 AND2_X1 \V4/V3/V4/A1/M3/M2/_0_  (.A1(\V4/V3/V4/A1/M3/s1 ),
    .A2(\V4/V3/V4/A1/c2 ),
    .ZN(\V4/V3/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M3/M2/_1_  (.A(\V4/V3/V4/A1/M3/s1 ),
    .B(\V4/V3/V4/A1/c2 ),
    .Z(\V4/V3/V4/s1 [2]));
 OR2_X1 \V4/V3/V4/A1/M3/_0_  (.A1(\V4/V3/V4/A1/M3/c1 ),
    .A2(\V4/V3/V4/A1/M3/c2 ),
    .ZN(\V4/V3/V4/A1/c3 ));
 AND2_X1 \V4/V3/V4/A1/M4/M1/_0_  (.A1(\V4/V3/V4/v2 [3]),
    .A2(\V4/V3/V4/v3 [3]),
    .ZN(\V4/V3/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A1/M4/M1/_1_  (.A(\V4/V3/V4/v2 [3]),
    .B(\V4/V3/V4/v3 [3]),
    .Z(\V4/V3/V4/A1/M4/s1 ));
 AND2_X1 \V4/V3/V4/A1/M4/M2/_0_  (.A1(\V4/V3/V4/A1/M4/s1 ),
    .A2(\V4/V3/V4/A1/c3 ),
    .ZN(\V4/V3/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A1/M4/M2/_1_  (.A(\V4/V3/V4/A1/M4/s1 ),
    .B(\V4/V3/V4/A1/c3 ),
    .Z(\V4/V3/V4/s1 [3]));
 OR2_X1 \V4/V3/V4/A1/M4/_0_  (.A1(\V4/V3/V4/A1/M4/c1 ),
    .A2(\V4/V3/V4/A1/M4/c2 ),
    .ZN(\V4/V3/V4/c1 ));
 AND2_X1 \V4/V3/V4/A2/M1/M1/_0_  (.A1(\V4/V3/V4/s1 [0]),
    .A2(\V4/V3/V4/v1 [2]),
    .ZN(\V4/V3/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M1/M1/_1_  (.A(\V4/V3/V4/s1 [0]),
    .B(\V4/V3/V4/v1 [2]),
    .Z(\V4/V3/V4/A2/M1/s1 ));
 AND2_X1 \V4/V3/V4/A2/M1/M2/_0_  (.A1(\V4/V3/V4/A2/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M1/M2/_1_  (.A(\V4/V3/V4/A2/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v4 [2]));
 OR2_X1 \V4/V3/V4/A2/M1/_0_  (.A1(\V4/V3/V4/A2/M1/c1 ),
    .A2(\V4/V3/V4/A2/M1/c2 ),
    .ZN(\V4/V3/V4/A2/c1 ));
 AND2_X1 \V4/V3/V4/A2/M2/M1/_0_  (.A1(\V4/V3/V4/s1 [1]),
    .A2(\V4/V3/V4/v1 [3]),
    .ZN(\V4/V3/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M2/M1/_1_  (.A(\V4/V3/V4/s1 [1]),
    .B(\V4/V3/V4/v1 [3]),
    .Z(\V4/V3/V4/A2/M2/s1 ));
 AND2_X1 \V4/V3/V4/A2/M2/M2/_0_  (.A1(\V4/V3/V4/A2/M2/s1 ),
    .A2(\V4/V3/V4/A2/c1 ),
    .ZN(\V4/V3/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M2/M2/_1_  (.A(\V4/V3/V4/A2/M2/s1 ),
    .B(\V4/V3/V4/A2/c1 ),
    .Z(\V4/V3/v4 [3]));
 OR2_X1 \V4/V3/V4/A2/M2/_0_  (.A1(\V4/V3/V4/A2/M2/c1 ),
    .A2(\V4/V3/V4/A2/M2/c2 ),
    .ZN(\V4/V3/V4/A2/c2 ));
 AND2_X1 \V4/V3/V4/A2/M3/M1/_0_  (.A1(\V4/V3/V4/s1 [2]),
    .A2(net10),
    .ZN(\V4/V3/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M3/M1/_1_  (.A(\V4/V3/V4/s1 [2]),
    .B(net10),
    .Z(\V4/V3/V4/A2/M3/s1 ));
 AND2_X1 \V4/V3/V4/A2/M3/M2/_0_  (.A1(\V4/V3/V4/A2/M3/s1 ),
    .A2(\V4/V3/V4/A2/c2 ),
    .ZN(\V4/V3/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M3/M2/_1_  (.A(\V4/V3/V4/A2/M3/s1 ),
    .B(\V4/V3/V4/A2/c2 ),
    .Z(\V4/V3/V4/s2 [2]));
 OR2_X1 \V4/V3/V4/A2/M3/_0_  (.A1(\V4/V3/V4/A2/M3/c1 ),
    .A2(\V4/V3/V4/A2/M3/c2 ),
    .ZN(\V4/V3/V4/A2/c3 ));
 AND2_X1 \V4/V3/V4/A2/M4/M1/_0_  (.A1(\V4/V3/V4/s1 [3]),
    .A2(net9),
    .ZN(\V4/V3/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A2/M4/M1/_1_  (.A(\V4/V3/V4/s1 [3]),
    .B(net9),
    .Z(\V4/V3/V4/A2/M4/s1 ));
 AND2_X1 \V4/V3/V4/A2/M4/M2/_0_  (.A1(\V4/V3/V4/A2/M4/s1 ),
    .A2(\V4/V3/V4/A2/c3 ),
    .ZN(\V4/V3/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A2/M4/M2/_1_  (.A(\V4/V3/V4/A2/M4/s1 ),
    .B(\V4/V3/V4/A2/c3 ),
    .Z(\V4/V3/V4/s2 [3]));
 OR2_X1 \V4/V3/V4/A2/M4/_0_  (.A1(\V4/V3/V4/A2/M4/c1 ),
    .A2(\V4/V3/V4/A2/M4/c2 ),
    .ZN(\V4/V3/V4/c2 ));
 AND2_X1 \V4/V3/V4/A3/M1/M1/_0_  (.A1(\V4/V3/V4/v4 [0]),
    .A2(\V4/V3/V4/s2 [2]),
    .ZN(\V4/V3/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M1/M1/_1_  (.A(\V4/V3/V4/v4 [0]),
    .B(\V4/V3/V4/s2 [2]),
    .Z(\V4/V3/V4/A3/M1/s1 ));
 AND2_X1 \V4/V3/V4/A3/M1/M2/_0_  (.A1(\V4/V3/V4/A3/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V3/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M1/M2/_1_  (.A(\V4/V3/V4/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V3/v4 [4]));
 OR2_X1 \V4/V3/V4/A3/M1/_0_  (.A1(\V4/V3/V4/A3/M1/c1 ),
    .A2(\V4/V3/V4/A3/M1/c2 ),
    .ZN(\V4/V3/V4/A3/c1 ));
 AND2_X1 \V4/V3/V4/A3/M2/M1/_0_  (.A1(\V4/V3/V4/v4 [1]),
    .A2(\V4/V3/V4/s2 [3]),
    .ZN(\V4/V3/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M2/M1/_1_  (.A(\V4/V3/V4/v4 [1]),
    .B(\V4/V3/V4/s2 [3]),
    .Z(\V4/V3/V4/A3/M2/s1 ));
 AND2_X1 \V4/V3/V4/A3/M2/M2/_0_  (.A1(\V4/V3/V4/A3/M2/s1 ),
    .A2(\V4/V3/V4/A3/c1 ),
    .ZN(\V4/V3/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M2/M2/_1_  (.A(\V4/V3/V4/A3/M2/s1 ),
    .B(\V4/V3/V4/A3/c1 ),
    .Z(\V4/V3/v4 [5]));
 OR2_X1 \V4/V3/V4/A3/M2/_0_  (.A1(\V4/V3/V4/A3/M2/c1 ),
    .A2(\V4/V3/V4/A3/M2/c2 ),
    .ZN(\V4/V3/V4/A3/c2 ));
 AND2_X1 \V4/V3/V4/A3/M3/M1/_0_  (.A1(\V4/V3/V4/v4 [2]),
    .A2(\V4/V3/V4/c3 ),
    .ZN(\V4/V3/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M3/M1/_1_  (.A(\V4/V3/V4/v4 [2]),
    .B(\V4/V3/V4/c3 ),
    .Z(\V4/V3/V4/A3/M3/s1 ));
 AND2_X1 \V4/V3/V4/A3/M3/M2/_0_  (.A1(\V4/V3/V4/A3/M3/s1 ),
    .A2(\V4/V3/V4/A3/c2 ),
    .ZN(\V4/V3/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M3/M2/_1_  (.A(\V4/V3/V4/A3/M3/s1 ),
    .B(\V4/V3/V4/A3/c2 ),
    .Z(\V4/V3/v4 [6]));
 OR2_X1 \V4/V3/V4/A3/M3/_0_  (.A1(\V4/V3/V4/A3/M3/c1 ),
    .A2(\V4/V3/V4/A3/M3/c2 ),
    .ZN(\V4/V3/V4/A3/c3 ));
 AND2_X1 \V4/V3/V4/A3/M4/M1/_0_  (.A1(\V4/V3/V4/v4 [3]),
    .A2(net10),
    .ZN(\V4/V3/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V3/V4/A3/M4/M1/_1_  (.A(\V4/V3/V4/v4 [3]),
    .B(net10),
    .Z(\V4/V3/V4/A3/M4/s1 ));
 AND2_X1 \V4/V3/V4/A3/M4/M2/_0_  (.A1(\V4/V3/V4/A3/M4/s1 ),
    .A2(\V4/V3/V4/A3/c3 ),
    .ZN(\V4/V3/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V3/V4/A3/M4/M2/_1_  (.A(\V4/V3/V4/A3/M4/s1 ),
    .B(\V4/V3/V4/A3/c3 ),
    .Z(\V4/V3/v4 [7]));
 OR2_X1 \V4/V3/V4/A3/M4/_0_  (.A1(\V4/V3/V4/A3/M4/c1 ),
    .A2(\V4/V3/V4/A3/M4/c2 ),
    .ZN(\V4/V3/V4/overflow ));
 AND2_X1 \V4/V3/V4/V1/HA1/_0_  (.A1(\V4/V3/V4/V1/w2 ),
    .A2(\V4/V3/V4/V1/w1 ),
    .ZN(\V4/V3/V4/V1/w4 ));
 XOR2_X2 \V4/V3/V4/V1/HA1/_1_  (.A(\V4/V3/V4/V1/w2 ),
    .B(\V4/V3/V4/V1/w1 ),
    .Z(\V4/V3/v4 [1]));
 AND2_X1 \V4/V3/V4/V1/HA2/_0_  (.A1(\V4/V3/V4/V1/w4 ),
    .A2(\V4/V3/V4/V1/w3 ),
    .ZN(\V4/V3/V4/v1 [3]));
 XOR2_X2 \V4/V3/V4/V1/HA2/_1_  (.A(\V4/V3/V4/V1/w4 ),
    .B(\V4/V3/V4/V1/w3 ),
    .Z(\V4/V3/V4/v1 [2]));
 AND2_X1 \V4/V3/V4/V1/_0_  (.A1(net37),
    .A2(B[28]),
    .ZN(\V4/V3/v4 [0]));
 AND2_X1 \V4/V3/V4/V1/_1_  (.A1(net37),
    .A2(B[29]),
    .ZN(\V4/V3/V4/V1/w1 ));
 AND2_X1 \V4/V3/V4/V1/_2_  (.A1(B[28]),
    .A2(net36),
    .ZN(\V4/V3/V4/V1/w2 ));
 AND2_X1 \V4/V3/V4/V1/_3_  (.A1(B[29]),
    .A2(net36),
    .ZN(\V4/V3/V4/V1/w3 ));
 AND2_X1 \V4/V3/V4/V2/HA1/_0_  (.A1(\V4/V3/V4/V2/w2 ),
    .A2(\V4/V3/V4/V2/w1 ),
    .ZN(\V4/V3/V4/V2/w4 ));
 XOR2_X2 \V4/V3/V4/V2/HA1/_1_  (.A(\V4/V3/V4/V2/w2 ),
    .B(\V4/V3/V4/V2/w1 ),
    .Z(\V4/V3/V4/v2 [1]));
 AND2_X1 \V4/V3/V4/V2/HA2/_0_  (.A1(\V4/V3/V4/V2/w4 ),
    .A2(\V4/V3/V4/V2/w3 ),
    .ZN(\V4/V3/V4/v2 [3]));
 XOR2_X2 \V4/V3/V4/V2/HA2/_1_  (.A(\V4/V3/V4/V2/w4 ),
    .B(\V4/V3/V4/V2/w3 ),
    .Z(\V4/V3/V4/v2 [2]));
 AND2_X1 \V4/V3/V4/V2/_0_  (.A1(net35),
    .A2(B[28]),
    .ZN(\V4/V3/V4/v2 [0]));
 AND2_X1 \V4/V3/V4/V2/_1_  (.A1(net35),
    .A2(B[29]),
    .ZN(\V4/V3/V4/V2/w1 ));
 AND2_X1 \V4/V3/V4/V2/_2_  (.A1(B[28]),
    .A2(net34),
    .ZN(\V4/V3/V4/V2/w2 ));
 AND2_X1 \V4/V3/V4/V2/_3_  (.A1(B[29]),
    .A2(net34),
    .ZN(\V4/V3/V4/V2/w3 ));
 AND2_X1 \V4/V3/V4/V3/HA1/_0_  (.A1(\V4/V3/V4/V3/w2 ),
    .A2(\V4/V3/V4/V3/w1 ),
    .ZN(\V4/V3/V4/V3/w4 ));
 XOR2_X2 \V4/V3/V4/V3/HA1/_1_  (.A(\V4/V3/V4/V3/w2 ),
    .B(\V4/V3/V4/V3/w1 ),
    .Z(\V4/V3/V4/v3 [1]));
 AND2_X1 \V4/V3/V4/V3/HA2/_0_  (.A1(\V4/V3/V4/V3/w4 ),
    .A2(\V4/V3/V4/V3/w3 ),
    .ZN(\V4/V3/V4/v3 [3]));
 XOR2_X2 \V4/V3/V4/V3/HA2/_1_  (.A(\V4/V3/V4/V3/w4 ),
    .B(\V4/V3/V4/V3/w3 ),
    .Z(\V4/V3/V4/v3 [2]));
 AND2_X1 \V4/V3/V4/V3/_0_  (.A1(net37),
    .A2(B[30]),
    .ZN(\V4/V3/V4/v3 [0]));
 AND2_X1 \V4/V3/V4/V3/_1_  (.A1(net37),
    .A2(B[31]),
    .ZN(\V4/V3/V4/V3/w1 ));
 AND2_X1 \V4/V3/V4/V3/_2_  (.A1(B[30]),
    .A2(net36),
    .ZN(\V4/V3/V4/V3/w2 ));
 AND2_X1 \V4/V3/V4/V3/_3_  (.A1(B[31]),
    .A2(net36),
    .ZN(\V4/V3/V4/V3/w3 ));
 AND2_X1 \V4/V3/V4/V4/HA1/_0_  (.A1(\V4/V3/V4/V4/w2 ),
    .A2(\V4/V3/V4/V4/w1 ),
    .ZN(\V4/V3/V4/V4/w4 ));
 XOR2_X2 \V4/V3/V4/V4/HA1/_1_  (.A(\V4/V3/V4/V4/w2 ),
    .B(\V4/V3/V4/V4/w1 ),
    .Z(\V4/V3/V4/v4 [1]));
 AND2_X1 \V4/V3/V4/V4/HA2/_0_  (.A1(\V4/V3/V4/V4/w4 ),
    .A2(\V4/V3/V4/V4/w3 ),
    .ZN(\V4/V3/V4/v4 [3]));
 XOR2_X2 \V4/V3/V4/V4/HA2/_1_  (.A(\V4/V3/V4/V4/w4 ),
    .B(\V4/V3/V4/V4/w3 ),
    .Z(\V4/V3/V4/v4 [2]));
 AND2_X1 \V4/V3/V4/V4/_0_  (.A1(net35),
    .A2(B[30]),
    .ZN(\V4/V3/V4/v4 [0]));
 AND2_X1 \V4/V3/V4/V4/_1_  (.A1(net35),
    .A2(B[31]),
    .ZN(\V4/V3/V4/V4/w1 ));
 AND2_X1 \V4/V3/V4/V4/_2_  (.A1(B[30]),
    .A2(net34),
    .ZN(\V4/V3/V4/V4/w2 ));
 AND2_X1 \V4/V3/V4/V4/_3_  (.A1(B[31]),
    .A2(net34),
    .ZN(\V4/V3/V4/V4/w3 ));
 OR2_X1 \V4/V3/V4/_0_  (.A1(\V4/V3/V4/c1 ),
    .A2(\V4/V3/V4/c2 ),
    .ZN(\V4/V3/V4/c3 ));
 OR2_X1 \V4/V3/_0_  (.A1(\V4/V3/c1 ),
    .A2(\V4/V3/c2 ),
    .ZN(\V4/V3/c3 ));
 AND2_X1 \V4/V4/A1/A1/M1/M1/_0_  (.A1(\V4/V4/v2 [0]),
    .A2(\V4/V4/v3 [0]),
    .ZN(\V4/V4/A1/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M1/M1/_1_  (.A(\V4/V4/v2 [0]),
    .B(\V4/V4/v3 [0]),
    .Z(\V4/V4/A1/A1/M1/s1 ));
 AND2_X1 \V4/V4/A1/A1/M1/M2/_0_  (.A1(\V4/V4/A1/A1/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V4/A1/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M1/M2/_1_  (.A(\V4/V4/A1/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V4/s1 [0]));
 OR2_X1 \V4/V4/A1/A1/M1/_0_  (.A1(\V4/V4/A1/A1/M1/c1 ),
    .A2(\V4/V4/A1/A1/M1/c2 ),
    .ZN(\V4/V4/A1/A1/c1 ));
 AND2_X1 \V4/V4/A1/A1/M2/M1/_0_  (.A1(\V4/V4/v2 [1]),
    .A2(\V4/V4/v3 [1]),
    .ZN(\V4/V4/A1/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M2/M1/_1_  (.A(\V4/V4/v2 [1]),
    .B(\V4/V4/v3 [1]),
    .Z(\V4/V4/A1/A1/M2/s1 ));
 AND2_X1 \V4/V4/A1/A1/M2/M2/_0_  (.A1(\V4/V4/A1/A1/M2/s1 ),
    .A2(\V4/V4/A1/A1/c1 ),
    .ZN(\V4/V4/A1/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M2/M2/_1_  (.A(\V4/V4/A1/A1/M2/s1 ),
    .B(\V4/V4/A1/A1/c1 ),
    .Z(\V4/V4/s1 [1]));
 OR2_X1 \V4/V4/A1/A1/M2/_0_  (.A1(\V4/V4/A1/A1/M2/c1 ),
    .A2(\V4/V4/A1/A1/M2/c2 ),
    .ZN(\V4/V4/A1/A1/c2 ));
 AND2_X1 \V4/V4/A1/A1/M3/M1/_0_  (.A1(\V4/V4/v2 [2]),
    .A2(\V4/V4/v3 [2]),
    .ZN(\V4/V4/A1/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M3/M1/_1_  (.A(\V4/V4/v2 [2]),
    .B(\V4/V4/v3 [2]),
    .Z(\V4/V4/A1/A1/M3/s1 ));
 AND2_X1 \V4/V4/A1/A1/M3/M2/_0_  (.A1(\V4/V4/A1/A1/M3/s1 ),
    .A2(\V4/V4/A1/A1/c2 ),
    .ZN(\V4/V4/A1/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M3/M2/_1_  (.A(\V4/V4/A1/A1/M3/s1 ),
    .B(\V4/V4/A1/A1/c2 ),
    .Z(\V4/V4/s1 [2]));
 OR2_X1 \V4/V4/A1/A1/M3/_0_  (.A1(\V4/V4/A1/A1/M3/c1 ),
    .A2(\V4/V4/A1/A1/M3/c2 ),
    .ZN(\V4/V4/A1/A1/c3 ));
 AND2_X1 \V4/V4/A1/A1/M4/M1/_0_  (.A1(\V4/V4/v2 [3]),
    .A2(\V4/V4/v3 [3]),
    .ZN(\V4/V4/A1/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A1/A1/M4/M1/_1_  (.A(\V4/V4/v2 [3]),
    .B(\V4/V4/v3 [3]),
    .Z(\V4/V4/A1/A1/M4/s1 ));
 AND2_X1 \V4/V4/A1/A1/M4/M2/_0_  (.A1(\V4/V4/A1/A1/M4/s1 ),
    .A2(\V4/V4/A1/A1/c3 ),
    .ZN(\V4/V4/A1/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A1/A1/M4/M2/_1_  (.A(\V4/V4/A1/A1/M4/s1 ),
    .B(\V4/V4/A1/A1/c3 ),
    .Z(\V4/V4/s1 [3]));
 OR2_X1 \V4/V4/A1/A1/M4/_0_  (.A1(\V4/V4/A1/A1/M4/c1 ),
    .A2(\V4/V4/A1/A1/M4/c2 ),
    .ZN(\V4/V4/A1/c1 ));
 AND2_X1 \V4/V4/A1/A2/M1/M1/_0_  (.A1(\V4/V4/v2 [4]),
    .A2(\V4/V4/v3 [4]),
    .ZN(\V4/V4/A1/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M1/M1/_1_  (.A(\V4/V4/v2 [4]),
    .B(\V4/V4/v3 [4]),
    .Z(\V4/V4/A1/A2/M1/s1 ));
 AND2_X1 \V4/V4/A1/A2/M1/M2/_0_  (.A1(\V4/V4/A1/A2/M1/s1 ),
    .A2(\V4/V4/A1/c1 ),
    .ZN(\V4/V4/A1/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M1/M2/_1_  (.A(\V4/V4/A1/A2/M1/s1 ),
    .B(\V4/V4/A1/c1 ),
    .Z(\V4/V4/s1 [4]));
 OR2_X1 \V4/V4/A1/A2/M1/_0_  (.A1(\V4/V4/A1/A2/M1/c1 ),
    .A2(\V4/V4/A1/A2/M1/c2 ),
    .ZN(\V4/V4/A1/A2/c1 ));
 AND2_X1 \V4/V4/A1/A2/M2/M1/_0_  (.A1(\V4/V4/v2 [5]),
    .A2(\V4/V4/v3 [5]),
    .ZN(\V4/V4/A1/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M2/M1/_1_  (.A(\V4/V4/v2 [5]),
    .B(\V4/V4/v3 [5]),
    .Z(\V4/V4/A1/A2/M2/s1 ));
 AND2_X1 \V4/V4/A1/A2/M2/M2/_0_  (.A1(\V4/V4/A1/A2/M2/s1 ),
    .A2(\V4/V4/A1/A2/c1 ),
    .ZN(\V4/V4/A1/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M2/M2/_1_  (.A(\V4/V4/A1/A2/M2/s1 ),
    .B(\V4/V4/A1/A2/c1 ),
    .Z(\V4/V4/s1 [5]));
 OR2_X1 \V4/V4/A1/A2/M2/_0_  (.A1(\V4/V4/A1/A2/M2/c1 ),
    .A2(\V4/V4/A1/A2/M2/c2 ),
    .ZN(\V4/V4/A1/A2/c2 ));
 AND2_X1 \V4/V4/A1/A2/M3/M1/_0_  (.A1(\V4/V4/v2 [6]),
    .A2(\V4/V4/v3 [6]),
    .ZN(\V4/V4/A1/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M3/M1/_1_  (.A(\V4/V4/v2 [6]),
    .B(\V4/V4/v3 [6]),
    .Z(\V4/V4/A1/A2/M3/s1 ));
 AND2_X1 \V4/V4/A1/A2/M3/M2/_0_  (.A1(\V4/V4/A1/A2/M3/s1 ),
    .A2(\V4/V4/A1/A2/c2 ),
    .ZN(\V4/V4/A1/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M3/M2/_1_  (.A(\V4/V4/A1/A2/M3/s1 ),
    .B(\V4/V4/A1/A2/c2 ),
    .Z(\V4/V4/s1 [6]));
 OR2_X1 \V4/V4/A1/A2/M3/_0_  (.A1(\V4/V4/A1/A2/M3/c1 ),
    .A2(\V4/V4/A1/A2/M3/c2 ),
    .ZN(\V4/V4/A1/A2/c3 ));
 AND2_X1 \V4/V4/A1/A2/M4/M1/_0_  (.A1(\V4/V4/v2 [7]),
    .A2(\V4/V4/v3 [7]),
    .ZN(\V4/V4/A1/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A1/A2/M4/M1/_1_  (.A(\V4/V4/v2 [7]),
    .B(\V4/V4/v3 [7]),
    .Z(\V4/V4/A1/A2/M4/s1 ));
 AND2_X1 \V4/V4/A1/A2/M4/M2/_0_  (.A1(\V4/V4/A1/A2/M4/s1 ),
    .A2(\V4/V4/A1/A2/c3 ),
    .ZN(\V4/V4/A1/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A1/A2/M4/M2/_1_  (.A(\V4/V4/A1/A2/M4/s1 ),
    .B(\V4/V4/A1/A2/c3 ),
    .Z(\V4/V4/s1 [7]));
 OR2_X1 \V4/V4/A1/A2/M4/_0_  (.A1(\V4/V4/A1/A2/M4/c1 ),
    .A2(\V4/V4/A1/A2/M4/c2 ),
    .ZN(\V4/V4/c1 ));
 AND2_X1 \V4/V4/A2/A1/M1/M1/_0_  (.A1(\V4/V4/s1 [0]),
    .A2(\V4/V4/v1 [4]),
    .ZN(\V4/V4/A2/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M1/M1/_1_  (.A(\V4/V4/s1 [0]),
    .B(\V4/V4/v1 [4]),
    .Z(\V4/V4/A2/A1/M1/s1 ));
 AND2_X1 \V4/V4/A2/A1/M1/M2/_0_  (.A1(\V4/V4/A2/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V4/A2/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M1/M2/_1_  (.A(\V4/V4/A2/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/v4 [4]));
 OR2_X1 \V4/V4/A2/A1/M1/_0_  (.A1(\V4/V4/A2/A1/M1/c1 ),
    .A2(\V4/V4/A2/A1/M1/c2 ),
    .ZN(\V4/V4/A2/A1/c1 ));
 AND2_X1 \V4/V4/A2/A1/M2/M1/_0_  (.A1(\V4/V4/s1 [1]),
    .A2(\V4/V4/v1 [5]),
    .ZN(\V4/V4/A2/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M2/M1/_1_  (.A(\V4/V4/s1 [1]),
    .B(\V4/V4/v1 [5]),
    .Z(\V4/V4/A2/A1/M2/s1 ));
 AND2_X1 \V4/V4/A2/A1/M2/M2/_0_  (.A1(\V4/V4/A2/A1/M2/s1 ),
    .A2(\V4/V4/A2/A1/c1 ),
    .ZN(\V4/V4/A2/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M2/M2/_1_  (.A(\V4/V4/A2/A1/M2/s1 ),
    .B(\V4/V4/A2/A1/c1 ),
    .Z(\V4/v4 [5]));
 OR2_X1 \V4/V4/A2/A1/M2/_0_  (.A1(\V4/V4/A2/A1/M2/c1 ),
    .A2(\V4/V4/A2/A1/M2/c2 ),
    .ZN(\V4/V4/A2/A1/c2 ));
 AND2_X1 \V4/V4/A2/A1/M3/M1/_0_  (.A1(\V4/V4/s1 [2]),
    .A2(\V4/V4/v1 [6]),
    .ZN(\V4/V4/A2/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M3/M1/_1_  (.A(\V4/V4/s1 [2]),
    .B(\V4/V4/v1 [6]),
    .Z(\V4/V4/A2/A1/M3/s1 ));
 AND2_X1 \V4/V4/A2/A1/M3/M2/_0_  (.A1(\V4/V4/A2/A1/M3/s1 ),
    .A2(\V4/V4/A2/A1/c2 ),
    .ZN(\V4/V4/A2/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M3/M2/_1_  (.A(\V4/V4/A2/A1/M3/s1 ),
    .B(\V4/V4/A2/A1/c2 ),
    .Z(\V4/v4 [6]));
 OR2_X1 \V4/V4/A2/A1/M3/_0_  (.A1(\V4/V4/A2/A1/M3/c1 ),
    .A2(\V4/V4/A2/A1/M3/c2 ),
    .ZN(\V4/V4/A2/A1/c3 ));
 AND2_X1 \V4/V4/A2/A1/M4/M1/_0_  (.A1(\V4/V4/s1 [3]),
    .A2(\V4/V4/v1 [7]),
    .ZN(\V4/V4/A2/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A2/A1/M4/M1/_1_  (.A(\V4/V4/s1 [3]),
    .B(\V4/V4/v1 [7]),
    .Z(\V4/V4/A2/A1/M4/s1 ));
 AND2_X1 \V4/V4/A2/A1/M4/M2/_0_  (.A1(\V4/V4/A2/A1/M4/s1 ),
    .A2(\V4/V4/A2/A1/c3 ),
    .ZN(\V4/V4/A2/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A2/A1/M4/M2/_1_  (.A(\V4/V4/A2/A1/M4/s1 ),
    .B(\V4/V4/A2/A1/c3 ),
    .Z(\V4/v4 [7]));
 OR2_X1 \V4/V4/A2/A1/M4/_0_  (.A1(\V4/V4/A2/A1/M4/c1 ),
    .A2(\V4/V4/A2/A1/M4/c2 ),
    .ZN(\V4/V4/A2/c1 ));
 AND2_X1 \V4/V4/A2/A2/M1/M1/_0_  (.A1(\V4/V4/s1 [4]),
    .A2(net9),
    .ZN(\V4/V4/A2/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M1/M1/_1_  (.A(\V4/V4/s1 [4]),
    .B(net9),
    .Z(\V4/V4/A2/A2/M1/s1 ));
 AND2_X1 \V4/V4/A2/A2/M1/M2/_0_  (.A1(\V4/V4/A2/A2/M1/s1 ),
    .A2(\V4/V4/A2/c1 ),
    .ZN(\V4/V4/A2/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M1/M2/_1_  (.A(\V4/V4/A2/A2/M1/s1 ),
    .B(\V4/V4/A2/c1 ),
    .Z(\V4/V4/s2 [4]));
 OR2_X1 \V4/V4/A2/A2/M1/_0_  (.A1(\V4/V4/A2/A2/M1/c1 ),
    .A2(\V4/V4/A2/A2/M1/c2 ),
    .ZN(\V4/V4/A2/A2/c1 ));
 AND2_X1 \V4/V4/A2/A2/M2/M1/_0_  (.A1(\V4/V4/s1 [5]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M2/M1/_1_  (.A(\V4/V4/s1 [5]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M2/s1 ));
 AND2_X1 \V4/V4/A2/A2/M2/M2/_0_  (.A1(\V4/V4/A2/A2/M2/s1 ),
    .A2(\V4/V4/A2/A2/c1 ),
    .ZN(\V4/V4/A2/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M2/M2/_1_  (.A(\V4/V4/A2/A2/M2/s1 ),
    .B(\V4/V4/A2/A2/c1 ),
    .Z(\V4/V4/s2 [5]));
 OR2_X1 \V4/V4/A2/A2/M2/_0_  (.A1(\V4/V4/A2/A2/M2/c1 ),
    .A2(\V4/V4/A2/A2/M2/c2 ),
    .ZN(\V4/V4/A2/A2/c2 ));
 AND2_X1 \V4/V4/A2/A2/M3/M1/_0_  (.A1(\V4/V4/s1 [6]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M3/M1/_1_  (.A(\V4/V4/s1 [6]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M3/s1 ));
 AND2_X1 \V4/V4/A2/A2/M3/M2/_0_  (.A1(\V4/V4/A2/A2/M3/s1 ),
    .A2(\V4/V4/A2/A2/c2 ),
    .ZN(\V4/V4/A2/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M3/M2/_1_  (.A(\V4/V4/A2/A2/M3/s1 ),
    .B(\V4/V4/A2/A2/c2 ),
    .Z(\V4/V4/s2 [6]));
 OR2_X1 \V4/V4/A2/A2/M3/_0_  (.A1(\V4/V4/A2/A2/M3/c1 ),
    .A2(\V4/V4/A2/A2/M3/c2 ),
    .ZN(\V4/V4/A2/A2/c3 ));
 AND2_X1 \V4/V4/A2/A2/M4/M1/_0_  (.A1(\V4/V4/s1 [7]),
    .A2(ground),
    .ZN(\V4/V4/A2/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A2/A2/M4/M1/_1_  (.A(\V4/V4/s1 [7]),
    .B(ground),
    .Z(\V4/V4/A2/A2/M4/s1 ));
 AND2_X1 \V4/V4/A2/A2/M4/M2/_0_  (.A1(\V4/V4/A2/A2/M4/s1 ),
    .A2(\V4/V4/A2/A2/c3 ),
    .ZN(\V4/V4/A2/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A2/A2/M4/M2/_1_  (.A(\V4/V4/A2/A2/M4/s1 ),
    .B(\V4/V4/A2/A2/c3 ),
    .Z(\V4/V4/s2 [7]));
 OR2_X1 \V4/V4/A2/A2/M4/_0_  (.A1(\V4/V4/A2/A2/M4/c1 ),
    .A2(\V4/V4/A2/A2/M4/c2 ),
    .ZN(\V4/V4/c2 ));
 AND2_X1 \V4/V4/A3/A1/M1/M1/_0_  (.A1(\V4/V4/v4 [0]),
    .A2(\V4/V4/s2 [4]),
    .ZN(\V4/V4/A3/A1/M1/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M1/M1/_1_  (.A(\V4/V4/v4 [0]),
    .B(\V4/V4/s2 [4]),
    .Z(\V4/V4/A3/A1/M1/s1 ));
 AND2_X1 \V4/V4/A3/A1/M1/M2/_0_  (.A1(\V4/V4/A3/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/A3/A1/M1/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M1/M2/_1_  (.A(\V4/V4/A3/A1/M1/s1 ),
    .B(net10),
    .Z(\V4/v4 [8]));
 OR2_X1 \V4/V4/A3/A1/M1/_0_  (.A1(\V4/V4/A3/A1/M1/c1 ),
    .A2(\V4/V4/A3/A1/M1/c2 ),
    .ZN(\V4/V4/A3/A1/c1 ));
 AND2_X1 \V4/V4/A3/A1/M2/M1/_0_  (.A1(\V4/V4/v4 [1]),
    .A2(\V4/V4/s2 [5]),
    .ZN(\V4/V4/A3/A1/M2/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M2/M1/_1_  (.A(\V4/V4/v4 [1]),
    .B(\V4/V4/s2 [5]),
    .Z(\V4/V4/A3/A1/M2/s1 ));
 AND2_X1 \V4/V4/A3/A1/M2/M2/_0_  (.A1(\V4/V4/A3/A1/M2/s1 ),
    .A2(\V4/V4/A3/A1/c1 ),
    .ZN(\V4/V4/A3/A1/M2/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M2/M2/_1_  (.A(\V4/V4/A3/A1/M2/s1 ),
    .B(\V4/V4/A3/A1/c1 ),
    .Z(\V4/v4 [9]));
 OR2_X1 \V4/V4/A3/A1/M2/_0_  (.A1(\V4/V4/A3/A1/M2/c1 ),
    .A2(\V4/V4/A3/A1/M2/c2 ),
    .ZN(\V4/V4/A3/A1/c2 ));
 AND2_X1 \V4/V4/A3/A1/M3/M1/_0_  (.A1(\V4/V4/v4 [2]),
    .A2(\V4/V4/s2 [6]),
    .ZN(\V4/V4/A3/A1/M3/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M3/M1/_1_  (.A(\V4/V4/v4 [2]),
    .B(\V4/V4/s2 [6]),
    .Z(\V4/V4/A3/A1/M3/s1 ));
 AND2_X1 \V4/V4/A3/A1/M3/M2/_0_  (.A1(\V4/V4/A3/A1/M3/s1 ),
    .A2(\V4/V4/A3/A1/c2 ),
    .ZN(\V4/V4/A3/A1/M3/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M3/M2/_1_  (.A(\V4/V4/A3/A1/M3/s1 ),
    .B(\V4/V4/A3/A1/c2 ),
    .Z(\V4/v4 [10]));
 OR2_X1 \V4/V4/A3/A1/M3/_0_  (.A1(\V4/V4/A3/A1/M3/c1 ),
    .A2(\V4/V4/A3/A1/M3/c2 ),
    .ZN(\V4/V4/A3/A1/c3 ));
 AND2_X1 \V4/V4/A3/A1/M4/M1/_0_  (.A1(\V4/V4/v4 [3]),
    .A2(\V4/V4/s2 [7]),
    .ZN(\V4/V4/A3/A1/M4/c1 ));
 XOR2_X2 \V4/V4/A3/A1/M4/M1/_1_  (.A(\V4/V4/v4 [3]),
    .B(\V4/V4/s2 [7]),
    .Z(\V4/V4/A3/A1/M4/s1 ));
 AND2_X1 \V4/V4/A3/A1/M4/M2/_0_  (.A1(\V4/V4/A3/A1/M4/s1 ),
    .A2(\V4/V4/A3/A1/c3 ),
    .ZN(\V4/V4/A3/A1/M4/c2 ));
 XOR2_X2 \V4/V4/A3/A1/M4/M2/_1_  (.A(\V4/V4/A3/A1/M4/s1 ),
    .B(\V4/V4/A3/A1/c3 ),
    .Z(\V4/v4 [11]));
 OR2_X1 \V4/V4/A3/A1/M4/_0_  (.A1(\V4/V4/A3/A1/M4/c1 ),
    .A2(\V4/V4/A3/A1/M4/c2 ),
    .ZN(\V4/V4/A3/c1 ));
 AND2_X1 \V4/V4/A3/A2/M1/M1/_0_  (.A1(\V4/V4/v4 [4]),
    .A2(\V4/V4/c3 ),
    .ZN(\V4/V4/A3/A2/M1/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M1/M1/_1_  (.A(\V4/V4/v4 [4]),
    .B(\V4/V4/c3 ),
    .Z(\V4/V4/A3/A2/M1/s1 ));
 AND2_X1 \V4/V4/A3/A2/M1/M2/_0_  (.A1(\V4/V4/A3/A2/M1/s1 ),
    .A2(\V4/V4/A3/c1 ),
    .ZN(\V4/V4/A3/A2/M1/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M1/M2/_1_  (.A(\V4/V4/A3/A2/M1/s1 ),
    .B(\V4/V4/A3/c1 ),
    .Z(\V4/v4 [12]));
 OR2_X1 \V4/V4/A3/A2/M1/_0_  (.A1(\V4/V4/A3/A2/M1/c1 ),
    .A2(\V4/V4/A3/A2/M1/c2 ),
    .ZN(\V4/V4/A3/A2/c1 ));
 AND2_X1 \V4/V4/A3/A2/M2/M1/_0_  (.A1(\V4/V4/v4 [5]),
    .A2(net10),
    .ZN(\V4/V4/A3/A2/M2/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M2/M1/_1_  (.A(\V4/V4/v4 [5]),
    .B(net10),
    .Z(\V4/V4/A3/A2/M2/s1 ));
 AND2_X1 \V4/V4/A3/A2/M2/M2/_0_  (.A1(\V4/V4/A3/A2/M2/s1 ),
    .A2(\V4/V4/A3/A2/c1 ),
    .ZN(\V4/V4/A3/A2/M2/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M2/M2/_1_  (.A(\V4/V4/A3/A2/M2/s1 ),
    .B(\V4/V4/A3/A2/c1 ),
    .Z(\V4/v4 [13]));
 OR2_X1 \V4/V4/A3/A2/M2/_0_  (.A1(\V4/V4/A3/A2/M2/c1 ),
    .A2(\V4/V4/A3/A2/M2/c2 ),
    .ZN(\V4/V4/A3/A2/c2 ));
 AND2_X1 \V4/V4/A3/A2/M3/M1/_0_  (.A1(\V4/V4/v4 [6]),
    .A2(ground),
    .ZN(\V4/V4/A3/A2/M3/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M3/M1/_1_  (.A(\V4/V4/v4 [6]),
    .B(ground),
    .Z(\V4/V4/A3/A2/M3/s1 ));
 AND2_X1 \V4/V4/A3/A2/M3/M2/_0_  (.A1(\V4/V4/A3/A2/M3/s1 ),
    .A2(\V4/V4/A3/A2/c2 ),
    .ZN(\V4/V4/A3/A2/M3/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M3/M2/_1_  (.A(\V4/V4/A3/A2/M3/s1 ),
    .B(\V4/V4/A3/A2/c2 ),
    .Z(\V4/v4 [14]));
 OR2_X1 \V4/V4/A3/A2/M3/_0_  (.A1(\V4/V4/A3/A2/M3/c1 ),
    .A2(\V4/V4/A3/A2/M3/c2 ),
    .ZN(\V4/V4/A3/A2/c3 ));
 AND2_X1 \V4/V4/A3/A2/M4/M1/_0_  (.A1(\V4/V4/v4 [7]),
    .A2(ground),
    .ZN(\V4/V4/A3/A2/M4/c1 ));
 XOR2_X2 \V4/V4/A3/A2/M4/M1/_1_  (.A(\V4/V4/v4 [7]),
    .B(ground),
    .Z(\V4/V4/A3/A2/M4/s1 ));
 AND2_X1 \V4/V4/A3/A2/M4/M2/_0_  (.A1(\V4/V4/A3/A2/M4/s1 ),
    .A2(\V4/V4/A3/A2/c3 ),
    .ZN(\V4/V4/A3/A2/M4/c2 ));
 XOR2_X2 \V4/V4/A3/A2/M4/M2/_1_  (.A(\V4/V4/A3/A2/M4/s1 ),
    .B(\V4/V4/A3/A2/c3 ),
    .Z(\V4/v4 [15]));
 OR2_X1 \V4/V4/A3/A2/M4/_0_  (.A1(\V4/V4/A3/A2/M4/c1 ),
    .A2(\V4/V4/A3/A2/M4/c2 ),
    .ZN(\V4/V4/overflow ));
 AND2_X1 \V4/V4/V1/A1/M1/M1/_0_  (.A1(\V4/V4/V1/v2 [0]),
    .A2(\V4/V4/V1/v3 [0]),
    .ZN(\V4/V4/V1/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M1/M1/_1_  (.A(\V4/V4/V1/v2 [0]),
    .B(\V4/V4/V1/v3 [0]),
    .Z(\V4/V4/V1/A1/M1/s1 ));
 AND2_X1 \V4/V4/V1/A1/M1/M2/_0_  (.A1(\V4/V4/V1/A1/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V4/V1/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M1/M2/_1_  (.A(\V4/V4/V1/A1/M1/s1 ),
    .B(net1),
    .Z(\V4/V4/V1/s1 [0]));
 OR2_X1 \V4/V4/V1/A1/M1/_0_  (.A1(\V4/V4/V1/A1/M1/c1 ),
    .A2(\V4/V4/V1/A1/M1/c2 ),
    .ZN(\V4/V4/V1/A1/c1 ));
 AND2_X1 \V4/V4/V1/A1/M2/M1/_0_  (.A1(\V4/V4/V1/v2 [1]),
    .A2(\V4/V4/V1/v3 [1]),
    .ZN(\V4/V4/V1/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M2/M1/_1_  (.A(\V4/V4/V1/v2 [1]),
    .B(\V4/V4/V1/v3 [1]),
    .Z(\V4/V4/V1/A1/M2/s1 ));
 AND2_X1 \V4/V4/V1/A1/M2/M2/_0_  (.A1(\V4/V4/V1/A1/M2/s1 ),
    .A2(\V4/V4/V1/A1/c1 ),
    .ZN(\V4/V4/V1/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M2/M2/_1_  (.A(\V4/V4/V1/A1/M2/s1 ),
    .B(\V4/V4/V1/A1/c1 ),
    .Z(\V4/V4/V1/s1 [1]));
 OR2_X1 \V4/V4/V1/A1/M2/_0_  (.A1(\V4/V4/V1/A1/M2/c1 ),
    .A2(\V4/V4/V1/A1/M2/c2 ),
    .ZN(\V4/V4/V1/A1/c2 ));
 AND2_X1 \V4/V4/V1/A1/M3/M1/_0_  (.A1(\V4/V4/V1/v2 [2]),
    .A2(\V4/V4/V1/v3 [2]),
    .ZN(\V4/V4/V1/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M3/M1/_1_  (.A(\V4/V4/V1/v2 [2]),
    .B(\V4/V4/V1/v3 [2]),
    .Z(\V4/V4/V1/A1/M3/s1 ));
 AND2_X1 \V4/V4/V1/A1/M3/M2/_0_  (.A1(\V4/V4/V1/A1/M3/s1 ),
    .A2(\V4/V4/V1/A1/c2 ),
    .ZN(\V4/V4/V1/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M3/M2/_1_  (.A(\V4/V4/V1/A1/M3/s1 ),
    .B(\V4/V4/V1/A1/c2 ),
    .Z(\V4/V4/V1/s1 [2]));
 OR2_X1 \V4/V4/V1/A1/M3/_0_  (.A1(\V4/V4/V1/A1/M3/c1 ),
    .A2(\V4/V4/V1/A1/M3/c2 ),
    .ZN(\V4/V4/V1/A1/c3 ));
 AND2_X1 \V4/V4/V1/A1/M4/M1/_0_  (.A1(\V4/V4/V1/v2 [3]),
    .A2(\V4/V4/V1/v3 [3]),
    .ZN(\V4/V4/V1/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A1/M4/M1/_1_  (.A(\V4/V4/V1/v2 [3]),
    .B(\V4/V4/V1/v3 [3]),
    .Z(\V4/V4/V1/A1/M4/s1 ));
 AND2_X1 \V4/V4/V1/A1/M4/M2/_0_  (.A1(\V4/V4/V1/A1/M4/s1 ),
    .A2(\V4/V4/V1/A1/c3 ),
    .ZN(\V4/V4/V1/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A1/M4/M2/_1_  (.A(\V4/V4/V1/A1/M4/s1 ),
    .B(\V4/V4/V1/A1/c3 ),
    .Z(\V4/V4/V1/s1 [3]));
 OR2_X1 \V4/V4/V1/A1/M4/_0_  (.A1(\V4/V4/V1/A1/M4/c1 ),
    .A2(\V4/V4/V1/A1/M4/c2 ),
    .ZN(\V4/V4/V1/c1 ));
 AND2_X1 \V4/V4/V1/A2/M1/M1/_0_  (.A1(\V4/V4/V1/s1 [0]),
    .A2(\V4/V4/V1/v1 [2]),
    .ZN(\V4/V4/V1/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M1/M1/_1_  (.A(\V4/V4/V1/s1 [0]),
    .B(\V4/V4/V1/v1 [2]),
    .Z(\V4/V4/V1/A2/M1/s1 ));
 AND2_X1 \V4/V4/V1/A2/M1/M2/_0_  (.A1(\V4/V4/V1/A2/M1/s1 ),
    .A2(net1),
    .ZN(\V4/V4/V1/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M1/M2/_1_  (.A(\V4/V4/V1/A2/M1/s1 ),
    .B(net1),
    .Z(\V4/v4 [2]));
 OR2_X1 \V4/V4/V1/A2/M1/_0_  (.A1(\V4/V4/V1/A2/M1/c1 ),
    .A2(\V4/V4/V1/A2/M1/c2 ),
    .ZN(\V4/V4/V1/A2/c1 ));
 AND2_X1 \V4/V4/V1/A2/M2/M1/_0_  (.A1(\V4/V4/V1/s1 [1]),
    .A2(\V4/V4/V1/v1 [3]),
    .ZN(\V4/V4/V1/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M2/M1/_1_  (.A(\V4/V4/V1/s1 [1]),
    .B(\V4/V4/V1/v1 [3]),
    .Z(\V4/V4/V1/A2/M2/s1 ));
 AND2_X1 \V4/V4/V1/A2/M2/M2/_0_  (.A1(\V4/V4/V1/A2/M2/s1 ),
    .A2(\V4/V4/V1/A2/c1 ),
    .ZN(\V4/V4/V1/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M2/M2/_1_  (.A(\V4/V4/V1/A2/M2/s1 ),
    .B(\V4/V4/V1/A2/c1 ),
    .Z(\V4/v4 [3]));
 OR2_X1 \V4/V4/V1/A2/M2/_0_  (.A1(\V4/V4/V1/A2/M2/c1 ),
    .A2(\V4/V4/V1/A2/M2/c2 ),
    .ZN(\V4/V4/V1/A2/c2 ));
 AND2_X1 \V4/V4/V1/A2/M3/M1/_0_  (.A1(\V4/V4/V1/s1 [2]),
    .A2(net1),
    .ZN(\V4/V4/V1/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M3/M1/_1_  (.A(\V4/V4/V1/s1 [2]),
    .B(net1),
    .Z(\V4/V4/V1/A2/M3/s1 ));
 AND2_X1 \V4/V4/V1/A2/M3/M2/_0_  (.A1(\V4/V4/V1/A2/M3/s1 ),
    .A2(\V4/V4/V1/A2/c2 ),
    .ZN(\V4/V4/V1/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M3/M2/_1_  (.A(\V4/V4/V1/A2/M3/s1 ),
    .B(\V4/V4/V1/A2/c2 ),
    .Z(\V4/V4/V1/s2 [2]));
 OR2_X1 \V4/V4/V1/A2/M3/_0_  (.A1(\V4/V4/V1/A2/M3/c1 ),
    .A2(\V4/V4/V1/A2/M3/c2 ),
    .ZN(\V4/V4/V1/A2/c3 ));
 AND2_X1 \V4/V4/V1/A2/M4/M1/_0_  (.A1(\V4/V4/V1/s1 [3]),
    .A2(net10),
    .ZN(\V4/V4/V1/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A2/M4/M1/_1_  (.A(\V4/V4/V1/s1 [3]),
    .B(net10),
    .Z(\V4/V4/V1/A2/M4/s1 ));
 AND2_X1 \V4/V4/V1/A2/M4/M2/_0_  (.A1(\V4/V4/V1/A2/M4/s1 ),
    .A2(\V4/V4/V1/A2/c3 ),
    .ZN(\V4/V4/V1/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A2/M4/M2/_1_  (.A(\V4/V4/V1/A2/M4/s1 ),
    .B(\V4/V4/V1/A2/c3 ),
    .Z(\V4/V4/V1/s2 [3]));
 OR2_X1 \V4/V4/V1/A2/M4/_0_  (.A1(\V4/V4/V1/A2/M4/c1 ),
    .A2(\V4/V4/V1/A2/M4/c2 ),
    .ZN(\V4/V4/V1/c2 ));
 AND2_X1 \V4/V4/V1/A3/M1/M1/_0_  (.A1(\V4/V4/V1/v4 [0]),
    .A2(\V4/V4/V1/s2 [2]),
    .ZN(\V4/V4/V1/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M1/M1/_1_  (.A(\V4/V4/V1/v4 [0]),
    .B(\V4/V4/V1/s2 [2]),
    .Z(\V4/V4/V1/A3/M1/s1 ));
 AND2_X1 \V4/V4/V1/A3/M1/M2/_0_  (.A1(\V4/V4/V1/A3/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V4/V1/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M1/M2/_1_  (.A(\V4/V4/V1/A3/M1/s1 ),
    .B(net1),
    .Z(\V4/V4/v1 [4]));
 OR2_X1 \V4/V4/V1/A3/M1/_0_  (.A1(\V4/V4/V1/A3/M1/c1 ),
    .A2(\V4/V4/V1/A3/M1/c2 ),
    .ZN(\V4/V4/V1/A3/c1 ));
 AND2_X1 \V4/V4/V1/A3/M2/M1/_0_  (.A1(\V4/V4/V1/v4 [1]),
    .A2(\V4/V4/V1/s2 [3]),
    .ZN(\V4/V4/V1/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M2/M1/_1_  (.A(\V4/V4/V1/v4 [1]),
    .B(\V4/V4/V1/s2 [3]),
    .Z(\V4/V4/V1/A3/M2/s1 ));
 AND2_X1 \V4/V4/V1/A3/M2/M2/_0_  (.A1(\V4/V4/V1/A3/M2/s1 ),
    .A2(\V4/V4/V1/A3/c1 ),
    .ZN(\V4/V4/V1/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M2/M2/_1_  (.A(\V4/V4/V1/A3/M2/s1 ),
    .B(\V4/V4/V1/A3/c1 ),
    .Z(\V4/V4/v1 [5]));
 OR2_X1 \V4/V4/V1/A3/M2/_0_  (.A1(\V4/V4/V1/A3/M2/c1 ),
    .A2(\V4/V4/V1/A3/M2/c2 ),
    .ZN(\V4/V4/V1/A3/c2 ));
 AND2_X1 \V4/V4/V1/A3/M3/M1/_0_  (.A1(\V4/V4/V1/v4 [2]),
    .A2(\V4/V4/V1/c3 ),
    .ZN(\V4/V4/V1/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M3/M1/_1_  (.A(\V4/V4/V1/v4 [2]),
    .B(\V4/V4/V1/c3 ),
    .Z(\V4/V4/V1/A3/M3/s1 ));
 AND2_X1 \V4/V4/V1/A3/M3/M2/_0_  (.A1(\V4/V4/V1/A3/M3/s1 ),
    .A2(\V4/V4/V1/A3/c2 ),
    .ZN(\V4/V4/V1/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M3/M2/_1_  (.A(\V4/V4/V1/A3/M3/s1 ),
    .B(\V4/V4/V1/A3/c2 ),
    .Z(\V4/V4/v1 [6]));
 OR2_X1 \V4/V4/V1/A3/M3/_0_  (.A1(\V4/V4/V1/A3/M3/c1 ),
    .A2(\V4/V4/V1/A3/M3/c2 ),
    .ZN(\V4/V4/V1/A3/c3 ));
 AND2_X1 \V4/V4/V1/A3/M4/M1/_0_  (.A1(\V4/V4/V1/v4 [3]),
    .A2(net9),
    .ZN(\V4/V4/V1/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V1/A3/M4/M1/_1_  (.A(\V4/V4/V1/v4 [3]),
    .B(net9),
    .Z(\V4/V4/V1/A3/M4/s1 ));
 AND2_X1 \V4/V4/V1/A3/M4/M2/_0_  (.A1(\V4/V4/V1/A3/M4/s1 ),
    .A2(\V4/V4/V1/A3/c3 ),
    .ZN(\V4/V4/V1/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V1/A3/M4/M2/_1_  (.A(\V4/V4/V1/A3/M4/s1 ),
    .B(\V4/V4/V1/A3/c3 ),
    .Z(\V4/V4/v1 [7]));
 OR2_X1 \V4/V4/V1/A3/M4/_0_  (.A1(\V4/V4/V1/A3/M4/c1 ),
    .A2(\V4/V4/V1/A3/M4/c2 ),
    .ZN(\V4/V4/V1/overflow ));
 AND2_X1 \V4/V4/V1/V1/HA1/_0_  (.A1(\V4/V4/V1/V1/w2 ),
    .A2(\V4/V4/V1/V1/w1 ),
    .ZN(\V4/V4/V1/V1/w4 ));
 XOR2_X2 \V4/V4/V1/V1/HA1/_1_  (.A(\V4/V4/V1/V1/w2 ),
    .B(\V4/V4/V1/V1/w1 ),
    .Z(\V4/v4 [1]));
 AND2_X1 \V4/V4/V1/V1/HA2/_0_  (.A1(\V4/V4/V1/V1/w4 ),
    .A2(\V4/V4/V1/V1/w3 ),
    .ZN(\V4/V4/V1/v1 [3]));
 XOR2_X2 \V4/V4/V1/V1/HA2/_1_  (.A(\V4/V4/V1/V1/w4 ),
    .B(\V4/V4/V1/V1/w3 ),
    .Z(\V4/V4/V1/v1 [2]));
 AND2_X1 \V4/V4/V1/V1/_0_  (.A1(net33),
    .A2(net14),
    .ZN(\V4/v4 [0]));
 AND2_X1 \V4/V4/V1/V1/_1_  (.A1(net33),
    .A2(B[25]),
    .ZN(\V4/V4/V1/V1/w1 ));
 AND2_X1 \V4/V4/V1/V1/_2_  (.A1(net14),
    .A2(net32),
    .ZN(\V4/V4/V1/V1/w2 ));
 AND2_X1 \V4/V4/V1/V1/_3_  (.A1(B[25]),
    .A2(net32),
    .ZN(\V4/V4/V1/V1/w3 ));
 AND2_X1 \V4/V4/V1/V2/HA1/_0_  (.A1(\V4/V4/V1/V2/w2 ),
    .A2(\V4/V4/V1/V2/w1 ),
    .ZN(\V4/V4/V1/V2/w4 ));
 XOR2_X2 \V4/V4/V1/V2/HA1/_1_  (.A(\V4/V4/V1/V2/w2 ),
    .B(\V4/V4/V1/V2/w1 ),
    .Z(\V4/V4/V1/v2 [1]));
 AND2_X1 \V4/V4/V1/V2/HA2/_0_  (.A1(\V4/V4/V1/V2/w4 ),
    .A2(\V4/V4/V1/V2/w3 ),
    .ZN(\V4/V4/V1/v2 [3]));
 XOR2_X2 \V4/V4/V1/V2/HA2/_1_  (.A(\V4/V4/V1/V2/w4 ),
    .B(\V4/V4/V1/V2/w3 ),
    .Z(\V4/V4/V1/v2 [2]));
 AND2_X1 \V4/V4/V1/V2/_0_  (.A1(net31),
    .A2(net14),
    .ZN(\V4/V4/V1/v2 [0]));
 AND2_X1 \V4/V4/V1/V2/_1_  (.A1(net31),
    .A2(B[25]),
    .ZN(\V4/V4/V1/V2/w1 ));
 AND2_X1 \V4/V4/V1/V2/_2_  (.A1(net14),
    .A2(net30),
    .ZN(\V4/V4/V1/V2/w2 ));
 AND2_X1 \V4/V4/V1/V2/_3_  (.A1(B[25]),
    .A2(net30),
    .ZN(\V4/V4/V1/V2/w3 ));
 AND2_X1 \V4/V4/V1/V3/HA1/_0_  (.A1(\V4/V4/V1/V3/w2 ),
    .A2(\V4/V4/V1/V3/w1 ),
    .ZN(\V4/V4/V1/V3/w4 ));
 XOR2_X2 \V4/V4/V1/V3/HA1/_1_  (.A(\V4/V4/V1/V3/w2 ),
    .B(\V4/V4/V1/V3/w1 ),
    .Z(\V4/V4/V1/v3 [1]));
 AND2_X1 \V4/V4/V1/V3/HA2/_0_  (.A1(\V4/V4/V1/V3/w4 ),
    .A2(\V4/V4/V1/V3/w3 ),
    .ZN(\V4/V4/V1/v3 [3]));
 XOR2_X2 \V4/V4/V1/V3/HA2/_1_  (.A(\V4/V4/V1/V3/w4 ),
    .B(\V4/V4/V1/V3/w3 ),
    .Z(\V4/V4/V1/v3 [2]));
 AND2_X1 \V4/V4/V1/V3/_0_  (.A1(net33),
    .A2(net13),
    .ZN(\V4/V4/V1/v3 [0]));
 AND2_X1 \V4/V4/V1/V3/_1_  (.A1(net33),
    .A2(B[27]),
    .ZN(\V4/V4/V1/V3/w1 ));
 AND2_X1 \V4/V4/V1/V3/_2_  (.A1(net13),
    .A2(net32),
    .ZN(\V4/V4/V1/V3/w2 ));
 AND2_X1 \V4/V4/V1/V3/_3_  (.A1(B[27]),
    .A2(net32),
    .ZN(\V4/V4/V1/V3/w3 ));
 AND2_X1 \V4/V4/V1/V4/HA1/_0_  (.A1(\V4/V4/V1/V4/w2 ),
    .A2(\V4/V4/V1/V4/w1 ),
    .ZN(\V4/V4/V1/V4/w4 ));
 XOR2_X2 \V4/V4/V1/V4/HA1/_1_  (.A(\V4/V4/V1/V4/w2 ),
    .B(\V4/V4/V1/V4/w1 ),
    .Z(\V4/V4/V1/v4 [1]));
 AND2_X1 \V4/V4/V1/V4/HA2/_0_  (.A1(\V4/V4/V1/V4/w4 ),
    .A2(\V4/V4/V1/V4/w3 ),
    .ZN(\V4/V4/V1/v4 [3]));
 XOR2_X2 \V4/V4/V1/V4/HA2/_1_  (.A(\V4/V4/V1/V4/w4 ),
    .B(\V4/V4/V1/V4/w3 ),
    .Z(\V4/V4/V1/v4 [2]));
 AND2_X1 \V4/V4/V1/V4/_0_  (.A1(net31),
    .A2(net13),
    .ZN(\V4/V4/V1/v4 [0]));
 AND2_X1 \V4/V4/V1/V4/_1_  (.A1(net31),
    .A2(B[27]),
    .ZN(\V4/V4/V1/V4/w1 ));
 AND2_X1 \V4/V4/V1/V4/_2_  (.A1(net13),
    .A2(net30),
    .ZN(\V4/V4/V1/V4/w2 ));
 AND2_X1 \V4/V4/V1/V4/_3_  (.A1(B[27]),
    .A2(net30),
    .ZN(\V4/V4/V1/V4/w3 ));
 OR2_X1 \V4/V4/V1/_0_  (.A1(\V4/V4/V1/c1 ),
    .A2(\V4/V4/V1/c2 ),
    .ZN(\V4/V4/V1/c3 ));
 AND2_X1 \V4/V4/V2/A1/M1/M1/_0_  (.A1(\V4/V4/V2/v2 [0]),
    .A2(\V4/V4/V2/v3 [0]),
    .ZN(\V4/V4/V2/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M1/M1/_1_  (.A(\V4/V4/V2/v2 [0]),
    .B(\V4/V4/V2/v3 [0]),
    .Z(\V4/V4/V2/A1/M1/s1 ));
 AND2_X1 \V4/V4/V2/A1/M1/M2/_0_  (.A1(\V4/V4/V2/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/V2/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M1/M2/_1_  (.A(\V4/V4/V2/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/V2/s1 [0]));
 OR2_X1 \V4/V4/V2/A1/M1/_0_  (.A1(\V4/V4/V2/A1/M1/c1 ),
    .A2(\V4/V4/V2/A1/M1/c2 ),
    .ZN(\V4/V4/V2/A1/c1 ));
 AND2_X1 \V4/V4/V2/A1/M2/M1/_0_  (.A1(\V4/V4/V2/v2 [1]),
    .A2(\V4/V4/V2/v3 [1]),
    .ZN(\V4/V4/V2/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M2/M1/_1_  (.A(\V4/V4/V2/v2 [1]),
    .B(\V4/V4/V2/v3 [1]),
    .Z(\V4/V4/V2/A1/M2/s1 ));
 AND2_X1 \V4/V4/V2/A1/M2/M2/_0_  (.A1(\V4/V4/V2/A1/M2/s1 ),
    .A2(\V4/V4/V2/A1/c1 ),
    .ZN(\V4/V4/V2/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M2/M2/_1_  (.A(\V4/V4/V2/A1/M2/s1 ),
    .B(\V4/V4/V2/A1/c1 ),
    .Z(\V4/V4/V2/s1 [1]));
 OR2_X1 \V4/V4/V2/A1/M2/_0_  (.A1(\V4/V4/V2/A1/M2/c1 ),
    .A2(\V4/V4/V2/A1/M2/c2 ),
    .ZN(\V4/V4/V2/A1/c2 ));
 AND2_X1 \V4/V4/V2/A1/M3/M1/_0_  (.A1(\V4/V4/V2/v2 [2]),
    .A2(\V4/V4/V2/v3 [2]),
    .ZN(\V4/V4/V2/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M3/M1/_1_  (.A(\V4/V4/V2/v2 [2]),
    .B(\V4/V4/V2/v3 [2]),
    .Z(\V4/V4/V2/A1/M3/s1 ));
 AND2_X1 \V4/V4/V2/A1/M3/M2/_0_  (.A1(\V4/V4/V2/A1/M3/s1 ),
    .A2(\V4/V4/V2/A1/c2 ),
    .ZN(\V4/V4/V2/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M3/M2/_1_  (.A(\V4/V4/V2/A1/M3/s1 ),
    .B(\V4/V4/V2/A1/c2 ),
    .Z(\V4/V4/V2/s1 [2]));
 OR2_X1 \V4/V4/V2/A1/M3/_0_  (.A1(\V4/V4/V2/A1/M3/c1 ),
    .A2(\V4/V4/V2/A1/M3/c2 ),
    .ZN(\V4/V4/V2/A1/c3 ));
 AND2_X1 \V4/V4/V2/A1/M4/M1/_0_  (.A1(\V4/V4/V2/v2 [3]),
    .A2(\V4/V4/V2/v3 [3]),
    .ZN(\V4/V4/V2/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A1/M4/M1/_1_  (.A(\V4/V4/V2/v2 [3]),
    .B(\V4/V4/V2/v3 [3]),
    .Z(\V4/V4/V2/A1/M4/s1 ));
 AND2_X1 \V4/V4/V2/A1/M4/M2/_0_  (.A1(\V4/V4/V2/A1/M4/s1 ),
    .A2(\V4/V4/V2/A1/c3 ),
    .ZN(\V4/V4/V2/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A1/M4/M2/_1_  (.A(\V4/V4/V2/A1/M4/s1 ),
    .B(\V4/V4/V2/A1/c3 ),
    .Z(\V4/V4/V2/s1 [3]));
 OR2_X1 \V4/V4/V2/A1/M4/_0_  (.A1(\V4/V4/V2/A1/M4/c1 ),
    .A2(\V4/V4/V2/A1/M4/c2 ),
    .ZN(\V4/V4/V2/c1 ));
 AND2_X1 \V4/V4/V2/A2/M1/M1/_0_  (.A1(\V4/V4/V2/s1 [0]),
    .A2(\V4/V4/V2/v1 [2]),
    .ZN(\V4/V4/V2/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M1/M1/_1_  (.A(\V4/V4/V2/s1 [0]),
    .B(\V4/V4/V2/v1 [2]),
    .Z(\V4/V4/V2/A2/M1/s1 ));
 AND2_X1 \V4/V4/V2/A2/M1/M2/_0_  (.A1(\V4/V4/V2/A2/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/V2/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M1/M2/_1_  (.A(\V4/V4/V2/A2/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/v2 [2]));
 OR2_X1 \V4/V4/V2/A2/M1/_0_  (.A1(\V4/V4/V2/A2/M1/c1 ),
    .A2(\V4/V4/V2/A2/M1/c2 ),
    .ZN(\V4/V4/V2/A2/c1 ));
 AND2_X1 \V4/V4/V2/A2/M2/M1/_0_  (.A1(\V4/V4/V2/s1 [1]),
    .A2(\V4/V4/V2/v1 [3]),
    .ZN(\V4/V4/V2/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M2/M1/_1_  (.A(\V4/V4/V2/s1 [1]),
    .B(\V4/V4/V2/v1 [3]),
    .Z(\V4/V4/V2/A2/M2/s1 ));
 AND2_X1 \V4/V4/V2/A2/M2/M2/_0_  (.A1(\V4/V4/V2/A2/M2/s1 ),
    .A2(\V4/V4/V2/A2/c1 ),
    .ZN(\V4/V4/V2/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M2/M2/_1_  (.A(\V4/V4/V2/A2/M2/s1 ),
    .B(\V4/V4/V2/A2/c1 ),
    .Z(\V4/V4/v2 [3]));
 OR2_X1 \V4/V4/V2/A2/M2/_0_  (.A1(\V4/V4/V2/A2/M2/c1 ),
    .A2(\V4/V4/V2/A2/M2/c2 ),
    .ZN(\V4/V4/V2/A2/c2 ));
 AND2_X1 \V4/V4/V2/A2/M3/M1/_0_  (.A1(\V4/V4/V2/s1 [2]),
    .A2(net9),
    .ZN(\V4/V4/V2/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M3/M1/_1_  (.A(\V4/V4/V2/s1 [2]),
    .B(net9),
    .Z(\V4/V4/V2/A2/M3/s1 ));
 AND2_X1 \V4/V4/V2/A2/M3/M2/_0_  (.A1(\V4/V4/V2/A2/M3/s1 ),
    .A2(\V4/V4/V2/A2/c2 ),
    .ZN(\V4/V4/V2/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M3/M2/_1_  (.A(\V4/V4/V2/A2/M3/s1 ),
    .B(\V4/V4/V2/A2/c2 ),
    .Z(\V4/V4/V2/s2 [2]));
 OR2_X1 \V4/V4/V2/A2/M3/_0_  (.A1(\V4/V4/V2/A2/M3/c1 ),
    .A2(\V4/V4/V2/A2/M3/c2 ),
    .ZN(\V4/V4/V2/A2/c3 ));
 AND2_X1 \V4/V4/V2/A2/M4/M1/_0_  (.A1(\V4/V4/V2/s1 [3]),
    .A2(net9),
    .ZN(\V4/V4/V2/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A2/M4/M1/_1_  (.A(\V4/V4/V2/s1 [3]),
    .B(net9),
    .Z(\V4/V4/V2/A2/M4/s1 ));
 AND2_X1 \V4/V4/V2/A2/M4/M2/_0_  (.A1(\V4/V4/V2/A2/M4/s1 ),
    .A2(\V4/V4/V2/A2/c3 ),
    .ZN(\V4/V4/V2/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A2/M4/M2/_1_  (.A(\V4/V4/V2/A2/M4/s1 ),
    .B(\V4/V4/V2/A2/c3 ),
    .Z(\V4/V4/V2/s2 [3]));
 OR2_X1 \V4/V4/V2/A2/M4/_0_  (.A1(\V4/V4/V2/A2/M4/c1 ),
    .A2(\V4/V4/V2/A2/M4/c2 ),
    .ZN(\V4/V4/V2/c2 ));
 AND2_X1 \V4/V4/V2/A3/M1/M1/_0_  (.A1(\V4/V4/V2/v4 [0]),
    .A2(\V4/V4/V2/s2 [2]),
    .ZN(\V4/V4/V2/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M1/M1/_1_  (.A(\V4/V4/V2/v4 [0]),
    .B(\V4/V4/V2/s2 [2]),
    .Z(\V4/V4/V2/A3/M1/s1 ));
 AND2_X1 \V4/V4/V2/A3/M1/M2/_0_  (.A1(\V4/V4/V2/A3/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/V2/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M1/M2/_1_  (.A(\V4/V4/V2/A3/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/v2 [4]));
 OR2_X1 \V4/V4/V2/A3/M1/_0_  (.A1(\V4/V4/V2/A3/M1/c1 ),
    .A2(\V4/V4/V2/A3/M1/c2 ),
    .ZN(\V4/V4/V2/A3/c1 ));
 AND2_X1 \V4/V4/V2/A3/M2/M1/_0_  (.A1(\V4/V4/V2/v4 [1]),
    .A2(\V4/V4/V2/s2 [3]),
    .ZN(\V4/V4/V2/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M2/M1/_1_  (.A(\V4/V4/V2/v4 [1]),
    .B(\V4/V4/V2/s2 [3]),
    .Z(\V4/V4/V2/A3/M2/s1 ));
 AND2_X1 \V4/V4/V2/A3/M2/M2/_0_  (.A1(\V4/V4/V2/A3/M2/s1 ),
    .A2(\V4/V4/V2/A3/c1 ),
    .ZN(\V4/V4/V2/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M2/M2/_1_  (.A(\V4/V4/V2/A3/M2/s1 ),
    .B(\V4/V4/V2/A3/c1 ),
    .Z(\V4/V4/v2 [5]));
 OR2_X1 \V4/V4/V2/A3/M2/_0_  (.A1(\V4/V4/V2/A3/M2/c1 ),
    .A2(\V4/V4/V2/A3/M2/c2 ),
    .ZN(\V4/V4/V2/A3/c2 ));
 AND2_X1 \V4/V4/V2/A3/M3/M1/_0_  (.A1(\V4/V4/V2/v4 [2]),
    .A2(\V4/V4/V2/c3 ),
    .ZN(\V4/V4/V2/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M3/M1/_1_  (.A(\V4/V4/V2/v4 [2]),
    .B(\V4/V4/V2/c3 ),
    .Z(\V4/V4/V2/A3/M3/s1 ));
 AND2_X1 \V4/V4/V2/A3/M3/M2/_0_  (.A1(\V4/V4/V2/A3/M3/s1 ),
    .A2(\V4/V4/V2/A3/c2 ),
    .ZN(\V4/V4/V2/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M3/M2/_1_  (.A(\V4/V4/V2/A3/M3/s1 ),
    .B(\V4/V4/V2/A3/c2 ),
    .Z(\V4/V4/v2 [6]));
 OR2_X1 \V4/V4/V2/A3/M3/_0_  (.A1(\V4/V4/V2/A3/M3/c1 ),
    .A2(\V4/V4/V2/A3/M3/c2 ),
    .ZN(\V4/V4/V2/A3/c3 ));
 AND2_X1 \V4/V4/V2/A3/M4/M1/_0_  (.A1(\V4/V4/V2/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V2/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V2/A3/M4/M1/_1_  (.A(\V4/V4/V2/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V2/A3/M4/s1 ));
 AND2_X1 \V4/V4/V2/A3/M4/M2/_0_  (.A1(\V4/V4/V2/A3/M4/s1 ),
    .A2(\V4/V4/V2/A3/c3 ),
    .ZN(\V4/V4/V2/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V2/A3/M4/M2/_1_  (.A(\V4/V4/V2/A3/M4/s1 ),
    .B(\V4/V4/V2/A3/c3 ),
    .Z(\V4/V4/v2 [7]));
 OR2_X1 \V4/V4/V2/A3/M4/_0_  (.A1(\V4/V4/V2/A3/M4/c1 ),
    .A2(\V4/V4/V2/A3/M4/c2 ),
    .ZN(\V4/V4/V2/overflow ));
 AND2_X1 \V4/V4/V2/V1/HA1/_0_  (.A1(\V4/V4/V2/V1/w2 ),
    .A2(\V4/V4/V2/V1/w1 ),
    .ZN(\V4/V4/V2/V1/w4 ));
 XOR2_X2 \V4/V4/V2/V1/HA1/_1_  (.A(\V4/V4/V2/V1/w2 ),
    .B(\V4/V4/V2/V1/w1 ),
    .Z(\V4/V4/v2 [1]));
 AND2_X1 \V4/V4/V2/V1/HA2/_0_  (.A1(\V4/V4/V2/V1/w4 ),
    .A2(\V4/V4/V2/V1/w3 ),
    .ZN(\V4/V4/V2/v1 [3]));
 XOR2_X2 \V4/V4/V2/V1/HA2/_1_  (.A(\V4/V4/V2/V1/w4 ),
    .B(\V4/V4/V2/V1/w3 ),
    .Z(\V4/V4/V2/v1 [2]));
 AND2_X1 \V4/V4/V2/V1/_0_  (.A1(net29),
    .A2(net14),
    .ZN(\V4/V4/v2 [0]));
 AND2_X1 \V4/V4/V2/V1/_1_  (.A1(net29),
    .A2(B[25]),
    .ZN(\V4/V4/V2/V1/w1 ));
 AND2_X1 \V4/V4/V2/V1/_2_  (.A1(net14),
    .A2(net28),
    .ZN(\V4/V4/V2/V1/w2 ));
 AND2_X1 \V4/V4/V2/V1/_3_  (.A1(B[25]),
    .A2(net28),
    .ZN(\V4/V4/V2/V1/w3 ));
 AND2_X1 \V4/V4/V2/V2/HA1/_0_  (.A1(\V4/V4/V2/V2/w2 ),
    .A2(\V4/V4/V2/V2/w1 ),
    .ZN(\V4/V4/V2/V2/w4 ));
 XOR2_X2 \V4/V4/V2/V2/HA1/_1_  (.A(\V4/V4/V2/V2/w2 ),
    .B(\V4/V4/V2/V2/w1 ),
    .Z(\V4/V4/V2/v2 [1]));
 AND2_X1 \V4/V4/V2/V2/HA2/_0_  (.A1(\V4/V4/V2/V2/w4 ),
    .A2(\V4/V4/V2/V2/w3 ),
    .ZN(\V4/V4/V2/v2 [3]));
 XOR2_X2 \V4/V4/V2/V2/HA2/_1_  (.A(\V4/V4/V2/V2/w4 ),
    .B(\V4/V4/V2/V2/w3 ),
    .Z(\V4/V4/V2/v2 [2]));
 AND2_X1 \V4/V4/V2/V2/_0_  (.A1(net27),
    .A2(net14),
    .ZN(\V4/V4/V2/v2 [0]));
 AND2_X1 \V4/V4/V2/V2/_1_  (.A1(net27),
    .A2(B[25]),
    .ZN(\V4/V4/V2/V2/w1 ));
 AND2_X1 \V4/V4/V2/V2/_2_  (.A1(net14),
    .A2(net26),
    .ZN(\V4/V4/V2/V2/w2 ));
 AND2_X1 \V4/V4/V2/V2/_3_  (.A1(B[25]),
    .A2(net26),
    .ZN(\V4/V4/V2/V2/w3 ));
 AND2_X1 \V4/V4/V2/V3/HA1/_0_  (.A1(\V4/V4/V2/V3/w2 ),
    .A2(\V4/V4/V2/V3/w1 ),
    .ZN(\V4/V4/V2/V3/w4 ));
 XOR2_X2 \V4/V4/V2/V3/HA1/_1_  (.A(\V4/V4/V2/V3/w2 ),
    .B(\V4/V4/V2/V3/w1 ),
    .Z(\V4/V4/V2/v3 [1]));
 AND2_X1 \V4/V4/V2/V3/HA2/_0_  (.A1(\V4/V4/V2/V3/w4 ),
    .A2(\V4/V4/V2/V3/w3 ),
    .ZN(\V4/V4/V2/v3 [3]));
 XOR2_X2 \V4/V4/V2/V3/HA2/_1_  (.A(\V4/V4/V2/V3/w4 ),
    .B(\V4/V4/V2/V3/w3 ),
    .Z(\V4/V4/V2/v3 [2]));
 AND2_X1 \V4/V4/V2/V3/_0_  (.A1(net29),
    .A2(net13),
    .ZN(\V4/V4/V2/v3 [0]));
 AND2_X1 \V4/V4/V2/V3/_1_  (.A1(net29),
    .A2(B[27]),
    .ZN(\V4/V4/V2/V3/w1 ));
 AND2_X1 \V4/V4/V2/V3/_2_  (.A1(net13),
    .A2(net28),
    .ZN(\V4/V4/V2/V3/w2 ));
 AND2_X1 \V4/V4/V2/V3/_3_  (.A1(B[27]),
    .A2(net28),
    .ZN(\V4/V4/V2/V3/w3 ));
 AND2_X1 \V4/V4/V2/V4/HA1/_0_  (.A1(\V4/V4/V2/V4/w2 ),
    .A2(\V4/V4/V2/V4/w1 ),
    .ZN(\V4/V4/V2/V4/w4 ));
 XOR2_X2 \V4/V4/V2/V4/HA1/_1_  (.A(\V4/V4/V2/V4/w2 ),
    .B(\V4/V4/V2/V4/w1 ),
    .Z(\V4/V4/V2/v4 [1]));
 AND2_X1 \V4/V4/V2/V4/HA2/_0_  (.A1(\V4/V4/V2/V4/w4 ),
    .A2(\V4/V4/V2/V4/w3 ),
    .ZN(\V4/V4/V2/v4 [3]));
 XOR2_X2 \V4/V4/V2/V4/HA2/_1_  (.A(\V4/V4/V2/V4/w4 ),
    .B(\V4/V4/V2/V4/w3 ),
    .Z(\V4/V4/V2/v4 [2]));
 AND2_X1 \V4/V4/V2/V4/_0_  (.A1(net27),
    .A2(net13),
    .ZN(\V4/V4/V2/v4 [0]));
 AND2_X1 \V4/V4/V2/V4/_1_  (.A1(net27),
    .A2(B[27]),
    .ZN(\V4/V4/V2/V4/w1 ));
 AND2_X1 \V4/V4/V2/V4/_2_  (.A1(net13),
    .A2(net26),
    .ZN(\V4/V4/V2/V4/w2 ));
 AND2_X1 \V4/V4/V2/V4/_3_  (.A1(B[27]),
    .A2(net26),
    .ZN(\V4/V4/V2/V4/w3 ));
 OR2_X1 \V4/V4/V2/_0_  (.A1(\V4/V4/V2/c1 ),
    .A2(\V4/V4/V2/c2 ),
    .ZN(\V4/V4/V2/c3 ));
 AND2_X1 \V4/V4/V3/A1/M1/M1/_0_  (.A1(\V4/V4/V3/v2 [0]),
    .A2(\V4/V4/V3/v3 [0]),
    .ZN(\V4/V4/V3/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M1/M1/_1_  (.A(\V4/V4/V3/v2 [0]),
    .B(\V4/V4/V3/v3 [0]),
    .Z(\V4/V4/V3/A1/M1/s1 ));
 AND2_X1 \V4/V4/V3/A1/M1/M2/_0_  (.A1(\V4/V4/V3/A1/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V3/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M1/M2/_1_  (.A(\V4/V4/V3/A1/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/V3/s1 [0]));
 OR2_X1 \V4/V4/V3/A1/M1/_0_  (.A1(\V4/V4/V3/A1/M1/c1 ),
    .A2(\V4/V4/V3/A1/M1/c2 ),
    .ZN(\V4/V4/V3/A1/c1 ));
 AND2_X1 \V4/V4/V3/A1/M2/M1/_0_  (.A1(\V4/V4/V3/v2 [1]),
    .A2(\V4/V4/V3/v3 [1]),
    .ZN(\V4/V4/V3/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M2/M1/_1_  (.A(\V4/V4/V3/v2 [1]),
    .B(\V4/V4/V3/v3 [1]),
    .Z(\V4/V4/V3/A1/M2/s1 ));
 AND2_X1 \V4/V4/V3/A1/M2/M2/_0_  (.A1(\V4/V4/V3/A1/M2/s1 ),
    .A2(\V4/V4/V3/A1/c1 ),
    .ZN(\V4/V4/V3/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M2/M2/_1_  (.A(\V4/V4/V3/A1/M2/s1 ),
    .B(\V4/V4/V3/A1/c1 ),
    .Z(\V4/V4/V3/s1 [1]));
 OR2_X1 \V4/V4/V3/A1/M2/_0_  (.A1(\V4/V4/V3/A1/M2/c1 ),
    .A2(\V4/V4/V3/A1/M2/c2 ),
    .ZN(\V4/V4/V3/A1/c2 ));
 AND2_X1 \V4/V4/V3/A1/M3/M1/_0_  (.A1(\V4/V4/V3/v2 [2]),
    .A2(\V4/V4/V3/v3 [2]),
    .ZN(\V4/V4/V3/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M3/M1/_1_  (.A(\V4/V4/V3/v2 [2]),
    .B(\V4/V4/V3/v3 [2]),
    .Z(\V4/V4/V3/A1/M3/s1 ));
 AND2_X1 \V4/V4/V3/A1/M3/M2/_0_  (.A1(\V4/V4/V3/A1/M3/s1 ),
    .A2(\V4/V4/V3/A1/c2 ),
    .ZN(\V4/V4/V3/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M3/M2/_1_  (.A(\V4/V4/V3/A1/M3/s1 ),
    .B(\V4/V4/V3/A1/c2 ),
    .Z(\V4/V4/V3/s1 [2]));
 OR2_X1 \V4/V4/V3/A1/M3/_0_  (.A1(\V4/V4/V3/A1/M3/c1 ),
    .A2(\V4/V4/V3/A1/M3/c2 ),
    .ZN(\V4/V4/V3/A1/c3 ));
 AND2_X1 \V4/V4/V3/A1/M4/M1/_0_  (.A1(\V4/V4/V3/v2 [3]),
    .A2(\V4/V4/V3/v3 [3]),
    .ZN(\V4/V4/V3/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A1/M4/M1/_1_  (.A(\V4/V4/V3/v2 [3]),
    .B(\V4/V4/V3/v3 [3]),
    .Z(\V4/V4/V3/A1/M4/s1 ));
 AND2_X1 \V4/V4/V3/A1/M4/M2/_0_  (.A1(\V4/V4/V3/A1/M4/s1 ),
    .A2(\V4/V4/V3/A1/c3 ),
    .ZN(\V4/V4/V3/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A1/M4/M2/_1_  (.A(\V4/V4/V3/A1/M4/s1 ),
    .B(\V4/V4/V3/A1/c3 ),
    .Z(\V4/V4/V3/s1 [3]));
 OR2_X1 \V4/V4/V3/A1/M4/_0_  (.A1(\V4/V4/V3/A1/M4/c1 ),
    .A2(\V4/V4/V3/A1/M4/c2 ),
    .ZN(\V4/V4/V3/c1 ));
 AND2_X1 \V4/V4/V3/A2/M1/M1/_0_  (.A1(\V4/V4/V3/s1 [0]),
    .A2(\V4/V4/V3/v1 [2]),
    .ZN(\V4/V4/V3/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M1/M1/_1_  (.A(\V4/V4/V3/s1 [0]),
    .B(\V4/V4/V3/v1 [2]),
    .Z(\V4/V4/V3/A2/M1/s1 ));
 AND2_X1 \V4/V4/V3/A2/M1/M2/_0_  (.A1(\V4/V4/V3/A2/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/V3/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M1/M2/_1_  (.A(\V4/V4/V3/A2/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/v3 [2]));
 OR2_X1 \V4/V4/V3/A2/M1/_0_  (.A1(\V4/V4/V3/A2/M1/c1 ),
    .A2(\V4/V4/V3/A2/M1/c2 ),
    .ZN(\V4/V4/V3/A2/c1 ));
 AND2_X1 \V4/V4/V3/A2/M2/M1/_0_  (.A1(\V4/V4/V3/s1 [1]),
    .A2(\V4/V4/V3/v1 [3]),
    .ZN(\V4/V4/V3/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M2/M1/_1_  (.A(\V4/V4/V3/s1 [1]),
    .B(\V4/V4/V3/v1 [3]),
    .Z(\V4/V4/V3/A2/M2/s1 ));
 AND2_X1 \V4/V4/V3/A2/M2/M2/_0_  (.A1(\V4/V4/V3/A2/M2/s1 ),
    .A2(\V4/V4/V3/A2/c1 ),
    .ZN(\V4/V4/V3/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M2/M2/_1_  (.A(\V4/V4/V3/A2/M2/s1 ),
    .B(\V4/V4/V3/A2/c1 ),
    .Z(\V4/V4/v3 [3]));
 OR2_X1 \V4/V4/V3/A2/M2/_0_  (.A1(\V4/V4/V3/A2/M2/c1 ),
    .A2(\V4/V4/V3/A2/M2/c2 ),
    .ZN(\V4/V4/V3/A2/c2 ));
 AND2_X1 \V4/V4/V3/A2/M3/M1/_0_  (.A1(\V4/V4/V3/s1 [2]),
    .A2(ground),
    .ZN(\V4/V4/V3/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M3/M1/_1_  (.A(\V4/V4/V3/s1 [2]),
    .B(ground),
    .Z(\V4/V4/V3/A2/M3/s1 ));
 AND2_X1 \V4/V4/V3/A2/M3/M2/_0_  (.A1(\V4/V4/V3/A2/M3/s1 ),
    .A2(\V4/V4/V3/A2/c2 ),
    .ZN(\V4/V4/V3/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M3/M2/_1_  (.A(\V4/V4/V3/A2/M3/s1 ),
    .B(\V4/V4/V3/A2/c2 ),
    .Z(\V4/V4/V3/s2 [2]));
 OR2_X1 \V4/V4/V3/A2/M3/_0_  (.A1(\V4/V4/V3/A2/M3/c1 ),
    .A2(\V4/V4/V3/A2/M3/c2 ),
    .ZN(\V4/V4/V3/A2/c3 ));
 AND2_X1 \V4/V4/V3/A2/M4/M1/_0_  (.A1(\V4/V4/V3/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V3/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A2/M4/M1/_1_  (.A(\V4/V4/V3/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V3/A2/M4/s1 ));
 AND2_X1 \V4/V4/V3/A2/M4/M2/_0_  (.A1(\V4/V4/V3/A2/M4/s1 ),
    .A2(\V4/V4/V3/A2/c3 ),
    .ZN(\V4/V4/V3/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A2/M4/M2/_1_  (.A(\V4/V4/V3/A2/M4/s1 ),
    .B(\V4/V4/V3/A2/c3 ),
    .Z(\V4/V4/V3/s2 [3]));
 OR2_X1 \V4/V4/V3/A2/M4/_0_  (.A1(\V4/V4/V3/A2/M4/c1 ),
    .A2(\V4/V4/V3/A2/M4/c2 ),
    .ZN(\V4/V4/V3/c2 ));
 AND2_X1 \V4/V4/V3/A3/M1/M1/_0_  (.A1(\V4/V4/V3/v4 [0]),
    .A2(\V4/V4/V3/s2 [2]),
    .ZN(\V4/V4/V3/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M1/M1/_1_  (.A(\V4/V4/V3/v4 [0]),
    .B(\V4/V4/V3/s2 [2]),
    .Z(\V4/V4/V3/A3/M1/s1 ));
 AND2_X1 \V4/V4/V3/A3/M1/M2/_0_  (.A1(\V4/V4/V3/A3/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V3/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M1/M2/_1_  (.A(\V4/V4/V3/A3/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/v3 [4]));
 OR2_X1 \V4/V4/V3/A3/M1/_0_  (.A1(\V4/V4/V3/A3/M1/c1 ),
    .A2(\V4/V4/V3/A3/M1/c2 ),
    .ZN(\V4/V4/V3/A3/c1 ));
 AND2_X1 \V4/V4/V3/A3/M2/M1/_0_  (.A1(\V4/V4/V3/v4 [1]),
    .A2(\V4/V4/V3/s2 [3]),
    .ZN(\V4/V4/V3/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M2/M1/_1_  (.A(\V4/V4/V3/v4 [1]),
    .B(\V4/V4/V3/s2 [3]),
    .Z(\V4/V4/V3/A3/M2/s1 ));
 AND2_X1 \V4/V4/V3/A3/M2/M2/_0_  (.A1(\V4/V4/V3/A3/M2/s1 ),
    .A2(\V4/V4/V3/A3/c1 ),
    .ZN(\V4/V4/V3/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M2/M2/_1_  (.A(\V4/V4/V3/A3/M2/s1 ),
    .B(\V4/V4/V3/A3/c1 ),
    .Z(\V4/V4/v3 [5]));
 OR2_X1 \V4/V4/V3/A3/M2/_0_  (.A1(\V4/V4/V3/A3/M2/c1 ),
    .A2(\V4/V4/V3/A3/M2/c2 ),
    .ZN(\V4/V4/V3/A3/c2 ));
 AND2_X1 \V4/V4/V3/A3/M3/M1/_0_  (.A1(\V4/V4/V3/v4 [2]),
    .A2(\V4/V4/V3/c3 ),
    .ZN(\V4/V4/V3/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M3/M1/_1_  (.A(\V4/V4/V3/v4 [2]),
    .B(\V4/V4/V3/c3 ),
    .Z(\V4/V4/V3/A3/M3/s1 ));
 AND2_X1 \V4/V4/V3/A3/M3/M2/_0_  (.A1(\V4/V4/V3/A3/M3/s1 ),
    .A2(\V4/V4/V3/A3/c2 ),
    .ZN(\V4/V4/V3/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M3/M2/_1_  (.A(\V4/V4/V3/A3/M3/s1 ),
    .B(\V4/V4/V3/A3/c2 ),
    .Z(\V4/V4/v3 [6]));
 OR2_X1 \V4/V4/V3/A3/M3/_0_  (.A1(\V4/V4/V3/A3/M3/c1 ),
    .A2(\V4/V4/V3/A3/M3/c2 ),
    .ZN(\V4/V4/V3/A3/c3 ));
 AND2_X1 \V4/V4/V3/A3/M4/M1/_0_  (.A1(\V4/V4/V3/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V3/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V3/A3/M4/M1/_1_  (.A(\V4/V4/V3/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V3/A3/M4/s1 ));
 AND2_X1 \V4/V4/V3/A3/M4/M2/_0_  (.A1(\V4/V4/V3/A3/M4/s1 ),
    .A2(\V4/V4/V3/A3/c3 ),
    .ZN(\V4/V4/V3/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V3/A3/M4/M2/_1_  (.A(\V4/V4/V3/A3/M4/s1 ),
    .B(\V4/V4/V3/A3/c3 ),
    .Z(\V4/V4/v3 [7]));
 OR2_X1 \V4/V4/V3/A3/M4/_0_  (.A1(\V4/V4/V3/A3/M4/c1 ),
    .A2(\V4/V4/V3/A3/M4/c2 ),
    .ZN(\V4/V4/V3/overflow ));
 AND2_X1 \V4/V4/V3/V1/HA1/_0_  (.A1(\V4/V4/V3/V1/w2 ),
    .A2(\V4/V4/V3/V1/w1 ),
    .ZN(\V4/V4/V3/V1/w4 ));
 XOR2_X2 \V4/V4/V3/V1/HA1/_1_  (.A(\V4/V4/V3/V1/w2 ),
    .B(\V4/V4/V3/V1/w1 ),
    .Z(\V4/V4/v3 [1]));
 AND2_X1 \V4/V4/V3/V1/HA2/_0_  (.A1(\V4/V4/V3/V1/w4 ),
    .A2(\V4/V4/V3/V1/w3 ),
    .ZN(\V4/V4/V3/v1 [3]));
 XOR2_X2 \V4/V4/V3/V1/HA2/_1_  (.A(\V4/V4/V3/V1/w4 ),
    .B(\V4/V4/V3/V1/w3 ),
    .Z(\V4/V4/V3/v1 [2]));
 AND2_X1 \V4/V4/V3/V1/_0_  (.A1(net33),
    .A2(B[28]),
    .ZN(\V4/V4/v3 [0]));
 AND2_X1 \V4/V4/V3/V1/_1_  (.A1(net33),
    .A2(B[29]),
    .ZN(\V4/V4/V3/V1/w1 ));
 AND2_X1 \V4/V4/V3/V1/_2_  (.A1(B[28]),
    .A2(net32),
    .ZN(\V4/V4/V3/V1/w2 ));
 AND2_X1 \V4/V4/V3/V1/_3_  (.A1(B[29]),
    .A2(net32),
    .ZN(\V4/V4/V3/V1/w3 ));
 AND2_X1 \V4/V4/V3/V2/HA1/_0_  (.A1(\V4/V4/V3/V2/w2 ),
    .A2(\V4/V4/V3/V2/w1 ),
    .ZN(\V4/V4/V3/V2/w4 ));
 XOR2_X2 \V4/V4/V3/V2/HA1/_1_  (.A(\V4/V4/V3/V2/w2 ),
    .B(\V4/V4/V3/V2/w1 ),
    .Z(\V4/V4/V3/v2 [1]));
 AND2_X1 \V4/V4/V3/V2/HA2/_0_  (.A1(\V4/V4/V3/V2/w4 ),
    .A2(\V4/V4/V3/V2/w3 ),
    .ZN(\V4/V4/V3/v2 [3]));
 XOR2_X2 \V4/V4/V3/V2/HA2/_1_  (.A(\V4/V4/V3/V2/w4 ),
    .B(\V4/V4/V3/V2/w3 ),
    .Z(\V4/V4/V3/v2 [2]));
 AND2_X1 \V4/V4/V3/V2/_0_  (.A1(net31),
    .A2(B[28]),
    .ZN(\V4/V4/V3/v2 [0]));
 AND2_X1 \V4/V4/V3/V2/_1_  (.A1(net31),
    .A2(B[29]),
    .ZN(\V4/V4/V3/V2/w1 ));
 AND2_X1 \V4/V4/V3/V2/_2_  (.A1(B[28]),
    .A2(net30),
    .ZN(\V4/V4/V3/V2/w2 ));
 AND2_X1 \V4/V4/V3/V2/_3_  (.A1(B[29]),
    .A2(net30),
    .ZN(\V4/V4/V3/V2/w3 ));
 AND2_X1 \V4/V4/V3/V3/HA1/_0_  (.A1(\V4/V4/V3/V3/w2 ),
    .A2(\V4/V4/V3/V3/w1 ),
    .ZN(\V4/V4/V3/V3/w4 ));
 XOR2_X2 \V4/V4/V3/V3/HA1/_1_  (.A(\V4/V4/V3/V3/w2 ),
    .B(\V4/V4/V3/V3/w1 ),
    .Z(\V4/V4/V3/v3 [1]));
 AND2_X1 \V4/V4/V3/V3/HA2/_0_  (.A1(\V4/V4/V3/V3/w4 ),
    .A2(\V4/V4/V3/V3/w3 ),
    .ZN(\V4/V4/V3/v3 [3]));
 XOR2_X2 \V4/V4/V3/V3/HA2/_1_  (.A(\V4/V4/V3/V3/w4 ),
    .B(\V4/V4/V3/V3/w3 ),
    .Z(\V4/V4/V3/v3 [2]));
 AND2_X1 \V4/V4/V3/V3/_0_  (.A1(net33),
    .A2(B[30]),
    .ZN(\V4/V4/V3/v3 [0]));
 AND2_X1 \V4/V4/V3/V3/_1_  (.A1(net33),
    .A2(B[31]),
    .ZN(\V4/V4/V3/V3/w1 ));
 AND2_X1 \V4/V4/V3/V3/_2_  (.A1(B[30]),
    .A2(net32),
    .ZN(\V4/V4/V3/V3/w2 ));
 AND2_X1 \V4/V4/V3/V3/_3_  (.A1(B[31]),
    .A2(net32),
    .ZN(\V4/V4/V3/V3/w3 ));
 AND2_X1 \V4/V4/V3/V4/HA1/_0_  (.A1(\V4/V4/V3/V4/w2 ),
    .A2(\V4/V4/V3/V4/w1 ),
    .ZN(\V4/V4/V3/V4/w4 ));
 XOR2_X2 \V4/V4/V3/V4/HA1/_1_  (.A(\V4/V4/V3/V4/w2 ),
    .B(\V4/V4/V3/V4/w1 ),
    .Z(\V4/V4/V3/v4 [1]));
 AND2_X1 \V4/V4/V3/V4/HA2/_0_  (.A1(\V4/V4/V3/V4/w4 ),
    .A2(\V4/V4/V3/V4/w3 ),
    .ZN(\V4/V4/V3/v4 [3]));
 XOR2_X2 \V4/V4/V3/V4/HA2/_1_  (.A(\V4/V4/V3/V4/w4 ),
    .B(\V4/V4/V3/V4/w3 ),
    .Z(\V4/V4/V3/v4 [2]));
 AND2_X1 \V4/V4/V3/V4/_0_  (.A1(net31),
    .A2(B[30]),
    .ZN(\V4/V4/V3/v4 [0]));
 AND2_X1 \V4/V4/V3/V4/_1_  (.A1(net31),
    .A2(B[31]),
    .ZN(\V4/V4/V3/V4/w1 ));
 AND2_X1 \V4/V4/V3/V4/_2_  (.A1(B[30]),
    .A2(net30),
    .ZN(\V4/V4/V3/V4/w2 ));
 AND2_X1 \V4/V4/V3/V4/_3_  (.A1(B[31]),
    .A2(net30),
    .ZN(\V4/V4/V3/V4/w3 ));
 OR2_X1 \V4/V4/V3/_0_  (.A1(\V4/V4/V3/c1 ),
    .A2(\V4/V4/V3/c2 ),
    .ZN(\V4/V4/V3/c3 ));
 AND2_X1 \V4/V4/V4/A1/M1/M1/_0_  (.A1(\V4/V4/V4/v2 [0]),
    .A2(\V4/V4/V4/v3 [0]),
    .ZN(\V4/V4/V4/A1/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M1/M1/_1_  (.A(\V4/V4/V4/v2 [0]),
    .B(\V4/V4/V4/v3 [0]),
    .Z(\V4/V4/V4/A1/M1/s1 ));
 AND2_X1 \V4/V4/V4/A1/M1/M2/_0_  (.A1(\V4/V4/V4/A1/M1/s1 ),
    .A2(net9),
    .ZN(\V4/V4/V4/A1/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M1/M2/_1_  (.A(\V4/V4/V4/A1/M1/s1 ),
    .B(net9),
    .Z(\V4/V4/V4/s1 [0]));
 OR2_X1 \V4/V4/V4/A1/M1/_0_  (.A1(\V4/V4/V4/A1/M1/c1 ),
    .A2(\V4/V4/V4/A1/M1/c2 ),
    .ZN(\V4/V4/V4/A1/c1 ));
 AND2_X1 \V4/V4/V4/A1/M2/M1/_0_  (.A1(\V4/V4/V4/v2 [1]),
    .A2(\V4/V4/V4/v3 [1]),
    .ZN(\V4/V4/V4/A1/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M2/M1/_1_  (.A(\V4/V4/V4/v2 [1]),
    .B(\V4/V4/V4/v3 [1]),
    .Z(\V4/V4/V4/A1/M2/s1 ));
 AND2_X1 \V4/V4/V4/A1/M2/M2/_0_  (.A1(\V4/V4/V4/A1/M2/s1 ),
    .A2(\V4/V4/V4/A1/c1 ),
    .ZN(\V4/V4/V4/A1/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M2/M2/_1_  (.A(\V4/V4/V4/A1/M2/s1 ),
    .B(\V4/V4/V4/A1/c1 ),
    .Z(\V4/V4/V4/s1 [1]));
 OR2_X1 \V4/V4/V4/A1/M2/_0_  (.A1(\V4/V4/V4/A1/M2/c1 ),
    .A2(\V4/V4/V4/A1/M2/c2 ),
    .ZN(\V4/V4/V4/A1/c2 ));
 AND2_X1 \V4/V4/V4/A1/M3/M1/_0_  (.A1(\V4/V4/V4/v2 [2]),
    .A2(\V4/V4/V4/v3 [2]),
    .ZN(\V4/V4/V4/A1/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M3/M1/_1_  (.A(\V4/V4/V4/v2 [2]),
    .B(\V4/V4/V4/v3 [2]),
    .Z(\V4/V4/V4/A1/M3/s1 ));
 AND2_X1 \V4/V4/V4/A1/M3/M2/_0_  (.A1(\V4/V4/V4/A1/M3/s1 ),
    .A2(\V4/V4/V4/A1/c2 ),
    .ZN(\V4/V4/V4/A1/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M3/M2/_1_  (.A(\V4/V4/V4/A1/M3/s1 ),
    .B(\V4/V4/V4/A1/c2 ),
    .Z(\V4/V4/V4/s1 [2]));
 OR2_X1 \V4/V4/V4/A1/M3/_0_  (.A1(\V4/V4/V4/A1/M3/c1 ),
    .A2(\V4/V4/V4/A1/M3/c2 ),
    .ZN(\V4/V4/V4/A1/c3 ));
 AND2_X1 \V4/V4/V4/A1/M4/M1/_0_  (.A1(\V4/V4/V4/v2 [3]),
    .A2(\V4/V4/V4/v3 [3]),
    .ZN(\V4/V4/V4/A1/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A1/M4/M1/_1_  (.A(\V4/V4/V4/v2 [3]),
    .B(\V4/V4/V4/v3 [3]),
    .Z(\V4/V4/V4/A1/M4/s1 ));
 AND2_X1 \V4/V4/V4/A1/M4/M2/_0_  (.A1(\V4/V4/V4/A1/M4/s1 ),
    .A2(\V4/V4/V4/A1/c3 ),
    .ZN(\V4/V4/V4/A1/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A1/M4/M2/_1_  (.A(\V4/V4/V4/A1/M4/s1 ),
    .B(\V4/V4/V4/A1/c3 ),
    .Z(\V4/V4/V4/s1 [3]));
 OR2_X1 \V4/V4/V4/A1/M4/_0_  (.A1(\V4/V4/V4/A1/M4/c1 ),
    .A2(\V4/V4/V4/A1/M4/c2 ),
    .ZN(\V4/V4/V4/c1 ));
 AND2_X1 \V4/V4/V4/A2/M1/M1/_0_  (.A1(\V4/V4/V4/s1 [0]),
    .A2(\V4/V4/V4/v1 [2]),
    .ZN(\V4/V4/V4/A2/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M1/M1/_1_  (.A(\V4/V4/V4/s1 [0]),
    .B(\V4/V4/V4/v1 [2]),
    .Z(\V4/V4/V4/A2/M1/s1 ));
 AND2_X1 \V4/V4/V4/A2/M1/M2/_0_  (.A1(\V4/V4/V4/A2/M1/s1 ),
    .A2(ground),
    .ZN(\V4/V4/V4/A2/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M1/M2/_1_  (.A(\V4/V4/V4/A2/M1/s1 ),
    .B(ground),
    .Z(\V4/V4/v4 [2]));
 OR2_X1 \V4/V4/V4/A2/M1/_0_  (.A1(\V4/V4/V4/A2/M1/c1 ),
    .A2(\V4/V4/V4/A2/M1/c2 ),
    .ZN(\V4/V4/V4/A2/c1 ));
 AND2_X1 \V4/V4/V4/A2/M2/M1/_0_  (.A1(\V4/V4/V4/s1 [1]),
    .A2(\V4/V4/V4/v1 [3]),
    .ZN(\V4/V4/V4/A2/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M2/M1/_1_  (.A(\V4/V4/V4/s1 [1]),
    .B(\V4/V4/V4/v1 [3]),
    .Z(\V4/V4/V4/A2/M2/s1 ));
 AND2_X1 \V4/V4/V4/A2/M2/M2/_0_  (.A1(\V4/V4/V4/A2/M2/s1 ),
    .A2(\V4/V4/V4/A2/c1 ),
    .ZN(\V4/V4/V4/A2/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M2/M2/_1_  (.A(\V4/V4/V4/A2/M2/s1 ),
    .B(\V4/V4/V4/A2/c1 ),
    .Z(\V4/V4/v4 [3]));
 OR2_X1 \V4/V4/V4/A2/M2/_0_  (.A1(\V4/V4/V4/A2/M2/c1 ),
    .A2(\V4/V4/V4/A2/M2/c2 ),
    .ZN(\V4/V4/V4/A2/c2 ));
 AND2_X1 \V4/V4/V4/A2/M3/M1/_0_  (.A1(\V4/V4/V4/s1 [2]),
    .A2(net10),
    .ZN(\V4/V4/V4/A2/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M3/M1/_1_  (.A(\V4/V4/V4/s1 [2]),
    .B(net10),
    .Z(\V4/V4/V4/A2/M3/s1 ));
 AND2_X1 \V4/V4/V4/A2/M3/M2/_0_  (.A1(\V4/V4/V4/A2/M3/s1 ),
    .A2(\V4/V4/V4/A2/c2 ),
    .ZN(\V4/V4/V4/A2/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M3/M2/_1_  (.A(\V4/V4/V4/A2/M3/s1 ),
    .B(\V4/V4/V4/A2/c2 ),
    .Z(\V4/V4/V4/s2 [2]));
 OR2_X1 \V4/V4/V4/A2/M3/_0_  (.A1(\V4/V4/V4/A2/M3/c1 ),
    .A2(\V4/V4/V4/A2/M3/c2 ),
    .ZN(\V4/V4/V4/A2/c3 ));
 AND2_X1 \V4/V4/V4/A2/M4/M1/_0_  (.A1(\V4/V4/V4/s1 [3]),
    .A2(ground),
    .ZN(\V4/V4/V4/A2/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A2/M4/M1/_1_  (.A(\V4/V4/V4/s1 [3]),
    .B(ground),
    .Z(\V4/V4/V4/A2/M4/s1 ));
 AND2_X1 \V4/V4/V4/A2/M4/M2/_0_  (.A1(\V4/V4/V4/A2/M4/s1 ),
    .A2(\V4/V4/V4/A2/c3 ),
    .ZN(\V4/V4/V4/A2/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A2/M4/M2/_1_  (.A(\V4/V4/V4/A2/M4/s1 ),
    .B(\V4/V4/V4/A2/c3 ),
    .Z(\V4/V4/V4/s2 [3]));
 OR2_X1 \V4/V4/V4/A2/M4/_0_  (.A1(\V4/V4/V4/A2/M4/c1 ),
    .A2(\V4/V4/V4/A2/M4/c2 ),
    .ZN(\V4/V4/V4/c2 ));
 AND2_X1 \V4/V4/V4/A3/M1/M1/_0_  (.A1(\V4/V4/V4/v4 [0]),
    .A2(\V4/V4/V4/s2 [2]),
    .ZN(\V4/V4/V4/A3/M1/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M1/M1/_1_  (.A(\V4/V4/V4/v4 [0]),
    .B(\V4/V4/V4/s2 [2]),
    .Z(\V4/V4/V4/A3/M1/s1 ));
 AND2_X1 \V4/V4/V4/A3/M1/M2/_0_  (.A1(\V4/V4/V4/A3/M1/s1 ),
    .A2(net10),
    .ZN(\V4/V4/V4/A3/M1/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M1/M2/_1_  (.A(\V4/V4/V4/A3/M1/s1 ),
    .B(net10),
    .Z(\V4/V4/v4 [4]));
 OR2_X1 \V4/V4/V4/A3/M1/_0_  (.A1(\V4/V4/V4/A3/M1/c1 ),
    .A2(\V4/V4/V4/A3/M1/c2 ),
    .ZN(\V4/V4/V4/A3/c1 ));
 AND2_X1 \V4/V4/V4/A3/M2/M1/_0_  (.A1(\V4/V4/V4/v4 [1]),
    .A2(\V4/V4/V4/s2 [3]),
    .ZN(\V4/V4/V4/A3/M2/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M2/M1/_1_  (.A(\V4/V4/V4/v4 [1]),
    .B(\V4/V4/V4/s2 [3]),
    .Z(\V4/V4/V4/A3/M2/s1 ));
 AND2_X1 \V4/V4/V4/A3/M2/M2/_0_  (.A1(\V4/V4/V4/A3/M2/s1 ),
    .A2(\V4/V4/V4/A3/c1 ),
    .ZN(\V4/V4/V4/A3/M2/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M2/M2/_1_  (.A(\V4/V4/V4/A3/M2/s1 ),
    .B(\V4/V4/V4/A3/c1 ),
    .Z(\V4/V4/v4 [5]));
 OR2_X1 \V4/V4/V4/A3/M2/_0_  (.A1(\V4/V4/V4/A3/M2/c1 ),
    .A2(\V4/V4/V4/A3/M2/c2 ),
    .ZN(\V4/V4/V4/A3/c2 ));
 AND2_X1 \V4/V4/V4/A3/M3/M1/_0_  (.A1(\V4/V4/V4/v4 [2]),
    .A2(\V4/V4/V4/c3 ),
    .ZN(\V4/V4/V4/A3/M3/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M3/M1/_1_  (.A(\V4/V4/V4/v4 [2]),
    .B(\V4/V4/V4/c3 ),
    .Z(\V4/V4/V4/A3/M3/s1 ));
 AND2_X1 \V4/V4/V4/A3/M3/M2/_0_  (.A1(\V4/V4/V4/A3/M3/s1 ),
    .A2(\V4/V4/V4/A3/c2 ),
    .ZN(\V4/V4/V4/A3/M3/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M3/M2/_1_  (.A(\V4/V4/V4/A3/M3/s1 ),
    .B(\V4/V4/V4/A3/c2 ),
    .Z(\V4/V4/v4 [6]));
 OR2_X1 \V4/V4/V4/A3/M3/_0_  (.A1(\V4/V4/V4/A3/M3/c1 ),
    .A2(\V4/V4/V4/A3/M3/c2 ),
    .ZN(\V4/V4/V4/A3/c3 ));
 AND2_X1 \V4/V4/V4/A3/M4/M1/_0_  (.A1(\V4/V4/V4/v4 [3]),
    .A2(ground),
    .ZN(\V4/V4/V4/A3/M4/c1 ));
 XOR2_X2 \V4/V4/V4/A3/M4/M1/_1_  (.A(\V4/V4/V4/v4 [3]),
    .B(ground),
    .Z(\V4/V4/V4/A3/M4/s1 ));
 AND2_X1 \V4/V4/V4/A3/M4/M2/_0_  (.A1(\V4/V4/V4/A3/M4/s1 ),
    .A2(\V4/V4/V4/A3/c3 ),
    .ZN(\V4/V4/V4/A3/M4/c2 ));
 XOR2_X2 \V4/V4/V4/A3/M4/M2/_1_  (.A(\V4/V4/V4/A3/M4/s1 ),
    .B(\V4/V4/V4/A3/c3 ),
    .Z(\V4/V4/v4 [7]));
 OR2_X1 \V4/V4/V4/A3/M4/_0_  (.A1(\V4/V4/V4/A3/M4/c1 ),
    .A2(\V4/V4/V4/A3/M4/c2 ),
    .ZN(\V4/V4/V4/overflow ));
 AND2_X1 \V4/V4/V4/V1/HA1/_0_  (.A1(\V4/V4/V4/V1/w2 ),
    .A2(\V4/V4/V4/V1/w1 ),
    .ZN(\V4/V4/V4/V1/w4 ));
 XOR2_X2 \V4/V4/V4/V1/HA1/_1_  (.A(\V4/V4/V4/V1/w2 ),
    .B(\V4/V4/V4/V1/w1 ),
    .Z(\V4/V4/v4 [1]));
 AND2_X1 \V4/V4/V4/V1/HA2/_0_  (.A1(\V4/V4/V4/V1/w4 ),
    .A2(\V4/V4/V4/V1/w3 ),
    .ZN(\V4/V4/V4/v1 [3]));
 XOR2_X2 \V4/V4/V4/V1/HA2/_1_  (.A(\V4/V4/V4/V1/w4 ),
    .B(\V4/V4/V4/V1/w3 ),
    .Z(\V4/V4/V4/v1 [2]));
 AND2_X1 \V4/V4/V4/V1/_0_  (.A1(net29),
    .A2(B[28]),
    .ZN(\V4/V4/v4 [0]));
 AND2_X1 \V4/V4/V4/V1/_1_  (.A1(net29),
    .A2(B[29]),
    .ZN(\V4/V4/V4/V1/w1 ));
 AND2_X1 \V4/V4/V4/V1/_2_  (.A1(B[28]),
    .A2(net28),
    .ZN(\V4/V4/V4/V1/w2 ));
 AND2_X1 \V4/V4/V4/V1/_3_  (.A1(B[29]),
    .A2(net28),
    .ZN(\V4/V4/V4/V1/w3 ));
 AND2_X1 \V4/V4/V4/V2/HA1/_0_  (.A1(\V4/V4/V4/V2/w2 ),
    .A2(\V4/V4/V4/V2/w1 ),
    .ZN(\V4/V4/V4/V2/w4 ));
 XOR2_X2 \V4/V4/V4/V2/HA1/_1_  (.A(\V4/V4/V4/V2/w2 ),
    .B(\V4/V4/V4/V2/w1 ),
    .Z(\V4/V4/V4/v2 [1]));
 AND2_X1 \V4/V4/V4/V2/HA2/_0_  (.A1(\V4/V4/V4/V2/w4 ),
    .A2(\V4/V4/V4/V2/w3 ),
    .ZN(\V4/V4/V4/v2 [3]));
 XOR2_X2 \V4/V4/V4/V2/HA2/_1_  (.A(\V4/V4/V4/V2/w4 ),
    .B(\V4/V4/V4/V2/w3 ),
    .Z(\V4/V4/V4/v2 [2]));
 AND2_X1 \V4/V4/V4/V2/_0_  (.A1(net27),
    .A2(B[28]),
    .ZN(\V4/V4/V4/v2 [0]));
 AND2_X1 \V4/V4/V4/V2/_1_  (.A1(net27),
    .A2(B[29]),
    .ZN(\V4/V4/V4/V2/w1 ));
 AND2_X1 \V4/V4/V4/V2/_2_  (.A1(B[28]),
    .A2(net26),
    .ZN(\V4/V4/V4/V2/w2 ));
 AND2_X1 \V4/V4/V4/V2/_3_  (.A1(B[29]),
    .A2(net26),
    .ZN(\V4/V4/V4/V2/w3 ));
 AND2_X1 \V4/V4/V4/V3/HA1/_0_  (.A1(\V4/V4/V4/V3/w2 ),
    .A2(\V4/V4/V4/V3/w1 ),
    .ZN(\V4/V4/V4/V3/w4 ));
 XOR2_X2 \V4/V4/V4/V3/HA1/_1_  (.A(\V4/V4/V4/V3/w2 ),
    .B(\V4/V4/V4/V3/w1 ),
    .Z(\V4/V4/V4/v3 [1]));
 AND2_X1 \V4/V4/V4/V3/HA2/_0_  (.A1(\V4/V4/V4/V3/w4 ),
    .A2(\V4/V4/V4/V3/w3 ),
    .ZN(\V4/V4/V4/v3 [3]));
 XOR2_X2 \V4/V4/V4/V3/HA2/_1_  (.A(\V4/V4/V4/V3/w4 ),
    .B(\V4/V4/V4/V3/w3 ),
    .Z(\V4/V4/V4/v3 [2]));
 AND2_X1 \V4/V4/V4/V3/_0_  (.A1(net29),
    .A2(B[30]),
    .ZN(\V4/V4/V4/v3 [0]));
 AND2_X1 \V4/V4/V4/V3/_1_  (.A1(net29),
    .A2(B[31]),
    .ZN(\V4/V4/V4/V3/w1 ));
 AND2_X1 \V4/V4/V4/V3/_2_  (.A1(B[30]),
    .A2(net28),
    .ZN(\V4/V4/V4/V3/w2 ));
 AND2_X1 \V4/V4/V4/V3/_3_  (.A1(B[31]),
    .A2(net28),
    .ZN(\V4/V4/V4/V3/w3 ));
 AND2_X1 \V4/V4/V4/V4/HA1/_0_  (.A1(\V4/V4/V4/V4/w2 ),
    .A2(\V4/V4/V4/V4/w1 ),
    .ZN(\V4/V4/V4/V4/w4 ));
 XOR2_X2 \V4/V4/V4/V4/HA1/_1_  (.A(\V4/V4/V4/V4/w2 ),
    .B(\V4/V4/V4/V4/w1 ),
    .Z(\V4/V4/V4/v4 [1]));
 AND2_X1 \V4/V4/V4/V4/HA2/_0_  (.A1(\V4/V4/V4/V4/w4 ),
    .A2(\V4/V4/V4/V4/w3 ),
    .ZN(\V4/V4/V4/v4 [3]));
 XOR2_X2 \V4/V4/V4/V4/HA2/_1_  (.A(\V4/V4/V4/V4/w4 ),
    .B(\V4/V4/V4/V4/w3 ),
    .Z(\V4/V4/V4/v4 [2]));
 AND2_X1 \V4/V4/V4/V4/_0_  (.A1(net27),
    .A2(B[30]),
    .ZN(\V4/V4/V4/v4 [0]));
 AND2_X1 \V4/V4/V4/V4/_1_  (.A1(net27),
    .A2(B[31]),
    .ZN(\V4/V4/V4/V4/w1 ));
 AND2_X1 \V4/V4/V4/V4/_2_  (.A1(B[30]),
    .A2(net26),
    .ZN(\V4/V4/V4/V4/w2 ));
 AND2_X1 \V4/V4/V4/V4/_3_  (.A1(B[31]),
    .A2(net26),
    .ZN(\V4/V4/V4/V4/w3 ));
 OR2_X1 \V4/V4/V4/_0_  (.A1(\V4/V4/V4/c1 ),
    .A2(\V4/V4/V4/c2 ),
    .ZN(\V4/V4/V4/c3 ));
 OR2_X1 \V4/V4/_0_  (.A1(\V4/V4/c1 ),
    .A2(\V4/V4/c2 ),
    .ZN(\V4/V4/c3 ));
 OR2_X1 \V4/_0_  (.A1(\V4/c1 ),
    .A2(\V4/c2 ),
    .ZN(\V4/c3 ));
 OR2_X2 _0_ (.A1(c1),
    .A2(c2),
    .ZN(c3));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Right_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Right_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Right_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Right_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Right_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Right_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Right_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Right_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Right_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Right_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Right_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Right_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Right_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Right_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Right_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Right_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Right_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Right_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Right_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Right_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Right_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Right_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Right_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Right_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Right_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Right_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Right_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Right_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_353_Right_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_354_Right_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_355_Right_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_356_Right_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_357_Right_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_358_Right_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_359_Right_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_360_Right_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_361_Right_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_362_Right_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_363_Right_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_364_Right_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_365_Right_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_366_Right_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_367_Right_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_368_Right_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_369_Right_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_370_Right_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_371_Right_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_372_Right_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_373_Right_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_374_Right_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_375_Right_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_376_Right_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_377_Right_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_378_Right_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_379_Right_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_380_Right_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_381_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_382_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_383_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_384_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_385_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_386_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_387_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_388_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_389_Right_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_390_Right_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_391_Right_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_392_Right_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_393_Right_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_394_Right_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_395_Right_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_396_Right_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_397_Right_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_398_Right_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_399_Right_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_400_Right_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_401_Right_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_402_Right_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_403_Right_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_404_Right_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_405_Right_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_406_Right_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_407_Right_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_408_Right_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_409_Right_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_410_Right_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_411_Right_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_412_Right_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_413_Right_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_414_Right_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_415_Right_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_416_Right_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_417_Right_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_418_Right_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_419_Right_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_420_Right_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_421_Right_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_422_Right_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_423_Right_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_424_Right_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_425_Right_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_426_Right_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_427_Right_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_428_Right_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_429_Right_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_430_Right_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_431_Right_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_432_Right_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_433_Right_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_434_Right_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_435_Right_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_436_Right_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_437_Right_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_438_Right_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_439_Right_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_440_Right_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_441_Right_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_442_Right_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_443_Right_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_444_Right_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_445_Right_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_446_Right_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_447_Right_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_448_Right_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_449_Right_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_450_Right_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_451_Right_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_452_Right_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_453_Right_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_454_Right_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_455_Right_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_456_Right_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_457_Right_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_458_Right_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_459_Right_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_460_Right_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_461_Right_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_462_Right_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_463_Right_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_464_Right_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_465_Right_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_466_Right_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_467_Right_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_468_Right_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_469_Right_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_470_Right_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_471_Right_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_472_Right_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_473_Right_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_474_Right_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_475_Right_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_476_Right_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_477_Right_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_478_Right_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_479_Right_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_480_Right_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_481_Right_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_482_Right_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_483_Right_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_484_Right_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_485_Right_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_486_Right_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_487_Right_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_488_Right_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_489_Right_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_490_Right_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_491_Right_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_492_Right_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_493_Right_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_494_Right_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_495_Right_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_496_Right_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_497_Right_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_498_Right_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_499_Right_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_500_Right_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_501_Right_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_502_Right_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_503_Right_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_504_Right_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_505_Right_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_506_Right_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_507_Right_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_508_Right_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_509_Right_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_510_Right_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_511_Right_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_512_Right_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_513_Right_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_514_Right_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_515_Right_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_516_Right_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_517_Right_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_518_Right_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_519_Right_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_520_Right_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_521_Right_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_522_Right_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_523_Right_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_524_Right_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_525_Right_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_526_Right_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_527_Right_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_528_Right_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_529_Right_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_530_Right_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_531_Right_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_532_Right_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_533_Right_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_534_Right_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_535_Right_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_536_Right_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_537_Right_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_538_Right_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_539_Right_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_540_Right_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_541_Right_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_542_Right_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_543_Right_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_544_Right_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_545_Right_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_546_Right_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_547_Right_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_548_Right_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_549_Right_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_550_Right_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_551_Right_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_552_Right_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_553_Right_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_554_Right_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_555_Right_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_556_Right_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_557_Right_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_558_Right_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_559_Right_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_560_Right_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_561_Right_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_562_Right_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_563_Right_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_564_Right_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_565_Right_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_566_Right_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_567_Right_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_568_Right_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_569_Right_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_570_Right_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_571_Right_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_572_Right_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_573_Right_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_574_Right_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_575_Right_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_576_Right_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_577_Right_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_578_Right_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_579_Right_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_580_Right_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_581_Right_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_582_Right_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_583_Right_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_584_Right_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_585_Right_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_586_Right_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_587_Right_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_588_Right_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_589_Right_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_590_Right_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_591_Right_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_592_Right_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_593_Right_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_594_Right_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_595_Right_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_596_Right_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_597_Right_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_598_Right_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_599_Right_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_600_Right_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_601_Right_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_602_Right_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_603_Right_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_604_Right_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_605_Right_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_606_Right_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_607_Right_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_608_Right_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_609_Right_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_610_Right_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_611_Right_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_612_Right_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_613_Right_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_614_Right_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_615_Right_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_616_Right_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_617_Right_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_618_Right_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_619_Right_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_620_Right_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_621_Right_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_622_Right_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_623_Right_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_624_Right_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_625_Right_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_626_Right_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_627_Right_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_628_Right_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_629_Right_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_630_Right_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_631_Right_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_632_Right_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_633_Right_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_634_Right_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_635_Right_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_636_Right_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_637_Right_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_638_Right_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_639_Right_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_640_Right_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_641_Right_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_642_Right_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_643_Right_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_644_Right_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_645_Right_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_646_Right_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_647_Right_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_648_Right_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_649_Right_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_650_Right_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_651_Right_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_652_Right_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_653_Right_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_654_Right_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_655_Right_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_656_Right_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_657_Right_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_658_Right_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_659_Right_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_660_Right_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_661_Right_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_662_Right_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_663_Right_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_664_Right_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_665_Right_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_666_Right_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_667_Right_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_668_Right_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_669_Right_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_670_Right_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_671_Right_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_672_Right_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_673_Right_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_674_Right_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_675_Right_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_676_Right_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_795 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_796 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_797 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_798 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_799 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_800 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_801 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_802 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_803 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_804 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_805 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_806 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_807 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_808 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_809 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_810 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_811 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_812 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_813 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_814 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_815 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_816 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_817 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_818 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_819 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_820 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_821 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_822 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_823 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_824 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_825 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_826 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_827 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_828 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_829 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_830 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_831 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_832 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_833 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_834 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_835 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_836 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_837 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_838 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_839 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_840 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_841 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_842 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_843 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_844 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_845 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_846 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_847 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_848 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_849 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_850 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_851 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_852 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_853 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_854 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_855 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_856 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_857 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_858 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_859 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_860 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_861 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_862 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_863 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_864 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_865 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_866 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_867 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_868 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_869 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_870 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_871 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_872 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_873 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_874 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_875 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_876 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_877 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_878 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_879 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_880 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_881 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_882 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_883 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_884 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_885 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_886 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_887 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_888 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_889 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_890 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_891 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_892 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_893 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_894 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_895 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_896 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_897 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_898 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_899 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_900 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_901 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_902 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_903 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_904 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_905 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_906 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_907 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_908 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_909 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_910 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_911 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_912 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_913 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_914 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_915 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_916 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_917 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_918 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_919 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_920 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_921 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_922 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_923 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_924 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_925 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_926 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_927 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_928 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_929 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_930 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_931 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_932 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_933 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Left_934 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Left_935 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Left_936 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Left_937 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Left_938 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Left_939 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Left_940 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Left_941 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Left_942 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Left_943 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Left_944 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Left_945 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Left_946 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Left_947 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Left_948 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Left_949 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Left_950 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Left_951 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Left_952 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Left_953 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Left_954 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Left_955 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Left_956 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Left_957 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Left_958 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Left_959 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Left_960 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Left_961 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Left_962 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Left_963 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Left_964 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Left_965 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Left_966 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Left_967 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Left_968 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Left_969 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Left_970 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Left_971 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Left_972 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Left_973 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Left_974 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Left_975 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Left_976 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Left_977 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Left_978 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Left_979 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Left_980 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Left_981 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Left_982 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Left_983 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Left_984 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Left_985 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Left_986 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Left_987 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Left_988 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Left_989 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Left_990 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Left_991 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Left_992 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Left_993 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Left_994 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Left_995 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Left_996 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Left_997 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Left_998 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Left_999 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Left_1000 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Left_1001 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Left_1002 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Left_1003 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Left_1004 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Left_1005 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Left_1006 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Left_1007 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Left_1008 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Left_1009 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Left_1010 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Left_1011 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Left_1012 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Left_1013 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Left_1014 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Left_1015 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Left_1016 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Left_1017 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Left_1018 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Left_1019 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Left_1020 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Left_1021 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Left_1022 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Left_1023 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Left_1024 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Left_1025 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Left_1026 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Left_1027 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Left_1028 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Left_1029 ();
 TAPCELL_X1 PHY_EDGE_ROW_353_Left_1030 ();
 TAPCELL_X1 PHY_EDGE_ROW_354_Left_1031 ();
 TAPCELL_X1 PHY_EDGE_ROW_355_Left_1032 ();
 TAPCELL_X1 PHY_EDGE_ROW_356_Left_1033 ();
 TAPCELL_X1 PHY_EDGE_ROW_357_Left_1034 ();
 TAPCELL_X1 PHY_EDGE_ROW_358_Left_1035 ();
 TAPCELL_X1 PHY_EDGE_ROW_359_Left_1036 ();
 TAPCELL_X1 PHY_EDGE_ROW_360_Left_1037 ();
 TAPCELL_X1 PHY_EDGE_ROW_361_Left_1038 ();
 TAPCELL_X1 PHY_EDGE_ROW_362_Left_1039 ();
 TAPCELL_X1 PHY_EDGE_ROW_363_Left_1040 ();
 TAPCELL_X1 PHY_EDGE_ROW_364_Left_1041 ();
 TAPCELL_X1 PHY_EDGE_ROW_365_Left_1042 ();
 TAPCELL_X1 PHY_EDGE_ROW_366_Left_1043 ();
 TAPCELL_X1 PHY_EDGE_ROW_367_Left_1044 ();
 TAPCELL_X1 PHY_EDGE_ROW_368_Left_1045 ();
 TAPCELL_X1 PHY_EDGE_ROW_369_Left_1046 ();
 TAPCELL_X1 PHY_EDGE_ROW_370_Left_1047 ();
 TAPCELL_X1 PHY_EDGE_ROW_371_Left_1048 ();
 TAPCELL_X1 PHY_EDGE_ROW_372_Left_1049 ();
 TAPCELL_X1 PHY_EDGE_ROW_373_Left_1050 ();
 TAPCELL_X1 PHY_EDGE_ROW_374_Left_1051 ();
 TAPCELL_X1 PHY_EDGE_ROW_375_Left_1052 ();
 TAPCELL_X1 PHY_EDGE_ROW_376_Left_1053 ();
 TAPCELL_X1 PHY_EDGE_ROW_377_Left_1054 ();
 TAPCELL_X1 PHY_EDGE_ROW_378_Left_1055 ();
 TAPCELL_X1 PHY_EDGE_ROW_379_Left_1056 ();
 TAPCELL_X1 PHY_EDGE_ROW_380_Left_1057 ();
 TAPCELL_X1 PHY_EDGE_ROW_381_Left_1058 ();
 TAPCELL_X1 PHY_EDGE_ROW_382_Left_1059 ();
 TAPCELL_X1 PHY_EDGE_ROW_383_Left_1060 ();
 TAPCELL_X1 PHY_EDGE_ROW_384_Left_1061 ();
 TAPCELL_X1 PHY_EDGE_ROW_385_Left_1062 ();
 TAPCELL_X1 PHY_EDGE_ROW_386_Left_1063 ();
 TAPCELL_X1 PHY_EDGE_ROW_387_Left_1064 ();
 TAPCELL_X1 PHY_EDGE_ROW_388_Left_1065 ();
 TAPCELL_X1 PHY_EDGE_ROW_389_Left_1066 ();
 TAPCELL_X1 PHY_EDGE_ROW_390_Left_1067 ();
 TAPCELL_X1 PHY_EDGE_ROW_391_Left_1068 ();
 TAPCELL_X1 PHY_EDGE_ROW_392_Left_1069 ();
 TAPCELL_X1 PHY_EDGE_ROW_393_Left_1070 ();
 TAPCELL_X1 PHY_EDGE_ROW_394_Left_1071 ();
 TAPCELL_X1 PHY_EDGE_ROW_395_Left_1072 ();
 TAPCELL_X1 PHY_EDGE_ROW_396_Left_1073 ();
 TAPCELL_X1 PHY_EDGE_ROW_397_Left_1074 ();
 TAPCELL_X1 PHY_EDGE_ROW_398_Left_1075 ();
 TAPCELL_X1 PHY_EDGE_ROW_399_Left_1076 ();
 TAPCELL_X1 PHY_EDGE_ROW_400_Left_1077 ();
 TAPCELL_X1 PHY_EDGE_ROW_401_Left_1078 ();
 TAPCELL_X1 PHY_EDGE_ROW_402_Left_1079 ();
 TAPCELL_X1 PHY_EDGE_ROW_403_Left_1080 ();
 TAPCELL_X1 PHY_EDGE_ROW_404_Left_1081 ();
 TAPCELL_X1 PHY_EDGE_ROW_405_Left_1082 ();
 TAPCELL_X1 PHY_EDGE_ROW_406_Left_1083 ();
 TAPCELL_X1 PHY_EDGE_ROW_407_Left_1084 ();
 TAPCELL_X1 PHY_EDGE_ROW_408_Left_1085 ();
 TAPCELL_X1 PHY_EDGE_ROW_409_Left_1086 ();
 TAPCELL_X1 PHY_EDGE_ROW_410_Left_1087 ();
 TAPCELL_X1 PHY_EDGE_ROW_411_Left_1088 ();
 TAPCELL_X1 PHY_EDGE_ROW_412_Left_1089 ();
 TAPCELL_X1 PHY_EDGE_ROW_413_Left_1090 ();
 TAPCELL_X1 PHY_EDGE_ROW_414_Left_1091 ();
 TAPCELL_X1 PHY_EDGE_ROW_415_Left_1092 ();
 TAPCELL_X1 PHY_EDGE_ROW_416_Left_1093 ();
 TAPCELL_X1 PHY_EDGE_ROW_417_Left_1094 ();
 TAPCELL_X1 PHY_EDGE_ROW_418_Left_1095 ();
 TAPCELL_X1 PHY_EDGE_ROW_419_Left_1096 ();
 TAPCELL_X1 PHY_EDGE_ROW_420_Left_1097 ();
 TAPCELL_X1 PHY_EDGE_ROW_421_Left_1098 ();
 TAPCELL_X1 PHY_EDGE_ROW_422_Left_1099 ();
 TAPCELL_X1 PHY_EDGE_ROW_423_Left_1100 ();
 TAPCELL_X1 PHY_EDGE_ROW_424_Left_1101 ();
 TAPCELL_X1 PHY_EDGE_ROW_425_Left_1102 ();
 TAPCELL_X1 PHY_EDGE_ROW_426_Left_1103 ();
 TAPCELL_X1 PHY_EDGE_ROW_427_Left_1104 ();
 TAPCELL_X1 PHY_EDGE_ROW_428_Left_1105 ();
 TAPCELL_X1 PHY_EDGE_ROW_429_Left_1106 ();
 TAPCELL_X1 PHY_EDGE_ROW_430_Left_1107 ();
 TAPCELL_X1 PHY_EDGE_ROW_431_Left_1108 ();
 TAPCELL_X1 PHY_EDGE_ROW_432_Left_1109 ();
 TAPCELL_X1 PHY_EDGE_ROW_433_Left_1110 ();
 TAPCELL_X1 PHY_EDGE_ROW_434_Left_1111 ();
 TAPCELL_X1 PHY_EDGE_ROW_435_Left_1112 ();
 TAPCELL_X1 PHY_EDGE_ROW_436_Left_1113 ();
 TAPCELL_X1 PHY_EDGE_ROW_437_Left_1114 ();
 TAPCELL_X1 PHY_EDGE_ROW_438_Left_1115 ();
 TAPCELL_X1 PHY_EDGE_ROW_439_Left_1116 ();
 TAPCELL_X1 PHY_EDGE_ROW_440_Left_1117 ();
 TAPCELL_X1 PHY_EDGE_ROW_441_Left_1118 ();
 TAPCELL_X1 PHY_EDGE_ROW_442_Left_1119 ();
 TAPCELL_X1 PHY_EDGE_ROW_443_Left_1120 ();
 TAPCELL_X1 PHY_EDGE_ROW_444_Left_1121 ();
 TAPCELL_X1 PHY_EDGE_ROW_445_Left_1122 ();
 TAPCELL_X1 PHY_EDGE_ROW_446_Left_1123 ();
 TAPCELL_X1 PHY_EDGE_ROW_447_Left_1124 ();
 TAPCELL_X1 PHY_EDGE_ROW_448_Left_1125 ();
 TAPCELL_X1 PHY_EDGE_ROW_449_Left_1126 ();
 TAPCELL_X1 PHY_EDGE_ROW_450_Left_1127 ();
 TAPCELL_X1 PHY_EDGE_ROW_451_Left_1128 ();
 TAPCELL_X1 PHY_EDGE_ROW_452_Left_1129 ();
 TAPCELL_X1 PHY_EDGE_ROW_453_Left_1130 ();
 TAPCELL_X1 PHY_EDGE_ROW_454_Left_1131 ();
 TAPCELL_X1 PHY_EDGE_ROW_455_Left_1132 ();
 TAPCELL_X1 PHY_EDGE_ROW_456_Left_1133 ();
 TAPCELL_X1 PHY_EDGE_ROW_457_Left_1134 ();
 TAPCELL_X1 PHY_EDGE_ROW_458_Left_1135 ();
 TAPCELL_X1 PHY_EDGE_ROW_459_Left_1136 ();
 TAPCELL_X1 PHY_EDGE_ROW_460_Left_1137 ();
 TAPCELL_X1 PHY_EDGE_ROW_461_Left_1138 ();
 TAPCELL_X1 PHY_EDGE_ROW_462_Left_1139 ();
 TAPCELL_X1 PHY_EDGE_ROW_463_Left_1140 ();
 TAPCELL_X1 PHY_EDGE_ROW_464_Left_1141 ();
 TAPCELL_X1 PHY_EDGE_ROW_465_Left_1142 ();
 TAPCELL_X1 PHY_EDGE_ROW_466_Left_1143 ();
 TAPCELL_X1 PHY_EDGE_ROW_467_Left_1144 ();
 TAPCELL_X1 PHY_EDGE_ROW_468_Left_1145 ();
 TAPCELL_X1 PHY_EDGE_ROW_469_Left_1146 ();
 TAPCELL_X1 PHY_EDGE_ROW_470_Left_1147 ();
 TAPCELL_X1 PHY_EDGE_ROW_471_Left_1148 ();
 TAPCELL_X1 PHY_EDGE_ROW_472_Left_1149 ();
 TAPCELL_X1 PHY_EDGE_ROW_473_Left_1150 ();
 TAPCELL_X1 PHY_EDGE_ROW_474_Left_1151 ();
 TAPCELL_X1 PHY_EDGE_ROW_475_Left_1152 ();
 TAPCELL_X1 PHY_EDGE_ROW_476_Left_1153 ();
 TAPCELL_X1 PHY_EDGE_ROW_477_Left_1154 ();
 TAPCELL_X1 PHY_EDGE_ROW_478_Left_1155 ();
 TAPCELL_X1 PHY_EDGE_ROW_479_Left_1156 ();
 TAPCELL_X1 PHY_EDGE_ROW_480_Left_1157 ();
 TAPCELL_X1 PHY_EDGE_ROW_481_Left_1158 ();
 TAPCELL_X1 PHY_EDGE_ROW_482_Left_1159 ();
 TAPCELL_X1 PHY_EDGE_ROW_483_Left_1160 ();
 TAPCELL_X1 PHY_EDGE_ROW_484_Left_1161 ();
 TAPCELL_X1 PHY_EDGE_ROW_485_Left_1162 ();
 TAPCELL_X1 PHY_EDGE_ROW_486_Left_1163 ();
 TAPCELL_X1 PHY_EDGE_ROW_487_Left_1164 ();
 TAPCELL_X1 PHY_EDGE_ROW_488_Left_1165 ();
 TAPCELL_X1 PHY_EDGE_ROW_489_Left_1166 ();
 TAPCELL_X1 PHY_EDGE_ROW_490_Left_1167 ();
 TAPCELL_X1 PHY_EDGE_ROW_491_Left_1168 ();
 TAPCELL_X1 PHY_EDGE_ROW_492_Left_1169 ();
 TAPCELL_X1 PHY_EDGE_ROW_493_Left_1170 ();
 TAPCELL_X1 PHY_EDGE_ROW_494_Left_1171 ();
 TAPCELL_X1 PHY_EDGE_ROW_495_Left_1172 ();
 TAPCELL_X1 PHY_EDGE_ROW_496_Left_1173 ();
 TAPCELL_X1 PHY_EDGE_ROW_497_Left_1174 ();
 TAPCELL_X1 PHY_EDGE_ROW_498_Left_1175 ();
 TAPCELL_X1 PHY_EDGE_ROW_499_Left_1176 ();
 TAPCELL_X1 PHY_EDGE_ROW_500_Left_1177 ();
 TAPCELL_X1 PHY_EDGE_ROW_501_Left_1178 ();
 TAPCELL_X1 PHY_EDGE_ROW_502_Left_1179 ();
 TAPCELL_X1 PHY_EDGE_ROW_503_Left_1180 ();
 TAPCELL_X1 PHY_EDGE_ROW_504_Left_1181 ();
 TAPCELL_X1 PHY_EDGE_ROW_505_Left_1182 ();
 TAPCELL_X1 PHY_EDGE_ROW_506_Left_1183 ();
 TAPCELL_X1 PHY_EDGE_ROW_507_Left_1184 ();
 TAPCELL_X1 PHY_EDGE_ROW_508_Left_1185 ();
 TAPCELL_X1 PHY_EDGE_ROW_509_Left_1186 ();
 TAPCELL_X1 PHY_EDGE_ROW_510_Left_1187 ();
 TAPCELL_X1 PHY_EDGE_ROW_511_Left_1188 ();
 TAPCELL_X1 PHY_EDGE_ROW_512_Left_1189 ();
 TAPCELL_X1 PHY_EDGE_ROW_513_Left_1190 ();
 TAPCELL_X1 PHY_EDGE_ROW_514_Left_1191 ();
 TAPCELL_X1 PHY_EDGE_ROW_515_Left_1192 ();
 TAPCELL_X1 PHY_EDGE_ROW_516_Left_1193 ();
 TAPCELL_X1 PHY_EDGE_ROW_517_Left_1194 ();
 TAPCELL_X1 PHY_EDGE_ROW_518_Left_1195 ();
 TAPCELL_X1 PHY_EDGE_ROW_519_Left_1196 ();
 TAPCELL_X1 PHY_EDGE_ROW_520_Left_1197 ();
 TAPCELL_X1 PHY_EDGE_ROW_521_Left_1198 ();
 TAPCELL_X1 PHY_EDGE_ROW_522_Left_1199 ();
 TAPCELL_X1 PHY_EDGE_ROW_523_Left_1200 ();
 TAPCELL_X1 PHY_EDGE_ROW_524_Left_1201 ();
 TAPCELL_X1 PHY_EDGE_ROW_525_Left_1202 ();
 TAPCELL_X1 PHY_EDGE_ROW_526_Left_1203 ();
 TAPCELL_X1 PHY_EDGE_ROW_527_Left_1204 ();
 TAPCELL_X1 PHY_EDGE_ROW_528_Left_1205 ();
 TAPCELL_X1 PHY_EDGE_ROW_529_Left_1206 ();
 TAPCELL_X1 PHY_EDGE_ROW_530_Left_1207 ();
 TAPCELL_X1 PHY_EDGE_ROW_531_Left_1208 ();
 TAPCELL_X1 PHY_EDGE_ROW_532_Left_1209 ();
 TAPCELL_X1 PHY_EDGE_ROW_533_Left_1210 ();
 TAPCELL_X1 PHY_EDGE_ROW_534_Left_1211 ();
 TAPCELL_X1 PHY_EDGE_ROW_535_Left_1212 ();
 TAPCELL_X1 PHY_EDGE_ROW_536_Left_1213 ();
 TAPCELL_X1 PHY_EDGE_ROW_537_Left_1214 ();
 TAPCELL_X1 PHY_EDGE_ROW_538_Left_1215 ();
 TAPCELL_X1 PHY_EDGE_ROW_539_Left_1216 ();
 TAPCELL_X1 PHY_EDGE_ROW_540_Left_1217 ();
 TAPCELL_X1 PHY_EDGE_ROW_541_Left_1218 ();
 TAPCELL_X1 PHY_EDGE_ROW_542_Left_1219 ();
 TAPCELL_X1 PHY_EDGE_ROW_543_Left_1220 ();
 TAPCELL_X1 PHY_EDGE_ROW_544_Left_1221 ();
 TAPCELL_X1 PHY_EDGE_ROW_545_Left_1222 ();
 TAPCELL_X1 PHY_EDGE_ROW_546_Left_1223 ();
 TAPCELL_X1 PHY_EDGE_ROW_547_Left_1224 ();
 TAPCELL_X1 PHY_EDGE_ROW_548_Left_1225 ();
 TAPCELL_X1 PHY_EDGE_ROW_549_Left_1226 ();
 TAPCELL_X1 PHY_EDGE_ROW_550_Left_1227 ();
 TAPCELL_X1 PHY_EDGE_ROW_551_Left_1228 ();
 TAPCELL_X1 PHY_EDGE_ROW_552_Left_1229 ();
 TAPCELL_X1 PHY_EDGE_ROW_553_Left_1230 ();
 TAPCELL_X1 PHY_EDGE_ROW_554_Left_1231 ();
 TAPCELL_X1 PHY_EDGE_ROW_555_Left_1232 ();
 TAPCELL_X1 PHY_EDGE_ROW_556_Left_1233 ();
 TAPCELL_X1 PHY_EDGE_ROW_557_Left_1234 ();
 TAPCELL_X1 PHY_EDGE_ROW_558_Left_1235 ();
 TAPCELL_X1 PHY_EDGE_ROW_559_Left_1236 ();
 TAPCELL_X1 PHY_EDGE_ROW_560_Left_1237 ();
 TAPCELL_X1 PHY_EDGE_ROW_561_Left_1238 ();
 TAPCELL_X1 PHY_EDGE_ROW_562_Left_1239 ();
 TAPCELL_X1 PHY_EDGE_ROW_563_Left_1240 ();
 TAPCELL_X1 PHY_EDGE_ROW_564_Left_1241 ();
 TAPCELL_X1 PHY_EDGE_ROW_565_Left_1242 ();
 TAPCELL_X1 PHY_EDGE_ROW_566_Left_1243 ();
 TAPCELL_X1 PHY_EDGE_ROW_567_Left_1244 ();
 TAPCELL_X1 PHY_EDGE_ROW_568_Left_1245 ();
 TAPCELL_X1 PHY_EDGE_ROW_569_Left_1246 ();
 TAPCELL_X1 PHY_EDGE_ROW_570_Left_1247 ();
 TAPCELL_X1 PHY_EDGE_ROW_571_Left_1248 ();
 TAPCELL_X1 PHY_EDGE_ROW_572_Left_1249 ();
 TAPCELL_X1 PHY_EDGE_ROW_573_Left_1250 ();
 TAPCELL_X1 PHY_EDGE_ROW_574_Left_1251 ();
 TAPCELL_X1 PHY_EDGE_ROW_575_Left_1252 ();
 TAPCELL_X1 PHY_EDGE_ROW_576_Left_1253 ();
 TAPCELL_X1 PHY_EDGE_ROW_577_Left_1254 ();
 TAPCELL_X1 PHY_EDGE_ROW_578_Left_1255 ();
 TAPCELL_X1 PHY_EDGE_ROW_579_Left_1256 ();
 TAPCELL_X1 PHY_EDGE_ROW_580_Left_1257 ();
 TAPCELL_X1 PHY_EDGE_ROW_581_Left_1258 ();
 TAPCELL_X1 PHY_EDGE_ROW_582_Left_1259 ();
 TAPCELL_X1 PHY_EDGE_ROW_583_Left_1260 ();
 TAPCELL_X1 PHY_EDGE_ROW_584_Left_1261 ();
 TAPCELL_X1 PHY_EDGE_ROW_585_Left_1262 ();
 TAPCELL_X1 PHY_EDGE_ROW_586_Left_1263 ();
 TAPCELL_X1 PHY_EDGE_ROW_587_Left_1264 ();
 TAPCELL_X1 PHY_EDGE_ROW_588_Left_1265 ();
 TAPCELL_X1 PHY_EDGE_ROW_589_Left_1266 ();
 TAPCELL_X1 PHY_EDGE_ROW_590_Left_1267 ();
 TAPCELL_X1 PHY_EDGE_ROW_591_Left_1268 ();
 TAPCELL_X1 PHY_EDGE_ROW_592_Left_1269 ();
 TAPCELL_X1 PHY_EDGE_ROW_593_Left_1270 ();
 TAPCELL_X1 PHY_EDGE_ROW_594_Left_1271 ();
 TAPCELL_X1 PHY_EDGE_ROW_595_Left_1272 ();
 TAPCELL_X1 PHY_EDGE_ROW_596_Left_1273 ();
 TAPCELL_X1 PHY_EDGE_ROW_597_Left_1274 ();
 TAPCELL_X1 PHY_EDGE_ROW_598_Left_1275 ();
 TAPCELL_X1 PHY_EDGE_ROW_599_Left_1276 ();
 TAPCELL_X1 PHY_EDGE_ROW_600_Left_1277 ();
 TAPCELL_X1 PHY_EDGE_ROW_601_Left_1278 ();
 TAPCELL_X1 PHY_EDGE_ROW_602_Left_1279 ();
 TAPCELL_X1 PHY_EDGE_ROW_603_Left_1280 ();
 TAPCELL_X1 PHY_EDGE_ROW_604_Left_1281 ();
 TAPCELL_X1 PHY_EDGE_ROW_605_Left_1282 ();
 TAPCELL_X1 PHY_EDGE_ROW_606_Left_1283 ();
 TAPCELL_X1 PHY_EDGE_ROW_607_Left_1284 ();
 TAPCELL_X1 PHY_EDGE_ROW_608_Left_1285 ();
 TAPCELL_X1 PHY_EDGE_ROW_609_Left_1286 ();
 TAPCELL_X1 PHY_EDGE_ROW_610_Left_1287 ();
 TAPCELL_X1 PHY_EDGE_ROW_611_Left_1288 ();
 TAPCELL_X1 PHY_EDGE_ROW_612_Left_1289 ();
 TAPCELL_X1 PHY_EDGE_ROW_613_Left_1290 ();
 TAPCELL_X1 PHY_EDGE_ROW_614_Left_1291 ();
 TAPCELL_X1 PHY_EDGE_ROW_615_Left_1292 ();
 TAPCELL_X1 PHY_EDGE_ROW_616_Left_1293 ();
 TAPCELL_X1 PHY_EDGE_ROW_617_Left_1294 ();
 TAPCELL_X1 PHY_EDGE_ROW_618_Left_1295 ();
 TAPCELL_X1 PHY_EDGE_ROW_619_Left_1296 ();
 TAPCELL_X1 PHY_EDGE_ROW_620_Left_1297 ();
 TAPCELL_X1 PHY_EDGE_ROW_621_Left_1298 ();
 TAPCELL_X1 PHY_EDGE_ROW_622_Left_1299 ();
 TAPCELL_X1 PHY_EDGE_ROW_623_Left_1300 ();
 TAPCELL_X1 PHY_EDGE_ROW_624_Left_1301 ();
 TAPCELL_X1 PHY_EDGE_ROW_625_Left_1302 ();
 TAPCELL_X1 PHY_EDGE_ROW_626_Left_1303 ();
 TAPCELL_X1 PHY_EDGE_ROW_627_Left_1304 ();
 TAPCELL_X1 PHY_EDGE_ROW_628_Left_1305 ();
 TAPCELL_X1 PHY_EDGE_ROW_629_Left_1306 ();
 TAPCELL_X1 PHY_EDGE_ROW_630_Left_1307 ();
 TAPCELL_X1 PHY_EDGE_ROW_631_Left_1308 ();
 TAPCELL_X1 PHY_EDGE_ROW_632_Left_1309 ();
 TAPCELL_X1 PHY_EDGE_ROW_633_Left_1310 ();
 TAPCELL_X1 PHY_EDGE_ROW_634_Left_1311 ();
 TAPCELL_X1 PHY_EDGE_ROW_635_Left_1312 ();
 TAPCELL_X1 PHY_EDGE_ROW_636_Left_1313 ();
 TAPCELL_X1 PHY_EDGE_ROW_637_Left_1314 ();
 TAPCELL_X1 PHY_EDGE_ROW_638_Left_1315 ();
 TAPCELL_X1 PHY_EDGE_ROW_639_Left_1316 ();
 TAPCELL_X1 PHY_EDGE_ROW_640_Left_1317 ();
 TAPCELL_X1 PHY_EDGE_ROW_641_Left_1318 ();
 TAPCELL_X1 PHY_EDGE_ROW_642_Left_1319 ();
 TAPCELL_X1 PHY_EDGE_ROW_643_Left_1320 ();
 TAPCELL_X1 PHY_EDGE_ROW_644_Left_1321 ();
 TAPCELL_X1 PHY_EDGE_ROW_645_Left_1322 ();
 TAPCELL_X1 PHY_EDGE_ROW_646_Left_1323 ();
 TAPCELL_X1 PHY_EDGE_ROW_647_Left_1324 ();
 TAPCELL_X1 PHY_EDGE_ROW_648_Left_1325 ();
 TAPCELL_X1 PHY_EDGE_ROW_649_Left_1326 ();
 TAPCELL_X1 PHY_EDGE_ROW_650_Left_1327 ();
 TAPCELL_X1 PHY_EDGE_ROW_651_Left_1328 ();
 TAPCELL_X1 PHY_EDGE_ROW_652_Left_1329 ();
 TAPCELL_X1 PHY_EDGE_ROW_653_Left_1330 ();
 TAPCELL_X1 PHY_EDGE_ROW_654_Left_1331 ();
 TAPCELL_X1 PHY_EDGE_ROW_655_Left_1332 ();
 TAPCELL_X1 PHY_EDGE_ROW_656_Left_1333 ();
 TAPCELL_X1 PHY_EDGE_ROW_657_Left_1334 ();
 TAPCELL_X1 PHY_EDGE_ROW_658_Left_1335 ();
 TAPCELL_X1 PHY_EDGE_ROW_659_Left_1336 ();
 TAPCELL_X1 PHY_EDGE_ROW_660_Left_1337 ();
 TAPCELL_X1 PHY_EDGE_ROW_661_Left_1338 ();
 TAPCELL_X1 PHY_EDGE_ROW_662_Left_1339 ();
 TAPCELL_X1 PHY_EDGE_ROW_663_Left_1340 ();
 TAPCELL_X1 PHY_EDGE_ROW_664_Left_1341 ();
 TAPCELL_X1 PHY_EDGE_ROW_665_Left_1342 ();
 TAPCELL_X1 PHY_EDGE_ROW_666_Left_1343 ();
 TAPCELL_X1 PHY_EDGE_ROW_667_Left_1344 ();
 TAPCELL_X1 PHY_EDGE_ROW_668_Left_1345 ();
 TAPCELL_X1 PHY_EDGE_ROW_669_Left_1346 ();
 TAPCELL_X1 PHY_EDGE_ROW_670_Left_1347 ();
 TAPCELL_X1 PHY_EDGE_ROW_671_Left_1348 ();
 TAPCELL_X1 PHY_EDGE_ROW_672_Left_1349 ();
 TAPCELL_X1 PHY_EDGE_ROW_673_Left_1350 ();
 TAPCELL_X1 PHY_EDGE_ROW_674_Left_1351 ();
 TAPCELL_X1 PHY_EDGE_ROW_675_Left_1352 ();
 TAPCELL_X1 PHY_EDGE_ROW_676_Left_1353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_2000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_2001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_2002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_2003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_2004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_2005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_2006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_2007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_2008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_2009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_2010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_2011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_2012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_2013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_2014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_2015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_2016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_2017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_2018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_2019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_2020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_2021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_2022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_2023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_2024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_2025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_2026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_2027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_2028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_2029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_2030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_2031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_2032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_2033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_2034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_2035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_2036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_2037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_2038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_2039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_2040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_2041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_2042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_2043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_2044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_2045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_2046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_2047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_2048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_2049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_2050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_2051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_2052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_2053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_2054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_2055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_2056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_2057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_2058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_2059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_2060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_2061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_2062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_2063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_2064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_2065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_2066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_2067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_2068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_2069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_2070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_2071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_2072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_2073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_2074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_2075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_2076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_2077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_2078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_2079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_2080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_2081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_2082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_2083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_2084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_2085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_2086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_2087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_2088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_2089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_2090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_2091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_2092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_2093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_2094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_2095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_2096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_2097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_2098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_2099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_2100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_2101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_2102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_2103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_2104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_2105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_2106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_2107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_2108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_2109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_2110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_2111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_2112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_2113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_2114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_2115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_2116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_2117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_2118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_2119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_2120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_2121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_2122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_2123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_2124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_2125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_2126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_2127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_2128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_2129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_2130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_2131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_2132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_2133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_2134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_2135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_2136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_2137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_2138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_2139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_2140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_2141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_2142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_2143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_2144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_2145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_2146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_2147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_2148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_2149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_2150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_2151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_2152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_2153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_2154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_2155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_2156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_2157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_2158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_2159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_2160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_2161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_2162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_2163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_2164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_2165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_2166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_2167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_2168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_2169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_2170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_2171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_2172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_2173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_2174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_2175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_2176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_2177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_2178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_2179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_2180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_2181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_2182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_2183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_2184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_2185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_2186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_2187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_2188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_2189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_2190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_2191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_2192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_2193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_2194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_2195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_2196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_2197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_2198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_2199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_2200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_2201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_2202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_2203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_2204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_2205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_2206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_2207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_2208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_2209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_2210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_2211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_2212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_2213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_2214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_2215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_2216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_2217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_2218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_2219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_2220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_2221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_2222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_2223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_2224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_2225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_2226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_2227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_2228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_2229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_2230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_2231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_2232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_2233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_2234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_2235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_2236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_2237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_2238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_2239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_2240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_2241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_2242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_2243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_2244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_2245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_2246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_2247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_2248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_2249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_2250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_2251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_2252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_2253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_2254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_2255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_2256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_2257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_2258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_2259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_2260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_2261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_2262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_2263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_2264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_2265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_2266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_2267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_2268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_2269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_2270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_2271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_2272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_2273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_2274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_2275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_2276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_2277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_2278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_2279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_2280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_2281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_2282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_2283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_2284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_2285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_2286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_2287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_2288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_2289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_2290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_2291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_2292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_2293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_2294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_2295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_2296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_2297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_2298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_2299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_2300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_2301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_2302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_2303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_2304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_2305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_2306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_2307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_2308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_2309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_2310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_2311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_2312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_2313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_2314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_2315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_2316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_2317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_2318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_2319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_2320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_2321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_2322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_2323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_2324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_2325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_2326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_2327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_2328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_2329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_2330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_2331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_2332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_2333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_2334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_2335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_2336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_2337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_2338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_2339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_2340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_2341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_2342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_2343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_2344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_2345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_2346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_2347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_2348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_2349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_2350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_2351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_2352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_2353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_2354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_2355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_2356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_2357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_2358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_2359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_2360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_2361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_2362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_2363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_2364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_2365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_2366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_2367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_2368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_2369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_2370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_2371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_2372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_2373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_2374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_2375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_2376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_2377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_2378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_2379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_2380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_2381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_2382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_2383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_2384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_2385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_2386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_2387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_2388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_2389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_2390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_2391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_2392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_2393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_2394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_2395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_2396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_2397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_2398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_2399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_2400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_2401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_2402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_2403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_2404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_2405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_2406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_2407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_2408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_2409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_2410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_2411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_2412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_2413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_2414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_2415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_2416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_2417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_2418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_2419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_2420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_2421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_2422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_2423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_2424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_2425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_2426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_2427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_2428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_2429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_2430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_2431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_2432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_2433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_2434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_2435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_2436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_2437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_2438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_2439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_2440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_2441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_2442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_2443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_2444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_2445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_2446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_2447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_2448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_2449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_2450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_2451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_2452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_2453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_2454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_2455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_2456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_2457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_2458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_2459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_2460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_2461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_2462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_2463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_2464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_2465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_2466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_2467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_2468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_2469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_2470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_2471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_2472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_2473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_2474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_2475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_2476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_2477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_2478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_2479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_2480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_2481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_2482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_2483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_2484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_2485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_2486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_2487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_2488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_2489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_2490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_2491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_2492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_2493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_2494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_2495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_2496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_2497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_2498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_2499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_2500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_2501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_2502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_2503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_2504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_2505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_2506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_2507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_2508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_2509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_2510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_2511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_2512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_2513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_2514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_2515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_2516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_2517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_2518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_2519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_2520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_2521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_2522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_2523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_2524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_2525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_2526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_2527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_2528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_2529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_2530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_2531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_2532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_2533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_2534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_2535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_2536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_2537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_2538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_2539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_2540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_2541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_2542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_2543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_2544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_2545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_2546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_2547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_2548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_2549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_2550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_2551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_2552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_2553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_2554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_2555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_2556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_2557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_2558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_2559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_2560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_2561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_2562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_2563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_2564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_2565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_2566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_2567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_2568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_2569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_2570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_2571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_2572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_2573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_2574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_2575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_2576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_2577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_2578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_2579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_2580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_2581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_2582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_2583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_2584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_2585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_2586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_2587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_2588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_2589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_2590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_2591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_2592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_2593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_2594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_2595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_2596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_2597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_2598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_2599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_2600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_2601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_2602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_2603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_2604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_2605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_2606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_2607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_2608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_2609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_2610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_2611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_2612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_2613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_2614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_2615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_2616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_2617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_2618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_2619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_2620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_2621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_2622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_2623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_2624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_2625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_2626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_2627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_2628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_2629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_2630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_2631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_2632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_2633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_2634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_2635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_2636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_2637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_2638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_2639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_2640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_2641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_2642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_2643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_2644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_2645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_2646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_2647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_2648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_2649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_2650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_2651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_2652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_2653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_2654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_2655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_2656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_2657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_2658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_2659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_2660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_2661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_2662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_2663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_2664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_2665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_2666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_2667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_2668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_2669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_2670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_2671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_2672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_2673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_2674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_2675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_2676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_2677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_2678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_2679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_2680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_2681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_2682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_2683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_2684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_2685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_2686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_2687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_2688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_2689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_2690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_2691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_2692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_2693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_2694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_2695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_2696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_2697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_2698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_2699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_2700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_2701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_2702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_2703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_2704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_2705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_2706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_2707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_2708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_2709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_2710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_2711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_2712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_2713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_2714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_2715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_2716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_2717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_2718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_2719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_2720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_2721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_2722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_2723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_2724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_2725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_2726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_2727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_2728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_2729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_2730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_2731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_2732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_2733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_2734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_2735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_2736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_2737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_2738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_2739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_2740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_2741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_2742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_2743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_2744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_2745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_2746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_2747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_2748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_2749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_2750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_2751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_2752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_2753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_2754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_2755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_2756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_2757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_2758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_2759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_2760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_2761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_2762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_2763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_2764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_2765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_2766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_2767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_2768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_2769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_2770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_2771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_2772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_2773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_2774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_2775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_2776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_2777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_2778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_2779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_2780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_2781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_2782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_2783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_2784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_2785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_2786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_2787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_2788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_2789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_2790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_2791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_2792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_2793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_2794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_2795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_2796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_2797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_2798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_2799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_2800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_2801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_2802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_2803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_2804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_2805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_2806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_2807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_2808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_2809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_2810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_2811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_2812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_2813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_2814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_2815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_2816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_2817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_2818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_2819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_2820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_2821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_2822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_2823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_2824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_2825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_2826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_2827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_2828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_2829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_2830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_2831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_2832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_2833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_2834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_2835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_2836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_2837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_2838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_2839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_2840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_2841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_2842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_2843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_2844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_2845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_2846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_2847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_2848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_2849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_2850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_2851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_2852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_2853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_2854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_2855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_2856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_2857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_2858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_2859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_2860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_2861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_2862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_2863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_2864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_2865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_2866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_2867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_2868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_2869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_2870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_2871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_2872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_2873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_2874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_2875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_2876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_2877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_2878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_2879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_2880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_2881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_2882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_2883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_2884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_2885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_2886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_2887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_2888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_2889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_2890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_2891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_2892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_2893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_2894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_2895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_2896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_2897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_2898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_2899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_2900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_2901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_2902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_2903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_2904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_2905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_2906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_2907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_2908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_2909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_2910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_2911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_2912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_2913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_2914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_2915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_2916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_2917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_2918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_2919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_2920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_2921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_2922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_2923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_2924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_2925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_2926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_2927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_2928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_2929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_2930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_2931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_2932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_2933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_2998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_2999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_3000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_3001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_3002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_3003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_3004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_3005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_3006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_3007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_3008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_3009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_3010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_3011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_3012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_3013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_3014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_3015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_3016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_3017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_3018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_3019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_3020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_3021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_3022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_3023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_3024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_3025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_3026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_3027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_3028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_3029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_3030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_3031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_3032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_3033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_3034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_3035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_3036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_3037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_3038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_3039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_3040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_3041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_3042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_3043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_3044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_3045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_3046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_3047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_3048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_3049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_3050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_3051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_3052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_3053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_3054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_3055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_3056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_3057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_3058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_3059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_3060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_3061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_3062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_3063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_3064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_3065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_3066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_3067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_3068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_3069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_3070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_3071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_3072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_3073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_3074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_3075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_3076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_3077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_3078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_3079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_3080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_3081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_3082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_3083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_3084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_3085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_3086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_3087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_3088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_3089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_3090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_3091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_3092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_3093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_3094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_3095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_3096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_3097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_3098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_3099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_3100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_3101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_3102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_3103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_3104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_3105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_3106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_3107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_3108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_3109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_3110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_3111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_3112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_3113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_3114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_3115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_3116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_3117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_3118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_3119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_3120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_3121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_3122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_3123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_3124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_3125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_3126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_3127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_3128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_3129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_3130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_3131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_3132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_3133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_3134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_3135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_3136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_3137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_3138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_3139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_3140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_3141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_3142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_3143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_3144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_3145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_3146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_3147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_3148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_3149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_3150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_3151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_3152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_3153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_3154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_3155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_3156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_3157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_3158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_3159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_3160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_3161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_3162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_3163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_3164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_3165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_3166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_3167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_3168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_3169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_3170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_3171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_3172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_3173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_3174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_3175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_3176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_3177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_3178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_3179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_3180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_3181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_3182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_3183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_3184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_3185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_3186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_3187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_3188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_3189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_3190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_3191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_3192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_3193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_3194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_3195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_3196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_3197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_3198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_3199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_3200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_3201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_3202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_3203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_3204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_3205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_3206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_3207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_3208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_3209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_3210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_3211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_3212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_3213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_3214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_3215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_3216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_3217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_3218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_3219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_3220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_3221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_3222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_3223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_3224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_3225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_3226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_3227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_3228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_3229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_3230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_3231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_3232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_3233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_3234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_3235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_3236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_3237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_3238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_3239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_3240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_3241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_3242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_3243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_3244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_3245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_3246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_3247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_3248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_3249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_3250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_3251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_3252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_3253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_3254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_3255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_3256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_3257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_3258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_3259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_3260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_3261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_3262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_3263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_3264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_3265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_3266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_3267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_3268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_3269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_3270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_3271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_3272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_3273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_3274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_3275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_3276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_3277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_3278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_3279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_3280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_3281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_3282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_3283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_3284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_3285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_3286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_3287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_3288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_3289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_3290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_3291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_3292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_3293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_3294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_3295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_3296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_3297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_3298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_3299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_3300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_3301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_3302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_3303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_3304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_3305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_3306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_3307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_3308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_3309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_3310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_3311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_3312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_3313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_3314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_3315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_3316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_3317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_3318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_3319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_3320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_3321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_3322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_3323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_3324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_3325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_3326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_3327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_3328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_3329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_3330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_3331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_3332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_3333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_3334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_3335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_3336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_3337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_3338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_3339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_3340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_3341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_3342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_3343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_3344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_3345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_3346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_3347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_3348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_3349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_3350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_3351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_3352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_3353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_3354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_3355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_3356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_3357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_3358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_3359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_3360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_3361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_3362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_3363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_3364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_3365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_3366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_3367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_3368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_3369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_3370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_3371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_3372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_3373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_3374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_3375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_3376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_3377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_3378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_3379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_3380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_3381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_3382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_3383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_3384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_3385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_507_3386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_507_3387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_507_3388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_507_3389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_508_3390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_508_3391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_508_3392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_508_3393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_509_3394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_509_3395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_509_3396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_509_3397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_510_3398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_510_3399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_510_3400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_510_3401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_511_3402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_511_3403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_511_3404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_511_3405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_512_3406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_512_3407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_512_3408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_512_3409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_513_3410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_513_3411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_513_3412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_513_3413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_514_3414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_514_3415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_514_3416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_514_3417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_515_3418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_515_3419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_515_3420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_515_3421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_516_3422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_516_3423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_516_3424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_516_3425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_517_3426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_517_3427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_517_3428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_517_3429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_518_3430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_518_3431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_518_3432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_518_3433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_519_3434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_519_3435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_519_3436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_519_3437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_520_3438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_520_3439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_520_3440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_520_3441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_521_3442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_521_3443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_521_3444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_521_3445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_522_3446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_522_3447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_522_3448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_522_3449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_523_3450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_523_3451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_523_3452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_523_3453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_524_3454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_524_3455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_524_3456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_524_3457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_525_3458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_525_3459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_525_3460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_525_3461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_526_3462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_526_3463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_526_3464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_526_3465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_527_3466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_527_3467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_527_3468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_527_3469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_528_3470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_528_3471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_528_3472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_528_3473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_529_3474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_529_3475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_529_3476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_529_3477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_530_3478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_530_3479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_530_3480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_530_3481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_531_3482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_531_3483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_531_3484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_531_3485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_532_3486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_532_3487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_532_3488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_532_3489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_533_3490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_533_3491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_533_3492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_533_3493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_534_3494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_534_3495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_534_3496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_534_3497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_535_3498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_535_3499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_535_3500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_535_3501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_536_3502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_536_3503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_536_3504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_536_3505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_537_3506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_537_3507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_537_3508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_537_3509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_538_3510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_538_3511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_538_3512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_538_3513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_539_3514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_539_3515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_539_3516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_539_3517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_540_3518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_540_3519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_540_3520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_540_3521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_541_3522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_541_3523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_541_3524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_541_3525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_542_3526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_542_3527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_542_3528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_542_3529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_543_3530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_543_3531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_543_3532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_543_3533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_544_3534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_544_3535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_544_3536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_544_3537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_545_3538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_545_3539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_545_3540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_545_3541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_546_3542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_546_3543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_546_3544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_546_3545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_547_3546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_547_3547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_547_3548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_547_3549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_548_3550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_548_3551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_548_3552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_548_3553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_549_3554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_549_3555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_549_3556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_549_3557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_550_3558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_550_3559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_550_3560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_550_3561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_551_3562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_551_3563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_551_3564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_551_3565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_552_3566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_552_3567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_552_3568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_552_3569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_553_3570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_553_3571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_553_3572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_553_3573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_554_3574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_554_3575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_554_3576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_554_3577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_555_3578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_555_3579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_555_3580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_555_3581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_556_3582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_556_3583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_556_3584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_556_3585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_557_3586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_557_3587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_557_3588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_557_3589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_558_3590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_558_3591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_558_3592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_558_3593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_559_3594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_559_3595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_559_3596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_559_3597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_560_3598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_560_3599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_560_3600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_560_3601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_561_3602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_561_3603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_561_3604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_561_3605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_562_3606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_562_3607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_562_3608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_562_3609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_563_3610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_563_3611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_563_3612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_563_3613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_564_3614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_564_3615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_564_3616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_564_3617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_565_3618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_565_3619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_565_3620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_565_3621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_566_3622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_566_3623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_566_3624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_566_3625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_567_3626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_567_3627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_567_3628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_567_3629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_568_3630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_568_3631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_568_3632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_568_3633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_569_3634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_569_3635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_569_3636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_569_3637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_570_3638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_570_3639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_570_3640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_570_3641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_571_3642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_571_3643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_571_3644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_571_3645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_572_3646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_572_3647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_572_3648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_572_3649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_573_3650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_573_3651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_573_3652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_573_3653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_574_3654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_574_3655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_574_3656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_574_3657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_575_3658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_575_3659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_575_3660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_575_3661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_576_3662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_576_3663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_576_3664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_576_3665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_577_3666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_577_3667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_577_3668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_577_3669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_578_3670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_578_3671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_578_3672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_578_3673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_579_3674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_579_3675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_579_3676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_579_3677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_580_3678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_580_3679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_580_3680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_580_3681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_581_3682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_581_3683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_581_3684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_581_3685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_582_3686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_582_3687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_582_3688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_582_3689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_583_3690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_583_3691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_583_3692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_583_3693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_584_3694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_584_3695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_584_3696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_584_3697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_585_3698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_585_3699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_585_3700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_585_3701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_586_3702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_586_3703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_586_3704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_586_3705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_587_3706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_587_3707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_587_3708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_587_3709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_588_3710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_588_3711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_588_3712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_588_3713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_589_3714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_589_3715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_589_3716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_589_3717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_590_3718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_590_3719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_590_3720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_590_3721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_591_3722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_591_3723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_591_3724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_591_3725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_592_3726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_592_3727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_592_3728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_592_3729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_593_3730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_593_3731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_593_3732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_593_3733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_594_3734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_594_3735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_594_3736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_594_3737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_595_3738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_595_3739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_595_3740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_595_3741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_596_3742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_596_3743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_596_3744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_596_3745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_597_3746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_597_3747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_597_3748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_597_3749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_598_3750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_598_3751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_598_3752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_598_3753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_599_3754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_599_3755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_599_3756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_599_3757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_600_3758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_600_3759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_600_3760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_600_3761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_601_3762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_601_3763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_601_3764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_601_3765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_602_3766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_602_3767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_602_3768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_602_3769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_603_3770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_603_3771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_603_3772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_603_3773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_604_3774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_604_3775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_604_3776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_604_3777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_605_3778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_605_3779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_605_3780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_605_3781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_606_3782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_606_3783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_606_3784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_606_3785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_607_3786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_607_3787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_607_3788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_607_3789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_608_3790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_608_3791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_608_3792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_608_3793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_609_3794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_609_3795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_609_3796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_609_3797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_610_3798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_610_3799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_610_3800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_610_3801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_611_3802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_611_3803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_611_3804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_611_3805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_612_3806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_612_3807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_612_3808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_612_3809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_613_3810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_613_3811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_613_3812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_613_3813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_614_3814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_614_3815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_614_3816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_614_3817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_615_3818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_615_3819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_615_3820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_615_3821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_616_3822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_616_3823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_616_3824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_616_3825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_617_3826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_617_3827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_617_3828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_617_3829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_618_3830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_618_3831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_618_3832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_618_3833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_619_3834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_619_3835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_619_3836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_619_3837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_620_3838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_620_3839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_620_3840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_620_3841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_621_3842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_621_3843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_621_3844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_621_3845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_622_3846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_622_3847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_622_3848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_622_3849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_623_3850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_623_3851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_623_3852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_623_3853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_624_3854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_624_3855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_624_3856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_624_3857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_625_3858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_625_3859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_625_3860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_625_3861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_626_3862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_626_3863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_626_3864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_626_3865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_627_3866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_627_3867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_627_3868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_627_3869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_628_3870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_628_3871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_628_3872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_628_3873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_629_3874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_629_3875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_629_3876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_629_3877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_630_3878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_630_3879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_630_3880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_630_3881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_631_3882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_631_3883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_631_3884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_631_3885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_632_3886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_632_3887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_632_3888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_632_3889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_633_3890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_633_3891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_633_3892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_633_3893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_634_3894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_634_3895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_634_3896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_634_3897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_635_3898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_635_3899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_635_3900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_635_3901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_636_3902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_636_3903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_636_3904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_636_3905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_637_3906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_637_3907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_637_3908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_637_3909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_638_3910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_638_3911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_638_3912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_638_3913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_639_3914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_639_3915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_639_3916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_639_3917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_640_3918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_640_3919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_640_3920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_640_3921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_641_3922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_641_3923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_641_3924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_641_3925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_642_3926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_642_3927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_642_3928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_642_3929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_643_3930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_643_3931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_643_3932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_643_3933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_644_3934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_644_3935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_644_3936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_644_3937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_645_3938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_645_3939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_645_3940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_645_3941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_646_3942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_646_3943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_646_3944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_646_3945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_647_3946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_647_3947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_647_3948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_647_3949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_648_3950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_648_3951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_648_3952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_648_3953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_649_3954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_649_3955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_649_3956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_649_3957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_650_3958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_650_3959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_650_3960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_650_3961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_651_3962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_651_3963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_651_3964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_651_3965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_652_3966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_652_3967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_652_3968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_652_3969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_653_3970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_653_3971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_653_3972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_653_3973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_654_3974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_654_3975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_654_3976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_654_3977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_655_3978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_655_3979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_655_3980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_655_3981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_656_3982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_656_3983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_656_3984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_656_3985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_657_3986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_657_3987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_657_3988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_657_3989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_658_3990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_658_3991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_658_3992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_658_3993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_659_3994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_659_3995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_659_3996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_659_3997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_660_3998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_660_3999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_660_4000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_660_4001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_661_4002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_661_4003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_661_4004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_661_4005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_662_4006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_662_4007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_662_4008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_662_4009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_663_4010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_663_4011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_663_4012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_663_4013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_664_4014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_664_4015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_664_4016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_664_4017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_665_4018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_665_4019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_665_4020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_665_4021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_666_4022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_666_4023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_666_4024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_666_4025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_667_4026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_667_4027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_667_4028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_667_4029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_668_4030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_668_4031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_668_4032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_668_4033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_669_4034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_669_4035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_669_4036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_669_4037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_670_4038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_670_4039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_670_4040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_670_4041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_671_4042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_671_4043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_671_4044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_671_4045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_672_4046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_672_4047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_672_4048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_672_4049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_673_4050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_673_4051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_673_4052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_673_4053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_674_4054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_674_4055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_674_4056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_674_4057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_675_4058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_675_4059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_675_4060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_675_4061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_676_4069 ();
 BUF_X32 max_length1 (.A(net10),
    .Z(net1));
 BUF_X32 wire2 (.A(net7),
    .Z(net2));
 BUF_X32 max_length3 (.A(net5),
    .Z(net3));
 BUF_X32 max_length4 (.A(net6),
    .Z(net4));
 BUF_X32 max_length5 (.A(net6),
    .Z(net5));
 BUF_X32 max_length6 (.A(net7),
    .Z(net6));
 BUF_X32 wire7 (.A(net8),
    .Z(net7));
 BUF_X32 max_length8 (.A(net9),
    .Z(net8));
 BUF_X32 max_length9 (.A(net10),
    .Z(net9));
 BUF_X32 max_length10 (.A(ground),
    .Z(net10));
 BUF_X16 wire11 (.A(B[9]),
    .Z(net11));
 BUF_X16 wire12 (.A(B[8]),
    .Z(net12));
 BUF_X16 wire13 (.A(B[26]),
    .Z(net13));
 BUF_X16 wire14 (.A(B[24]),
    .Z(net14));
 BUF_X8 max_length15 (.A(B[23]),
    .Z(net15));
 BUF_X8 max_length16 (.A(B[22]),
    .Z(net16));
 BUF_X8 max_length17 (.A(B[21]),
    .Z(net17));
 BUF_X8 wire18 (.A(B[20]),
    .Z(net18));
 BUF_X8 max_length19 (.A(B[19]),
    .Z(net19));
 BUF_X8 max_length20 (.A(B[18]),
    .Z(net20));
 BUF_X16 wire21 (.A(B[17]),
    .Z(net21));
 BUF_X8 max_length22 (.A(B[16]),
    .Z(net22));
 BUF_X8 max_length23 (.A(B[0]),
    .Z(net23));
 BUF_X16 wire24 (.A(A[9]),
    .Z(net24));
 BUF_X16 wire25 (.A(A[8]),
    .Z(net25));
 BUF_X16 wire26 (.A(A[31]),
    .Z(net26));
 BUF_X16 wire27 (.A(A[30]),
    .Z(net27));
 BUF_X16 wire28 (.A(A[29]),
    .Z(net28));
 BUF_X16 wire29 (.A(A[28]),
    .Z(net29));
 BUF_X16 wire30 (.A(A[27]),
    .Z(net30));
 BUF_X16 wire31 (.A(A[26]),
    .Z(net31));
 BUF_X16 wire32 (.A(A[25]),
    .Z(net32));
 BUF_X16 wire33 (.A(A[24]),
    .Z(net33));
 BUF_X16 wire34 (.A(A[23]),
    .Z(net34));
 BUF_X16 wire35 (.A(A[22]),
    .Z(net35));
 BUF_X8 wire36 (.A(A[21]),
    .Z(net36));
 BUF_X8 wire37 (.A(A[20]),
    .Z(net37));
 BUF_X16 wire38 (.A(A[19]),
    .Z(net38));
 BUF_X8 max_length39 (.A(A[18]),
    .Z(net39));
 BUF_X16 wire40 (.A(A[17]),
    .Z(net40));
 BUF_X16 wire41 (.A(A[16]),
    .Z(net41));
 BUF_X16 wire42 (.A(A[15]),
    .Z(net42));
 BUF_X16 wire43 (.A(A[14]),
    .Z(net43));
 BUF_X16 wire44 (.A(A[13]),
    .Z(net44));
 BUF_X16 wire45 (.A(A[12]),
    .Z(net45));
 BUF_X16 wire46 (.A(A[11]),
    .Z(net46));
 BUF_X16 wire47 (.A(A[10]),
    .Z(net47));
 BUF_X8 wire48 (.A(A[0]),
    .Z(net48));
 assign Prod[16] = s2[0];
 assign Prod[26] = s2[10];
 assign Prod[27] = s2[11];
 assign Prod[28] = s2[12];
 assign Prod[29] = s2[13];
 assign Prod[30] = s2[14];
 assign Prod[31] = s2[15];
 assign Prod[17] = s2[1];
 assign Prod[18] = s2[2];
 assign Prod[19] = s2[3];
 assign Prod[20] = s2[4];
 assign Prod[21] = s2[5];
 assign Prod[22] = s2[6];
 assign Prod[23] = s2[7];
 assign Prod[24] = s2[8];
 assign Prod[25] = s2[9];
 assign Prod[0] = v1[0];
 assign Prod[10] = v1[10];
 assign Prod[11] = v1[11];
 assign Prod[12] = v1[12];
 assign Prod[13] = v1[13];
 assign Prod[14] = v1[14];
 assign Prod[15] = v1[15];
 assign Prod[1] = v1[1];
 assign Prod[2] = v1[2];
 assign Prod[3] = v1[3];
 assign Prod[4] = v1[4];
 assign Prod[5] = v1[5];
 assign Prod[6] = v1[6];
 assign Prod[7] = v1[7];
 assign Prod[8] = v1[8];
 assign Prod[9] = v1[9];
endmodule
